`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAw1/4wNkWeivqsXy8ekYN1vJlV1Iod5PYGgK7SadacgKlh5usEz4jj3m5NqLPcS
qkbcUURT3eX7pA9K0TZp/C30DVAYDZfQInnTjfwy3EHKBjG6ynH/Ef0X6JxoYoFw
knnHBGgS7HgEhW1EG6ntcjoJKPqr2SIlPJiqd1Up2r1Q1gzmMGSGqJdjFRg2qiYD
tIyiQkWvkw9a7EbJqKivP41aU+lAVJMWDl3WtLdy/qVnKvq0NFXefgLeNINUAziw
AeRBVvj5x9qkmsdloxYE8NXi4fpvvvDD+IODgyz1FMB0IlWsXa9qoiguv//IpXXV
L0R24LgGUW1XkVXWCknmvs3Ffp3uBN7t6em6gcURiYAhM5vn3VzMQ+NhRwdTQ8DJ
TrHNGm5Vf4tIOXAB+Ywt33/vfi65aI3A9tpqMDzZWGAxlSxtFpAVBGN/nR0ssEmT
A2E8JNoQ2MpZ3HzDWSrMfQRgOXLgaBOxdl39U8nf9K0+sUAFHw6gv4d+LPBgDrqw
gsOC0xGwEoYY0iOK9QZKk4Y82twkWVd8tzsFMpMgXRpYdL7u83t7Pi0+dOjGYNIH
u7YHz2eRZ6Lzcqb2Bn0j6D/u/zOzzQPS/ViHDqqV+5wcibIO6FZZAG0zvvFftaNg
ah2foEmVqh3uyGFy7IQSSXNkhgfPc7WafHesHwCtitHQKQ0kT2gmVZ974ORnI34r
qrYhWxujYQiGqANnz6SPnarN0AswQPlOEJidqCLFVjgRSAnd8P9cfGmUJcfwIhki
OKokflTqVFEHgtvpOiuVVWozv8OUvoipJCnJHIl6C/nXlz8oYBGrOhjqitEwtGfZ
CtxHTbRza/SKNj4LBkM9ns2nNyLUxA9XA5r01CyNmmXWazBO27OjO39d/JmYGAQ0
eVvqNilc9BS3DK+kDklX+omzz44TlwXf1VkUiZewOAu6RYCV+ND+XUmzk6HD88s+
WrAQVHcm5hqdIntf06g85FTfHUwTad6tKz7cEa9d2a8=
`protect END_PROTECTED
