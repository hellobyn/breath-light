`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8AazN4y3O/EHqbKHSWL7JNzqFbQPt8KXiCsUY8P5ivTFofIW109Bmyj84mlVfsF
UuWZrOhXGzZm1prta78vKGrv+N/vUVu8st0mMos1ijA4NUsZj1c5atgRE1M7d/e5
+a7eZOVovupgszAahr3U0vDINKaQgiKGEHvvANufxDGeezMF0igPPsQQZvGDi/jo
gTnpgyTQemqrJfMaVZjWFb/z6L5FfkcyeM1Pjp1gjVkoY60lxjviX3CP5LiHZ6TP
mTL3929B7AVA1N+9/1D6qMflhredbm3IZ74PLPaj8zy7BbSZjxIGKShSDxNthGLG
VgYEUGhu+EIdR9SdjByiydmIlC/1mnyy49bL/scQ0vF16DX4t6zM8d2ezPgYVT27
98MeRsGkW1wnL8IFLFfjQZxgs4ZvtPr/hAfYnLj8e/yEW/TnByXqG+Vx+AE2u/io
97kTSYPScLRdfjUV16n7J8lExpv34ChKY6OLwPLMRa1SPoJpAxrT7wGtZLLec88v
T9sYWdw6uxUpWk+Rx11qMLwvH7bY/7ldQwRWsUP4Qt3dmpnraCTcV0bktZySDlrw
fiDi0Vhat/l1QGbK57ZjaccZNWqMD8DPybkqLd93StagltS2y11NKSzNNueBiiYQ
wzdTtwzChPQQohb6awAC/ovZSg4dDKWdRSfOqGf7CYhWIztAOkEiZBBfUYA1MVXh
WNx4o0RuRMl8qqkoou1uAKBfmfiRfqVXOQ35jc7UIUORORutHOjOPdSzTj2wpEDs
T9Jir//EBtf4mhUSapSDzFL/3eGzPKu82TYdmYUIUkBQL4jEIg17szXFZS4lOUwx
KUChEGpfsVx4WE9kFfFHaVP/+xy17w7bdzfZd+cIbhj1KNsd4VZ+7M/BY1YNLmZN
n7QmKConyo7lUgXm2v+L8s/Dob6Tgs89NP14fhjlDbfzmAX1LG9GYwI1fMx/cDvx
hKYDsfbiOFBJVz0MhJt3ANnhUllcI8Sw9YSjl9AAOi6gEGntHlxbSTiWMc3bDYYx
Yek8cg55aSDiAtJ88w9xhlOn3sXZz9U4s10vknghO/GEfRYBae8vIqkV2KHfG6Eo
nXp/sqg3bL76ejg0wDQdakWkKbpjzbDjnGR8gNjTRFS/TpZAWiUMO1bhWGBhrhbS
U86Qbk9oQDEqkpFOEK3+lzugcTx7xbkJSJXnf8h0a2ClmvXUrog5CSXlI1iFLZNd
V38So/swb65UXLfb5cYNvYLLMNEewIyUvYsIeoT6QTZ5mLJ5gDOnH2BKrXIzufaV
4kqg0cjbcq245YQrtxxfXBJdwCOqroidVvkWW9WSvLUdbb8orijAdYSKkyTPJMGk
FuuuI+L1Su2jkcAeIuw2EI6eDABvKEi+/nPffaTGLi1DfzNzSWSBpjGc1tb6gZ5q
Tsz4BRS2C86l5mCxtZDcDUH/gF88cqv0Z5Uc4MJFIhr86jc8phCN060luvqjbk0W
QJy06YBmm1I0OTdjuoHbdgcjp2tiWW8pOO4TbRkFp31LyzJZFapxcO8tGOeoWCNm
PkJQXTAa1ZDNUk72YCi9Frn2ikT0NkNTz1ZfxTuHXRF7jZl91sHEq/azN23MT86S
fMTt/JpJeqgnCuaMKW6x8z4BBprzEVcrMsuH6At+fOlaXsN6a6y8trDXzoS3mMvq
HRAd8M6jv86Lqgz54XGfgZPD/yLG+ikqsZ2Ffof65JlRPul7THauxSee15RY8FE7
QGPynfkaUHTIDyx7IlLwUO7ogSNWt05M53QPClK1K7IquyKGg7IBTFdmoudShWpU
mvJR+C1C0jIbgsZFo7rx5iQTaWCb9vGVHZYgC99qkqVE09pTVJivqczdO7kMiNzL
er+oAHO2s74tFoyrOb74iOsuC5obztFlm4yr8utoVUb+iZau/1BunaYjUEYZStoF
h0iHrbrBjCjNHCHcksKTw7heKIr+nVXBhLIqSFvXGATSJabUZeLpVCQ1zbUn4RIm
3Y4cLeATnQjJF1dHSd2TqV7J0RM957EJlkG/41fb2jYe7vn5ZYeTafKyiSnS70xR
akC1WSpoRTm7TJwbZ467i5CGctfAVjOJijrbYkjH8idtNgHvHzRHwnu6p+u9gmF4
UyStyWiLn24LNiZtSVugFjoswFhCyF3N22OVFtIUg3jen5nS3AIENWUAeONi2IR7
cJjPTfCMwXhdP+pkJMxEkGsWEtp9p+m046BSVBamUEYA38meENZU07asGHGqpjsy
ud7p8zPz55C3b7VJesk5/etQVQWjyzrT1jhB/hSDZsofCc7O1FbRqGkPgjxfS4Uu
lvBYGLBWE19jWzxVGKvyLdWshgzFsp8UiAfB9bVqJoxpzBI1jze/7+RVMiSuAZj+
XQSzmCIHs+bfgl4DJkfqx6lm6kuqOzpeUqUNiZG4ORYNTxzBKLzm+DkGXh5sGWNu
rAagcGKELtAjiGpS20xVHQ==
`protect END_PROTECTED
