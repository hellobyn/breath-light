`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXdLhLsJHkiiCD7iosQ6cotnDomrQZZP4CSaLu0/LSH7WSUCMv9O+A/3zh5sm4Vc
bcolL6DbIjKHC9g5RrliEELDgUusHKJ5C6sGerx/BaPuxlaw7/9swQ8BO4ne4wTj
fHuxI7AXAYHb/BuEHUr8Elzopq6QPidSxsKX/Nn0Nhdl/2l3w8mDX8cNTcFoJiE6
a7IhtoB48s6WDqk459HHYQAn3CTwBdhRIGYXCcg1Q8+X1bqr7CCLztT7EZmqvq8q
ObGZQbHuEuWjdzTnNnoC7rI+hhY8KHEZzi41PLcwm2jQLOJFKshYn1r0d3wI5qVd
UH0D9r0mKaDxrAJl4I7uT7/XgkfFjhnWrzSKaevySska3hteyIx2ZGKzMc8WaxJ9
uLjdnG0deQGH6B9yA+D1bTSxKxOAjMGJJ4dHb2gXLjU2tkfHYWGiOJOpkQLs1h8l
NdgkNJ8gDvsI3h/8KrQ+qS76/VAPEtyAEO9ZwrYAWrmlTxZXUPJjdLrwJs8Tdaes
XZ7oFezRKXcQgliStNC3wAcRYazTBiTGPaUXR3B7kHn1pwf0HXDOlLDmHa5D2kwb
NRSFU9COiAYCo1HwVSgzKb6sYRFDk53AsS7rBGb9D3o3fHjyD6ylUbero6Od42t5
z3R0GBsHkeTDj4gS0HcK0n3A+lD5go6oVyizDSqKMXRmSf13pOiOuWh37Z1YCe28
ClYG4G3xRsP5sldIzI9s0YcmUhK8ACwEhYZf/4T6p3zn2R1LsGjVM5LPnZPb3wo6
Xb4qPQ29Pwjjhpoc2YYkPeFNUCQ4OJBBVYukud8GAzIY3VomwwYjngeGCjHNzIwJ
PkFb2+SNFDK6zIIW4mtPtXfgOZCUHzAChWA7h46XhvNC0bEG4lNveLhkgJoUKixY
`protect END_PROTECTED
