`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEStOMUEUbiE8rxXe7MSr6TRmqLXzwTcw8H4HPuzd3N27a8d2+hWdjC347Cfdrm3
bAcdHp+as8tlYshvwH8uPs0Kc8YHkFFWtuXhLrQYDHoGeN6TEGRHlcMPzcu3oxnL
UuBQAe58nblbA/ex4oBy2W4kVSiIYMnX9U2+Q8EnLeA9Lt7DTb9WYNOIDkO+qQwg
ot32TnPyjGX79aByUOqdcwDPkC6Pcm6g/lWPsrCjF5vJ5vo5I6fEj8wUxhW22Ln/
1v8a6Bx9S6ECjIdW0PHFK/3SJb7TFUMh0sBZbeBT7olfDJNMWbN0qoDpBhd83Zhh
7o9iEp2yvhCF0F+dJlmS7SLbwg/YG0ABEetFcAz4ySC4EZYMCbvpNKX1t3BT58su
Ywj6vRqqthQHmpARrJkXh/NXAzEANtZqf/Ki4/EjxUNXLAeSyPA6tIF40HpNAPJ7
/2eMdAWUu0rqgCEA72GG49JuUYjiFomJd8qN7WIvXVWQ3fXvgdWERyK9EdeTSNE2
Cff8Upn7Z1iB4gObsoj2NQfUaQHjHiQny2jczfQUYVk1w2qiwjfZy0gr+CkezuDR
EDvuemRMgkfpF+wqGSOFqVGI2d3JXiW4PZF7GRXsiSWsVo/u4BavUgeoSrAkFXtd
dKVx/XYO9L0X8ep7Z+Bc8eNwTpaB1m9QG1TsTsR2T4Wejs1SCMZWjaNCYuDAvIFj
/f5AuW7OpfP8BU6M8P4nEEw+KoQ9qoum96Bttxfvy7XpRJ1ZXvmNYDLhnMsiQqlV
tDH7UIYeurN9hn7Xeydhww8XEHMCByZWGkDODWcJAw2oYjsiVK4GAt8zCcJvakjp
f27tsb64rGfFyfyvIjqigfwt1N40uHL2nmn81bX5f9jFnOE+b6o+GfUirRTklLR1
RrWIN50Lfbq3NUmmb+PYVp27HDQrV9ZgQyGjnD9NYloCCGD/DEIXQVp2i6D+ZqNh
9oqboZAot+qYERD9joNRdCzDscqGoNhbvvk5wNr5avBgDpW/a21DjamdidoYuDMH
`protect END_PROTECTED
