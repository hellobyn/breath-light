`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHeWR3mbchgHaEzidz4sK3k+jALXcbr6OvY/XqnKgQEU1GNWqwASmNNMPm/35h1b
fNZJvbC+SnQi66ZWbh1Gtk61MszbzBCKMDv0Sbn4YAFhXx2L4Rerd4Yf7uzla1ec
qv/epzPLv3wsxq03eg9NlQlwgDYUZvKfz0wrZmud5T6Qc3jnaSiJBV62MjHQrXYb
ncbWLntk4Br/PSwlikZ4xnWLCE3X+rSlq6Lti/rt6xeKnVpfiMYDreAUhkjx6sSR
BAFSzPe2FODafX0iEBLHTGnLYm/kvBMxzk6sXCUk+8WMJpF6MbVwLX2E9YPF+7Sz
NuWtPreo0hFVGRM/lxm8OhAyY2pfh2buXz7s0ViUGqFGEi/Dz29KamDm0yHm9vAw
KCaNAz+NQfSetmH9Dpx/HH9mGsoeMl6QdgcKfyZTAh+QSjhQpWs1N1p3alYKPBao
sYnEt42kbLXfEJxyoaVlkv0tFTde9NAX1WWONJDFYXOj17Tn5WRg2HBZnlk88nHM
kupk8xO8a7QurZ1fmQIwr3iCI5x+VshQMfptrXZyYRs7yKWqAStHIweuPGfSrJ5v
`protect END_PROTECTED
