`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRyKOJIplo/yor1fMff6s9fI1ZOjJAiGojLvExjqb6aX98CSVhsDol3ko1IdUE5C
9B1ymXDH82NinYuOpdp+ZLuRIp/62yFZ5rUIeuavSZGsWQiOQfW5htNDon5zfosJ
Trbw8QVzcFYExHVaAQwv0RIqI+sp24r2OqGwNl9dlEwHRZB0i4ESxND00tyl/+Ff
5WiTPJX1zMfZBbufoeoFX+wIf8f+9H8qDWkqTggoClKThJyDU+59Cp47JkQkKji8
N8xh3Y+uR//clzqiniQJxS2qaflRdcUP/Cp1CvfMCHhe+eUDD/UwxMh8BpSv630P
D9OhjXEveR+jtKHNqJp0BwOMWSMc6KS/9VeN7nxi5Vs+dFlgvCEL2Lj/GwCbZ4H9
O6XFn4M11Fs5Aya8kZ7pcb/3EAsvdorcN/T1sbgsGHIrRG+6uvLTYWiFW+aatCi+
x4zCmuzX4bBd32MKsiHs/88aXTHnlbbEq//evcnR4awp1YIDXXA2tNYb/CHLXSkF
RHdFWIlKBLWkAAOwIgICLaxRXuhmp4ms8LDX0DsudV+ncM8C09bSiGBJwa63j6GY
37kfhbgvhvix7hksUqpQH3+yJnj6K+YZ/kkVcOG6QBrBXMFKFf+1Cu7JKLKi95k0
ZM6xl1pAYRhDDaMcQJOY73NHQmHb/6EVxhjLuo0TBFKQnPp7uL3ryJs59mLLq9bx
JZX2oiQtsD+nq2P9ZwRHO+bKkWHlbsv43Eef3IoPTZdLJy5pcwgn1iOX8R50R/4Y
9wpzTx4exmZp86Yumc8+0zrtZU0ettCRMctRbrI2B9mECMSMmB+nDRw4qsT7Je4j
j8ogWXYMkqsweAdSv2hGBpS+BQ+wCjS65TKgcsLlEflIacEN8pfk5xbPtK82El7G
J4eJf1PamKHr2r+DCXM2V9IVBFz6jdP5vOcveIurw1U=
`protect END_PROTECTED
