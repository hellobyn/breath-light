`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hw3j04BMdlWE4vUw4CvjMS/Fvifma6QrE9HX89FZQJyWfNJxEQ4wan83y2N1wcGo
JZV4acMEeyEA17ciQ9/3eKffospQQsSFkIPNmqTADBwdT1HkJgbxh2KpWzxyKdVq
RzPXmm3LY3CooKg1T7pQzlKOAarIiUjrDOeBQ7mgZjeleSrWIpNQT+Wchu9QXVTd
TeEtyoRy89XfCmTO+zsvzROqO+82zJn5Qqv4rXg+cSLYtdI7RV/pn4AVHlKs2EQo
FhqjHoOgCkCaZGdzVs7SgNob/uIQyo0TguVEkPzWMYtjOsdLi5wewAY2YerWPNK0
TQe8+guePEkUL/QzldpLRdHsqLe+OqiVmTuGZDSO4pIkZid1IjwiojffUdel5y+d
9r6i1kdICwS7sIuZ/sw7wXa9JmPeOeb+OVYQrfxL5NY/ND0NpRtC+lPOTjfqRvXY
kHSupLIiTnd9/4Xu2kRLuKYfpK4iWbwpDtlgpNVsH++7cL8XTk9XZixdsn+elaiU
Jwfr1LFZ6eJZF1PnqxWpjA==
`protect END_PROTECTED
