`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gg8vQphQj0GgjmosxGTMxfmEdqCF2QIDEaExGzuy587T36Gpu4RIBksHB1wxuGDZ
mxMTC6QESV0Y8RUvJCCX3IpA+kmol1mjDsfiZKA0gWjl402lAYoxcEniTQeLTdUR
t5JEvln6lIORyiH/MudnwHh8jzdDKSaihr5C3IgQl0aO1V5bslO/NrBtDNq7Lm68
u29BoVHDiRoFDfk69TnIHYZfMn2MNR4RgNMX9x6FUe5Taii56scshdMN6f3hUrn2
W0ivmYO8nv7+5Qq6QAmvWylAFhRm26PzMp+R880UqBinWRMaSzmTIOXn4JAweIzS
aff+t4p023Bnw1WApX7n9M4CQ8oN7YdLTQKcpfcYjGux19GV1s3WOEcIuSCGjk+S
csXLtc0dnJJajR8Bj9YDu+V5o/yAo3uA1tr2P2In02eZM57TphlO3wq2CjimYCXt
57q04gSZO/ncWjWAI/L9WsvfsGKT9/Gmb4eBv/FllUAII/oUR1K5zpZGi48FcFnL
BijPnYwvdf6k7B8IbpkD8jMmK4Jp5weUnhki57ZYQ9DaWsCZyJtMds2qAIJvVSIs
4gNtr8P7IhKWCPlGVEx7VS6EiyEziRkP7/B1rfJ9bHFzZQtvF7nSzse46UcCIJeQ
RQ+OhcNQ7fZrqW5Aw2TAFdrDkIX+0Ix41N01+FMvJJ7a3N4w1Wkz7Eo8FNCQbEba
Sjd3strvVVBxRPURu4OlU+ughRkQ8lITHGK+kNTgOjlKaGL9dgIWHlk6MVicQOse
RZm73ckNMtajrYKFXk4V9FXm84wn8TzL36wUkcnShFGiXSiExdgJ7Pb//Ba9ZngA
hHAP+fO5v8b9mXUPn9eNkF+1ulGj5jTo3xe9KiLuj8oSeANvV4sX2NeeZzcCAKTv
1QYkxHKMnD8BjmvQcXr/KUcONNJG/RD6jYTN860+0dzf/ObkRCl2o6cN4tvBMl6o
V4pHwmlzjwB5Rx/qVKrtRM7EMeNun+z/UmNYcNgJYfvYNAwdZJaKmXFeYjjT18AI
obXsbDH3hbN/HcfX9epYqTFfh+eRn0NBsrqFF+psBlsaGdVtmr/+fCuECHeD020A
hRo8xhDFO/cVVs4B9/jcqBRwNFG9dMLfrn175OstHi4=
`protect END_PROTECTED
