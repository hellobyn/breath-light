`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glWo4QkXuiEzvRJ0mFCjG2nyyGW2l88wctBswQ45xGsYLEYuT5vzG4ugG6w8JUno
fpsXVmwHUrPCCX1FYRVqI0bI1JPooyJPX+dOOvEnWSWnFQzib9I0kgwv1haphuDz
p3riXfrE2hT0+NGV0fUSovajb5xts0zWxCm7FIUOzU/cJPUkIN9MXmIQ7SkMP5Fd
r44qd88ui9A0FadV/bh5VUnL1hhTpSvokE3iWg0SsiJcoFTX/eM3xAW6kCRsYM+P
NezYyMAUvV7pkUyZGbLuj7gPA505d32taexKYYCkn4yaa0EQEdzp9yo9Ie81OXz7
M6KmPct7t1CJvXkxbOAVUD6iDKLOubs2I1/kNHuo4+GSysp9AtrnyITr/37LeayV
cT2yNpVOIlAWJqkyfjaUVbAgpeYq7Oz5FyXVyOhNOi9RF0RJs+j7qKZ15kPakdQy
xwuF+kX5CCJjtAgdF4c7rp3sIh6BE+8ApvEazxNn5IX2YxJXds1Lowf/I9FXEnNU
Mpoga1RjfzgAJ4j8yUKnvKYNi5VQo+s3xphiViIR6m8Xqf2hGhli1AE6SN5IxBpT
tBM8b4ptt5qfRorW/LcnzSTPlKpLabYKQeoIIVx/ep4f0+kmbYkXwy0dfhN+EqvM
idGiryoPopHahgmI/9qlZ24KW/1cHiE3+7f8xPdIzd9RAtsy1GjYpk5IIcD6jnl9
ysXPlre2I60OvprjYAyoxlnlVt5Fti1OWEtAJLuAcWt0VseZrU6GS6f1B6/CDAG1
CG8x8RmFkAFU7mJ5yNESqAemRqwILkmXPSVo3N7LCz7mWA0/3KG+kSDipheXJhk7
odp70UVBFPl5thVooWx0MJ9lEMVhX6pbCzjIUvXJj2rYny1tu+K/AB4qxFw6+yDx
S6fRSDeOzCRWYTYYHhc25rde7pYBNOVJGFyyR4ZWxUTOIuUfFseKhh+caD/J7zFk
dshKGad11i5hk28F1ETrR+3Xz4mlmL8CQU6gtCy1OtLLMat8l4IIePwdSY1OeHB4
fQ6d9Wfzbf/D76nL113mzhBXKykzXm+s5HK/uogCrL6KgXN38wW449BmLrCoN370
CPs/nUEUGIJf3hTGK5uV9JXpoSQg5l62kWMQzayKKjt0mV+aQS35aWrj7IYukra1
nrJRyvjkw08dMpC1JVyMvw3dmw0v3NjctsX8ffAFubYa3eiW7mPkdF58UsM/o/YB
sW757Z/LiT68aIRI9H0iyE4dPPTkgrMBbDrFf3KIZ81j4A2XQt9/M5u6AeglKZ0f
ZZlDd8MlEOASy0DjWeSkDIFITLZUQkyWmDmK1oMS20RBaNM7hVWr8RYzGRHC0NTc
B4aZSLWnNvXeANeFXBnF5e/uyFfH82yqsJxVkWcKd4DObs6WsR51Hcv5Y5SCAOyN
mvmVcX+toduZ21790tJ4iihqw2nbF7QZmsjvD4VatcUhVhSBLSlswgN/6GzHGBSj
aosHFINtCBjku5OpjmnO4ueIEYuuhGkZQ9h6p3uoTQTx/cXw5jMvbn6lvZ+f0uY/
qMlEooPk/C0yHJitztwGOkCXPR8r/laUFLDpiR5wDvK546PuiqaYlpUhIG4UgtwT
kg2Odk6/k1yxbGHkvk+bTvpIyz2iUiyfa3pxAw0s1t7MI0s6v9C8X5qM3TSuAcLh
hUeCvzKrFKWGVltJpkt0qjNFQgi6oSYB2VU1QPxuvzb7I6K/s53fA8o0+wOzwsr+
b05I+t5FerZ/xtSZm1TdWBXZNwe3S0129e+lrWRp/ka0MiKrS4DBSmkGFrJZhvCT
/URBUX9KVO35GYrXED5LHvw6Tjh8zmedFPm3BpdLc5gfvyvLb0aZwywJJjMjTmjN
3tPHM5wueJijPCN+ro6YF6valOiG8oOuXWXnHjg/yzMJkDi8f7ION8Gd2tIVW78J
XbUgLIYKUWO+TZtRFWTrjpMPiQrcubM0jpaXSxSdBKs4i3m/cGp3DHTlh+pHA8X+
5XHnJUWxEmJmYnmz5MeyYP8Fe4oGPGnXXwX/NMpafwmiRtiqtSzC/1MOuV5uiHNP
jFmiLfH8joR3N3vYio23OX8/OuGExk59f/wnRQVSKhWmZqzywtDZr2Y2GKyG/TgO
j96AjgD5MoeXONpBFQ5ViOV8YWI54ILqd9xWcanACn0etCVjXuCywLkKpfGU7h3y
hTEzcecXdfa/PHhvhGCAsKlksfM5F87clBhbe4Ep6I56gX1L4hZzr2XodCGRZ4Sd
hkHXh5FDI+SuOTPz/ddDKoagJmsXI0RDbHbdcJY/zeakIi44uDsqQ1Ob6bq892oI
cmkmwvX4VW8CG2gslgZrd2qBNW8hDvL1guf4gSupMkzNHVAh9Ntm1/AWS1qhXUzX
jZum5dVgWK8i40baTc2Q8MTBAIwpJ2w14y1PRit1LD3T7DkyFeSsNlJE1+ti/Bfi
1EgE2zPlzm4AlrnebEX9D6d45mwEpG9ImLIzzQ6KtCa/ZI/9BG0iYLNfEpXvvsRI
jWWlsAcCm9xzVW3ckrE3L07lKuYhhJzsdr3iNqpApqGtqyyOtqH6BnjhXyoGKXg1
02r2RVaZF+yNoJy1xcS2YyOqltM/PjymLu/sKw/8YTOvqrBaBWS9iR+mrOJ8ie/I
Lzj1T8ct2/9EOtq18eKPtDuvlHrE8ULHBOvaflVUkwEKTohX8qpv6djKZc077WGs
Khjmu50ACGTCmp7HZ8/VD/kingWEbufY+qZWbNaCgBVapoNLWQ+r81r8FNMRyc9h
VYqYT+8MPsFgnppIHWIciHCIklowXjPY4GjdbvZdgd3aA+lJuxR8R59D9UPT8AXK
c9VBdXqneslla48vI3n/3FyN17aO8TXvAAjBEmMtWqhBULQBwVsX2O26G1AZYLwg
hyO1lZQAJCG++lo1xqQ4l9mSW0XIZ1YcEf9rpCbFI7dj7iXJCSHAsSQzBTByKtSS
UHtHbpgB4QTaxP84dVSNt5F2VvVdqpMT1MBBcGX6bRAkcWieYsshwNzJA3HsT+HB
QaOTw7Aa1m1gEHJi4YqNCk8rnQFOPrvlTCasBHRwL7iQc9Dror97KtbKQx+ZMw7M
wA7xGcrkzSYQwHNyUPNazlZ4ZcRne6sdaiNheyEwIEJq4JQG1UiuTBrYQJWxbxM9
DHiJGXB8QrHIM7X3m0ZNW/9tGNCNgTc3R7g+OW+0yLT9rs5+amPdDiy3/htNSTsg
JsIxfvy3NISkdzxb1tU0UfGzGOZunqK80dDU1NBwPNIctdLZyrMbuwNXEi/tVsHF
eVcGJC0LJxBGBNVFYJVl2pA5iQveRK8kDC/tKix3mLcOhNpIJZ8/F1sgCONoI+ZX
gzU8oj5nuct8oeah2tBv4XFxK/tcr6sMjEdNKIv7HMvJgan55NCJZb3Kbp3kda2C
+eKdgnhcOtFaSnn04+6CGCLqKl0yBOqbcbFJUCKhAF19jNNpDLcM56ZaixXKrvII
/bTpaO+0qyMHBEgyJAhA7BBUitFVfJC1aiyyEodjCRuM+E5hY4K1xSbuk1IUm6Ug
/5yLa3MGZblSb6+oLB6XnPbMkE8AtAI108BzTcAYHhdoo9xP4h4lyFGzR3m8LRgy
CSpdrBF4drFxqAbEzpOjpUfbHx78YdU6ECZUuAGZgnYtSV09Q2FZuns+wJfg496a
hlM2Mg5oLCs5fMWOCjmlFosc0Q9oFXqhlpu0pXjp7D8psISyp5oaPtvJHrLvXq5z
3OLDO3uAoQN10AtjQM95m3TH8mepLXwqTF+buUY25f2Q9hrgm7TpIYEL1vo/HNJX
MAav+B0t7VH1eZgIqp+INwe31rLIQ8fLnJbFrvbLH0wsP+swStH7azULeG4+Hmnb
loAQlaAIha8vh47DQHZTKAu4nee/wQgyNpYQQGfsbSTMvWCUN3VEjn52opMrsdDm
i12VQbUCTrQmsnBD1sF33Rg/FnG16PJDaqqgH5N6a8zlEDSRqKDtFRzruAnFhuVX
PDBg9GXmFapOUGd8I9/aJwEzAu0GmPnejZecanqcnXD/PjfD2qrl6oKOUpEG6Mb3
H22/qWgoKXuIlKB8Y/YptQ9FV1W1nHY5mEi++OV8lSBtglYCaQqvsTIEInBIb1Sy
T5F0uxhMBFy7DbWWx0frhrOq9Av6NoDOd1q96zQT04YmLKbvkCgNCBZnTGPazu2o
OKMied6PeyokgRECmf7i6gmtA+08v9vYBYVxgsZyiWsCxneRGCGB19rd/eZwRysE
lUujvy43XC6jSmQoHBeKcfCDubKeG/lc426KPn8IFBtdAN17Oonn9K0I5jfjAAWY
U9zzb5VjDWGw9931zmrXamf0PY9f1q4AkzBW2TCA1bUh7PDASAfwR23yYUKVe+R6
3yKwIaA3IDn9zlW2s3PWvFyKo3BUOa+Wf2E5rD8YXKa/IV3aawpQAjPC4wbcAzsB
vjQ34/n0UXaUZPIqcHmJF5O9cCtDKNkUFqIvnFZcYvEC0fvI5b446JvqYYG4nusR
CHYX/OgVmQCeekVfcaNCYS4nSwZMBXOhmGSv69d51Ok5otJ88T6BYTAHSMjGtwEE
sOoiojjsVid4L/bqcFtEIYGu0Z09ziiHL65heP8Ey5Xb/FEtIFa6arpw4LEOlwCD
CsMswsEonwKIe+Rd4fVsCyg6CiVLb20xQOmSK+QCSOn/D31t9M8jBM7SH9+mG/ry
jR6RNcX0tmDFXVQSgko46NlpDILIoBEx7JbkIUjCDzCzK9+kuuSlZc7anfPIU8fu
3FruB0hjk3/A5sZ2Q9ookVIAWpo2YrhGhAXj2C0w3YJeJcTIZCa+3VVzZD56apCM
H00p74snqda35WV8/Nh/OALpz+wR7yZFt2cuC+Njbv1PdwVZIMHjMOtKErXmabrj
LHdP+8SUoIj46LCsQ877O9qMyzo/hIIX262ekXzfPK8WyX1GhdN5/sEf9W8Amdpb
+Gck6/vcIr3kgYVOnMbe9pe9vZcQpfuOBYLEfdT5Pa4+ThAqh6WNriEhU3qk04pP
gTQkhEgDQpJLWi+oPycawEr1QqPuz7+1fN1yb2f2+fOtNaBzj19cBnOYu3sDinsM
/3WWXP37kowcir/8MAXjRcPYPl/TKurI7FPzo9hE58jl/GFRvQ14K4dBlv2h29jA
njBJZAvmk62qh+zppSmP+VCG2ngaqaFSn8VKWU7hZ3yCJvuDXMtboFiStQwPicVJ
qPjoDTqlj9N+usAk7nUF0sQ0z+44PYcpi9FlVXCZSHkPGWf9pak4xlnTDJ3rRWE+
Bl06Tv7w4BDXPHtu9GymObdIkk1mE8RK0qSAM1xR/a2oIMqfzxOCaZcPUr1JFL7G
P64nVkckIkX25eL7Ak29876B0ySVrCJqnXdb26/0IJb1BYD4HJIJBxiB9KM4w0/J
MwJUAyf9m4lU/fTA4u3sN5zPc3K/fdFG3nliqfYht2ude4bt5s7im0nWVcJMAQvR
SAnx4VaZZwKaUMhlbG0pjdbiSvkiWApaSYcGF2rmdYuR44aJAy2xUyNbgCSHhwG0
ZhLqpzy1/k/5XCqAYrH8TRIW8QBUSStaTobC9q2UFwzJkDEQZyamx+3yHHLQKL+q
CGJhDlSKwzuvpdyLKKhVazreyOBJgqE4QUrlxDZiTCx2VlEw/oe2OgmNkC9P097t
R+MteY5s8vDoUKtsJlFe6eK9lEiK3dARH9+lABpZMgnV7gKvECcFlTifTl4DDLFZ
VwQ6D1U6w1njojrlGrtFnUbu4Vgce/J5bmv7b/kSVPCAbSP30Oscpbv5sHFoWaLk
vnzgshFBv4KA8dscbcilYscU49b/jEposZ/3eaymE6vGzD5XoK83wHqnTolDtLYZ
ZeNMmLlLG3k5B7PVxMZArqR0fK435WNBzUGgwJp8D7MpkQlVUC5uPBm2WLJ1deoT
YwL5I5mrAb+rj7HmLeCWkTOiCGzhynZo8eboDlXKfPqZWeHbwxEJEE2bH3MY0yRg
NnSbKG1jyDyTgxOghjQ3YP1fNCco6zg7VfoMATrtycH541s1NiDVUGqIFbeDOjYE
gTA4F7UuX3RAnWWKSUEP762oWnTuSAdnnbyhirO9fzFduOBKjguf2TOea6QX15Za
Km8v+wbxOCK2G7YU1eDdHsYrqSS9CNH6prCw7etvnIvfljVCo/kzFP5gndIh0uou
2Sh09Ch75EZ05HIrxL8EqB4ZruE2LkTO3P+YYjq740BGHXfo7BSjeklCc8kK1EN0
sruvp/fwvhoLWvGP6AKAYB1VCXYsvtZTALExnJU8QzGPBg4AYjxrtntbnv7RTSpE
t2Kdj780Kh3pZq2151KOhuhPiV+LIu+biRG/5me5XncFldl3c3w5I0msUq+M5QA1
HN/x0Zrtfdu7pj4E5H2UQdO2eV0w1Km8cSZhRvH8Pdlbwd0vB1ljpweVw1e3XWuf
rSbY/kLD9VXZTgYF7wCcIlk/3asuxrWlvZ/V1ngnSdqfbZE3JEIb+ERAW8/5pBUq
lhMu+y1W/NcaJ9qP1Hq/5pRVrWFmTg0BOShmLZonWqt0I5rxlOvSwY7zIifo671O
Z15hGB0L4fxVJJWtXzJ4c47rcwW85HKOyi/B4XRQ72EFzCLEh1dnsp2fGeqnklLS
8Tg63ASseIneuiij8AnKYSLWtlj/wTwGe4a+KR0qH/BfKDXlrwQ233H54sW/EJE3
tjZcQpABmM3e1ojD8jrCXWdoJbEOeCyq8oLpj7F+ckzBAQhfnB0dbNFMc4yQH2hF
lbJ/EHTGWub54gaU8zrd8YSdlTi4E+agElHiqB80HEmkyEDHL92Ng5cMBZQXzF6C
dugJ7W8JWP8Gf4vQSIxubTd5y22ZLhwgcOPiV0F1LDa01bYXHVb7e2282nnBK+lw
0GMsb8J9ZfGhC5XR1XfNOgia6Kr5H8Rz6xkLtFa7SnAdqg0PoF+tjovmeyBuGXSc
XP8oM8ru1d9UKBEBAU9MHEDFMBYX6Fieoc9LoY9NoOCO8rugBlyLCnxA4lqlr1XQ
mJ5kD0p1CD4ewFt611xDNRaJQ4yra6whDvEitDysv1/NHXEUv92Nk2w4FRlb5yo5
MapCAn6AcB3DozoT8SY4XuMGmCCkTEgc2V+Z/pADfCnkc4gEUMSo7T6w+KXxE/Mp
y/MaZcRXaPYSH9Tv5eysCjgBTGzYx4wSv4T009ZVW+/0JTnVN6AoM5Ez/8muh61X
loXJTx29VK9i76Pb2SWyl7Q+rnyUKOkDfM6qsq3MYoRHbUPRufQGs3yN6kZxJqFx
2WRHySGXGqME8n3gYYJ7zuJ2vTFFoKN/cHrZLZwSnn7VVeVch+lmKq/Aj7gEcNW5
Zht1pjYTkZqGAEm3K6g01t3682bibxt1i44yKgLXxVRIbtgZ5hS+BGmOzRSRoR8Y
qFc1FgRn/pkq7nivYzw1BPdOFWe0ZBwdaNzONVZfrOvQRKkCjZ31OpeR4wtXWAmI
X++TaKitnvq/UUaZ5x8jWRWFX4+XX/6t8orDr4ZeRcA+4e5Q0xmjrhfbkmObMHQ6
oMd7FpmpB151iu26t6OoDO9GIUMwSj+qza+HnaOT58EC5wsgi6us7GiC0MMrSl5J
PXr1lOdVB/i5133iwQ5HXPfmy7ti61pZ14StEx0l798kQTDfIICw3xdsUBKeagQg
CkWO4Ksh0zNFdKpPqXT36o1odl5kdIPAEQF2MZmrfc1axklvhQ/J5lDJ4HOyalu9
4SiTeaRUzw8+F6cHGFJSltfbp75H6yQKo8ETUdqjbNUeNsa4ZeoeYjdedkcOZYcT
A56wUnLD6CTwHxtfe0SKdqf8YlCyNbyvXhX//yT0oe3IYxUiLvibFsXtIbjAF7pH
oE2gUeGzPX3lTmdPnz8Fgqny2BJuJG+9pU5NjWkJkDvwLkp5BReNIArvkzFXCaTs
P2aNlH39wu1DnL/9P1lAMPq4no2618rjXNqLYpOMPjze+eREh+O1GNYPQXJr2W1F
2F2ZKi1AQrmnck6DJZdfXCxfSHGvrdX1arES2K//666EAo1cRrMeYhsFXMZN/FES
4DdQ7xCE9bmS1jqVN4WmY3RU09CdFdy+mbsRcVtDnQvKWkU+0a8gbhcDU8mYkLEz
U4FQ2jdHHWdOb5JcnEa9/8wCMAPjzTqfVBTRwsVNGjw/YiTT19Iew4U+Pf6Vf5iR
lI9voKfSGpHKV7PhTiaIbgeHa+Z/OsCVHgGgM6MlCNjwMGz2wy3/xlBpAn/PjD4B
qkIQu+idRDW1QgMl6o6jZXUWyFQRnrDPU7QrTHV+kt+2i30d0AqUetiB0cOzE2o4
AI93Mx+VjOd9l1MWpI/rJqiHQ8xsgzSFq2Jw30VDx6vKxOuRGMe938/aE+vMlYh1
yxuOFIUoMnMsWC3Qd3gwS7OZtVaKs/2umyxZeBJHcM1PS5sk2JFwjhHRmDfQuV1f
Lv4xzpd+LDrsjZv9HwUODVU5Ss0PvREy2dKG/umshaK57czNR8BTlFhr9uuNdqoS
NdN1wye48fKOEtSxYRpGRBMNRp/oBb+k2QTR9yIfJtyyCuKFwOGbPB/Io+YxV4+w
Gfzry5W/rfOINWPLY3uzdCbzMRAfzkBrXoKn+MGLeJNwz13y3OOTnWQMg3weBW9i
4LpcuoqitiNl1oSZKonINzoJVUJ67f5BjEBlAuRw2Zk39OvPi3w4ydR4Y5WY70TG
JFaPCnzA0e2Mpmeg9Cag8a64VrfKfKBu3ChpAddXXXItGzRC7TCs2kaum8mbQ+qu
A7xjzgUJMHOtlTJnHOTsbYOmAy1oZUtIwVj5CVllX398yoV1P3098oTIb+X8tWFL
YLUBDTNNXkIigJm3x14tmTbgw292h1VR9ku9H9+Td9rCtwIMnoYEHHiD2w6fJ4Ku
OnYUwkz/NOKzngth7CW7SpJg1BDQcIBd1ZzkIv1wP5OGt4zIQrm65iCJvTBoOcB1
cvv1+fIcf46dbqb7NmZRUm3Wt7HarVOM96UxXockUCY2w4+V4VfFgyhK2X3nLN+Y
C9qvF19CvZKyoVfa7ot2ra18Cny1zYGYNyFiW0ikMBYX4iQp3o71nPral3g6O050
s6m6E93a4DuYRZwT9ozQ2bjdgFxUShhGS+wuPbCZQbj7aynkmyQ1oAytx+7LJfb7
ucanPvzA0ZFIa5wL4IKJz0AgyXVN4X48xkyiDSvrvWAMl6h9HUH+Ma2IgzbBSQMd
SK75Y1DsJIn5SFiJaab69x9sG8qNEv09fnmHxwHlFV+avlJRlybYypmfAGLJ4oc1
TE3v9Y1K5ZBaDWkUeluzA36nQ7D/G2wprpxwt+wGbHHWtaWRfwu8QCySWuSyKECJ
kkPyi9crStzKcDypI1aO/knRoAGLOKv4O8yWrUhQJKzMIelsGZ2xrCXoApvqCNpA
nXWrDFH4Duwic/wyZkpgncMgkt1sX9ZXbcL9qiQAOyf7Qu6D2KGQg9gtaeJ1f8MW
GR+1FQOvXMsQpvaYjBVc27StGCFm29zXkynCV9zfn+EZbygtmkBNQWzwXk+V/PkC
VEiRBMSQL4UbyGSfVua0QundEE3vG7qJ5NW0+k3OqrjhGaM+fOG9s6TGjGK3nrk2
grkLxXijQG1CbO/Y9TooMmsESdrul1oXLmZXS+bECpmzJuj+L04i/iewkhw2GdeD
sZZot7TcwSh8TsisvLocBr6ubxzGfC2lYPJt3Qhi5mAW6l6Ez/Mh/2iJryo6+6+N
eqE7P0oZ3mG4NRRBeKgqfwOiKVoKYekdpJUfHrUqA3UR1l58r00QVMLCV1HpKeK8
zZQCPzBCBq3q97qjQsrRkgF1Pzj2GEjEOiQOqal2N2pOpR3rBBED5gTRFQJWaFpE
RUxd5NAkYg7GyOxHf3ceSHHtXWaEW26VSmCz79gW+aV6fKpR+k018zrDikaodLjs
Ce2ckm/jVHi1QhcLwgXMiCAUmo7Yi9fOxHovx3QmsyhuodVSaTttLxyNRcsmTOmL
A81CD3ppC7jC7oi6rh5sjlIT4mgSKeIjduKLA1XaMlb9xqrWfW3qyYtYl7ARlLzD
j7W9/6lA4kC14npBSWmqaFjwbMTsIVqS92x/4OqRixoj6+s+eYbvnUOOMh8k1j8h
zqpRDT3IDcA32JxNAswMlwEgq5hCj7bPDbGZcy34h2p3ZwZNP8/vO3USCPj2QqCz
0hYHT5yVpdQ83afBde96ynjZZ8PhyIvUr4OJQaT1G2ydJ+WpmTm/ft98jxExTr5E
HqL0AZHnk6XR7M+vo3horhtMe0KtvCvNb6kPUhHU7EUlWs1kNiqa/bqDSnqBUbwK
yO08GKLcpk6ghTIeN160rC1257yVV2JVN6mSXEJEqFk=
`protect END_PROTECTED
