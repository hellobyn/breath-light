`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpjtBkzKW4hxsFM5wg1aVbUy2DtbA6l0IP+IzNQFP0xcloGMJyJ8cyNEfygfoA4g
e71+/FdIPDH2Wr+DgpXXbuOq54mN7eF6cYmsDzGXzYPNcp4WMdXEi6icYY+OSIY4
C3HlhZDnCva6E7e1gqaH+kK+wivyTs7Kf5erE8RXCgOyIxtTU2enTQJn2RSV7sF6
P2jijY5fFkEq5BH9/4BBQ6Cy1Do3lwVxxJhTY7UIeUAPdWEbELxYmrFKfStwjuwl
lt1cxkTqegELIw+eerS3an/LAoEN+cLwhlR0weodrYdTnpyQEnD2q5w2C3NY5C4Q
6jJE8zazB6F0yr+8RdVh/HcuAEilXcJD/GQXOsP1++4zvsn/WufoJTPfbximhhI/
LZg7W51bpGowkw5ntZF29lYBYXvLBiZE+vGXoRzHTijqclhAbDDGgBhzYJGnyEr6
AIWDG9J9/R4vexVLj2XDfC5tJ2xRH4M6m1iWHd04pMQwGuB/f1XcdgXCRTN4rFrn
ekyzG1MSJc/1N4iiObJS1yVvBIFurwgLA6hbXWzdb23qOYkLl+o2ZGxQ9asERCbH
ooHc4hCIi3t8kRnljScTITBM4GwQeO4cIoOr+L6MXZ0lXwayaMLK5XUS53G1qIuV
dE56DOBU+iubxdiwrvfClBs+em8ecqIT8eXrY3Jsu9Q6FCJp+FrDKufZRg/TbjME
P9hZEC8+vGKod/lLS2fafmt9tOCkhbAIxH1Z1WfSLvrCA1bfPTZTA7oz7DuNrSlA
UsKPeRx8YEzKvAxhnL/7xg7gzNAQa1hZmUz5oJeOSieEQgEUkERnxAj3vixP7BJc
jSmbWdjB7PVV4fRkRjVtEcIWZkzL+Xm4K2N4NbSmp58uFNI02YrRJnaGay8629oe
rgk5Eo03GG4OqUaZ0VINGubn25D6REhG0Ibd3ep65um0V4yBWXgLYB6b204irYcZ
eMXp4vQntGqRJzCtJ1gY5MTZaoKTFYNd7pK218W2r5nKhITf6phrJ+WG3ESfhy/N
K+GRVrR+6u2WmXRdZO/aH6yRUbg3MaPE/m3nROKc4VZ2Ng6oWavcwdX6qCZIULWt
ZKjHY8WO00ZHS+mv/28KzwHjNB9chkXC7yPt67E8lIEHFqfNCPZqfV/hAu5aeiRj
tprzCMOVf9VMDOoub/3k27Lk14yCYqUbqe8pQex5xRZb3+N0jwe7IgsaodlHBtjD
EMhoeDqRTS+RPA6TOhgORzVXPM1G3WcfGZi9r3vkUoygWFoRLkFi95dJu4qFf7O7
r0oBi75mBke88NZ6OWwfthrk/98H/0yQTDfshxJiJFnuAjP4wnsZKVEkd77T7cq+
JmSNAHtALrxOtdndt2NxwtERjhNM2WACcAvBgt6sGQaRsSN1le16npEuD1qwY3Z7
9aBOTslYdRloj1mbDj5VeUhFek2kbw9LzkUhFypYFJzWznaxTt4l41jfJpoXtMFE
31SSo7r4u7qc6Jj9XcV0IIyWq366nMvD4MZKcnyGADqIYlD0wWq9i6kMk6yX/Rjw
1UKg2k6QzQ9PCElVzVRInSoaA2Wmyq8cts3K5c7BiOrtZfPgO0OZ5sXPiG3+1v+i
/R2bOlDValZQcOnB4loI1BZxcY8mmiQDmWB8uJf2CGHkUHf0zKl0T2jV9oU8t5C8
TFeEkqNqGi8xhBxmxsrO+PWIfNs5Ys6DkZb2cySIpWX3FZ7tpDs1wXS+CoJ85ZRq
R+Vdtfn3NFBmAlv/AWOozEm7tygUqJw2SFuKcCoC9l9FyDRmWuE1XLdNwxv0m0PX
KoHSBsq14ZkdrbCovyFK8DZ/jywEU31B2e79skRmEfylzZ5DENWtzlO0/3fDM91t
Hti0iTiPCgFMxvEbrlN7uRYYP40ICD02BkBOTQjRkPUjDU18o1yOh9HG80in+RBe
xZqXMQfNmr3i2+pj4n44uV0uHfNbtSRHZXs6QPz2TNdk/PjNkyJlnxd8iroQK4CJ
kiRpRplRlm5+IKJbCDRyTX2P5HGNSa8OxdA8QmmLBif9hzKOkZ/hB97arG/Xv+YT
ECMUoQMS7IjUowCysHWJlzTEu4hwV+m0yXz3kmr95bv3x/VZLFvLkWoqWrkJTPLY
IPgFNNV4+6pYBJwcTuBxl6iDM82NhYLhL7E+kqxtbWBxxM+RwfWWtGhZbCJ0jVdD
bOlYWlpnclGCse4e9Hd4P+c7r0nIAf9ydADfUrm7jizY6UPU6pTctsALa+C4mqhc
Xw63xIce7u5+LASpt2r+bP72zcG1AB56m6i6d9/axOjAKfMzXlxNlYssHVi8ej5P
naJPN9xggoQihJKCNV1mPCKzOODdSR+zvc7oUU/E+weG2efWCqwhxg+zMzn1r+oM
gqjyj7WhBfazfZMnjITjuhyU1uzVFe3ejV82wRXWpIMswoif+SIAAcI48XsgHG1j
X7W8BXilyIsgUnATUxWgEoJqm0PClSzEfTaW8VaeGp2b/cRWYvUI3rleDAxYn5UJ
elY5KaaR/WnXE5u4l+tWoEwKP0OIByzhQQl5r75gfbljb8lm6Wbs29H0uA9Uzn05
iTR4IddF2WodLbdIy7HQd6fM91MnOvcw2MUAAibTCjHRu9hkoMkWWKH1LzguV+/d
28hcKYAnyoztePMnaKlKCBBWuuA/Zs9GHwtbwvM+GIppuRQ8l2L+h4NO7ZlyqzeU
sxCn/tgmIO7//7Q4FbPtyRBuuHkhuhyoyDpn4YOrQFWjZ/7ggtciDNT8ql//3X0m
jIwT/MHlThwIaO/CkdVXaDKte+5gULLLNZe7wSa5Tpajh2MQCaBvCi7YnYPagY0f
ype2uClD0MyeOpVLvOKjCBlMCMzcx2LiFCXW9SazLm9dGCELIw1qO1akBFPzUabD
EbWezxjrKj/hi3XsnBuY0wDBn0jkTjGsNJ+GJDw64nSXkYhK9ycTpCtk7UhPjyiF
KorwM9xNjYJ/vAo4mNE6S+5okv/tYEGuW6ETmkqcTsh3gLB3+/LdjD7lBBXr3BpP
yu7PX2GXSk03GA1hWIVOmO+IqvtBvNsQBOS4m6arhOv3dzSMOIeaVAwHsMaZVtyU
FZ8exck7H8ezte2kSfuDWe+7P7tG4h7O8jQxTf0z6q69dRBaFToJiY4NsqTAlboG
+VEVkymOOijdikeBP21KN+JWj9ue2ZodAg3STIGfd7lAr+dUb+hjwIiWoUkcCl0B
y5FZHwrydVSADZiFpi8WipJ0N0fpPES8O0aYdgZ5SMrz7pmcSztizZeLuG3AwkgT
v7ItsHLQ+krgq2TE37olxxZPgSMeyhPilmet9iso20a7IjxUK4nOAgJZFJdgVt4T
GK5VafnyIKhx4yt3hmJS2uHTnJsdq1TBo8K6vSSGQ6odzZs53FUxEbQi0pbtQYs8
kflmMvmwCETkl7s2qntN4CjMcZh39B2CluCc55/f0QMWp3WjYn4EcrhoHhIqLgX1
LASGdBl43rS7hi5PKWoOnAQd3+1kD+8A2cnsCG4zfW3oPtJ0PB9SiK7RiTNbTqi0
Bn576QUW1VEZTUmpQ3xdhYD2azrNM/oXKuTSIzvBK99YqdfzrT9qRRjcNHV2dLMx
2DjP7+sxtphcA6hiPYn5d2ES3byiGL2bh5E+XPQDHHvPQs7COAXoBOD2QlriKp/4
DJM70w4QXHvfeyi0qdW4gTANyw4EHKlgiYu5C+GGaqdZedKnaaaTfuXlLikTUTWa
WAw9wsrp40LmRfQzlk7cbl53iznMv2gRAON3PRLJ4n7tN/HZ/OEaZjTI2hxweWrK
UZ45CfGwxvw6XMtqWR0BovbvZMwuJgjTHZvxi3ob2ctTv7kOQXHjeh0bNc62HJuA
nWJenXDc+zOKiKBYevT1zfSjEBIFW7TFOkD/bpHh5T8a9jywLbZmsxFA43BwpqmB
CR2JrQiAcnyvqnd04J+0aPpalgEqhp0PK+U7ncizJYRCIIUrkGDOCSrKZ7BNejT9
oTocfS/r0eGNU3HT5Qz9ed1hnjpIhXlBBXKUH7lmpZEC/CTIy4c+kHM1YXxxgU/5
GKd2Crh8ZiCdkF2X9tjc+VG17lUhk3RXKnhzkOvFc2KBkVMWHLs4k5TqRb39Mcsx
`protect END_PROTECTED
