`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwxwFqbHo3Ko7DtQt/GJgVEWJarKgRQlzHi3LX80tmAKoZxTxpybto6LUK9eKp9Z
TLVKHH7Dnlnf7dn/zRa3MtYEZTpSh8mCVLxD9pyjPMyE7G6WsIw8HJMuBgdK6U0z
OX1wX9xKus2U+4aXPIZnLToIYaPq5mPFEdd9Qn6merZLNBw5MA6kTb3GXZRxnTSl
o86V2sWh4YxNSl11XllurdZMFaTaeOHBaLi26OmKfN2U3/Yj2DXkXcRW0bafb+Oa
4mCIyyb6KykpioVX9d+l5YtX9+RvIAEIkVTHIxQjjttXsv53KCzHMTXTBjNPCtUZ
Pqoy8ho2nqIbUcb3z33aK+obcfGZq7AAYyMWC6n95lrX3gqlL8IwenrXYLKfai46
fdvPO1JY4OWRpgCVCqnOLXg8YsiOCPPjcsHKgTuTzlNJiy+l57TmxEzCZpvE+RS/
QWq9MP33XKOU7BnxZts0nXjUdDBzaiyufepV/OEX+lzC4JBPpWIqqtXVkHIIAlQs
Bz6KiK2QmipJ5eBgczP92EKLkdTNeVuQKwmhrm28A3MkYknhQwOjuYEVy7m233V6
6Rf6m3bNiRk5XZWLTsePCPSfTuO9eJjjTMQ2UQWpnj13TXNj7dtpXAwls37KXdxc
uOSfXaZd9frCt+6PbASSGcZHlOzixEWNKueDWNfIo6qJUJRbAOr6ZPUXDij6KUDe
jFpepCQ8XZBgkBq3no3+1/zacwXwpVE1SoPB4S+pdtL8F6gX4UmqZvTt/m3r6Z3C
dQs6eZLYagsy5lwZrFPTKUoJMCJhoBnwFumckM3oJUKOtHfeGEL5APql32Jl4jLZ
MooDv3xqXeebXCCXaekmBrE8+RHw1nbqO52dt2mbOKD75xxyWmbeV0ZUOviC/1mY
BtKAhz2fm3RSBX8TQA10a7Y6QlmX7bMb9k+GhYyCJ8EJGu/TJ5ccucvE/gQzyvOW
+ejsd21busf6nFOmK1bwW1NzfPyK35jdilFzZG0xJZfeSx/+wCv8GZi2vry4Ahm0
HfAexSuK3N0um/JMixjQjM5+5ooj6X9aXrgA6U8Eez88ynNx/ZqQsD/hTBZIKela
UZB+atB05MtABOCKKkA+JCd2e5yoc/gqc36vB1i71ET2K2jrI+gGG4MUUy/qESs2
7ulnhZWf1Rf5+ECZw6jqe2ozymzZvWfzERoh0eXabQya7XXkJKXyRujUBrjdWGin
tpVA5DWy/wNCENReBAceCC/FEohU6l2SMBtNxMSWzHTrYOa+FKODzsRAatZEulIH
AMA05N28zT5e6Cv+tgqfBqeR+QM9jI47EXB7nWq8PWxKIw5ghvZ3ZhG8UYoZhWAm
mWlv3tmGQOy4N4gjSm2omL7LK3+51kcCzu49H+IiM9ubj97R7B3wqTUTumFB5d+Y
fw/5Cyf2n/z4IDJdz+v967PlgTQn/a6oklAaTH18jvOiZE3NfEwwc2kok8cJCS2c
hCGGj5r54Y22qavCeve4Sb4Xjeo2cVLkS01ClK4yF0iExSmV8rMs5T9KvXbD1t4d
8PKlm2GRca+GFv8+BtGbzVpYanvMmVLGGGJnkO3gQ3NNOq328nqOwZZ02MhKohkV
NdqLaGUN9qRPDC5UZDbrP8v6/aGQCggKv79vOilPDzzYxneTOYvn7OCxFoVjFAuJ
iJ5n93pEt7kd7mNEGL46XSVDCadchoPb3hn7z3lJK/ZOFuXAlDR2IVFjqZY3BFS6
0AXEu+bAK81PgM4/qhtPPVLd52V31vI69aZ/CDSD4+8PCBNjbYlMMrX9gjw2oESs
jmFlUEDeVdIl1Z/dJOyZApKpkm2nX03UNzst9WRXJFoYhsPqBRHLE2iTvTDprJzv
QTGXYpANq1FLE3mcZtyNbu2nCFQ8DDmbXyHxCr841w7tsQvwBvX0jAHC1fLSmcJm
Dwft93UQd6OwSRHalrHP9t+PwAzgaoKE0lNu3fnwP3874+R9xoHaJVnH6dRWjIa7
w4NNa5aCaVDXYZDztwh0Av4KjPtdOane9rN6uJn3+FFy/gdZK53Z/NSRUJ89z6iL
7iEJLJPz+QkXyPEJITnGrRMpGW3IugG+F3KEyq+zZykC0TTNE6vx79RHSvYnkAC0
0gukprcb0RdCl4OdFdhBwRQ/4F3jVtUqpgYWEE6b3gHXIM7NOLAzlw2n0Y/s3Q/+
IazsP4LAcSPpZ5G4Z4ODhr3fSbfjJrsk9eRiI0RFN1mtdjgXsiLWGwHSB1ETQqqq
LqTfazsxUvoydwWKF3O39KWHUgUDQtYHSauS1gSOJFKQniEht5lPDrKPTSQMuNiP
mbze3LZ2Zp9utUvmb3+AYI7KhIKUtHYaifrYnSeI89LXWtmM3Hz0zEqD1IANcLU+
EUVNCMAHjOAn0Oe7V57U4FYRsci8zQTR6amBFW3Y5NpomWzcT5nhS+yXDIXIh7PO
rogZ//9LRlfLnXK2aox+EFi59CTjoH18gLyQdP2lBOZPBseagB5sap/6aGtKgSQ2
IwOm2+yfp+3MGvxCElkguOzspf1oLckVcYho2fRGbTLQ44s2+0pxnp6C+Gy2AujR
Tiy2ECxwtczmoLhDUat+MTtRASutTIME8RUaw54nubzG4C8ijyxL7SUl+8sWuHy7
62IuT4G+urjfwcMizjXOxc53UGWynp5JVRYp40SufoWezd4GxZliKYRiroMXXfFH
NJN93oByucz0Hgi2+GGruTON5KIoqmgicJfEFOt8yHo6+5x+rOZjCRI09zzQcZe7
BmUICFize+vUVwdZipmbmYLRmgMfGWMTpjqiLrCgVG8r64EhzcARc/ElFV9Ot1pw
TI7LP87YA2StxfKmyTYcXo5813ovm99ru2llUJGwWygbc9Igv8wSIwiDWKJY6sYN
xULl/QlN7cpcOmoCNl/ZwZY2G42eA+BzRKm5gv37IepJ4VfNARXK4VUSgb+80jNR
LeW1RHRRJz3qsG7yVEaLtOO2Zb+bn05acYD67m626Hv3ilwFfE1NW3Y6d+nkfsMc
kj1y4KwDQMJBnzh3mO8y2s9ngCoRhbDnEG9gJFkqatBjXx1tsR+dlbqSovaUZOO5
upmPbPmBhMNG+7V8D0q5kiVBZk5iuIIEZNC9hI8QVg1nZxwUSP3DKXAKZ+z2JcpF
BfYP29U2vIHdg0mWEx8M5vXSg4oscZV6SIG7EqSzm/81ZZ+NCDjr6/egkBbxgLyg
/h/5to8Tyql4aG9hohnf6ib2l5IZ1AxM3FVx1DjtbDLJKPG53Fi6tY3lFAPo6GHh
tOsqjIvgCwaFxJASVVGfOSCp7QbfwQ9ojcmyxsI5ed/S3dVi5n4pJ+UAdqLLumAU
d/hjj/mN9TM/yRBeQFpw8dK6yhkO9sbdpX1zVMxdQWUhq/mpR4W75HrLLk6tP+9h
OVPz/jvJC9I7U6cAcV0IivxwWBbUy6aPvhLdkZkWQ7CxkVjTWJNGnhO1l87i4opj
ZhpqNrCDy2V2iWJSEMQbmQ8kyV2h6+h6ZbscbpVhdQ38jNcMpIMi400DVBvwLwvv
hiinZUZr+4o3BSp8nI1CZusqmjB8pFvbivqWeVyXA8U4rEYXsDoOUORAF0abk4NS
FNKmLxzRQoBSa/UTEdleDGtDZtSp0rCdqOK8Jnaw2F5oFOkm3o4FkUpiX61U5tEH
BXpkfI8NLCq9ZsBG7sSKo1c/wUtHts2304QV375vsalw5MMkHObjbxKw5wB/1lHg
ApQBtKr1wmfnZ3MYTPIxugTHtUgXbxwzokXCGmNUQVkzo61PIRWc4ilHi2vr0cd0
c6Dlil73T1UbaVopRNKqBBHKwVDi8SJEGEal1bt3QIqhtuO9FhcVpV4+LSAkDzg7
86iWeyTxSwLiXZC7+fu2dpwKviE/xqGkWVHdRDvRxCE5R+hdI/L1oHFVGxbHL2LK
5Q8cP0H1IC+Hc5uxj48hw6RCMivNE2d+sFHSCyuPDB4Qbnf3QlyR5dkykcyMj3Sw
aHPuY52u5PQ4prjW1OwFQ7a7648Q1o+VUJxiFfLzwqdCQnjDGa4CckwpjcOCPSLr
KcZwb9xd2koDEbPVy9Zg9DZuv1laNpuIqKJ9bSzWT3Ac6gaYMzyTjXFLX4yM679x
`protect END_PROTECTED
