`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwMJJprmoXobCN6rg3xhTG2DpLrESx0lcxVqFy72n+e9/Qd0lNzDmY4CdMmb3obc
YnlPtJpN2ZHdJ2dclm7pso+ymWwgPSOtBNyQx7QhAA30pHKp2I88fTlVcKalmFwm
Fzpn4LKhCiOJPcyt3qubUcq8hdIsDgYbjDAPBRrd2i0HRS0FDjuH+bevzAH1e8g3
EX8rr81zeuaFMUEvq39Th9M1ZzDm+QK/gIhUnsfS3d5BmoeASpUM7EssmZ3ZfO09
NXXBqT+FRoJVNa5cAgVkLK3MVMurIkLg3iHBacgFbGpNhXlzYVLBX8kgP/LYuwaI
AhX3OXAdup4zwRzirtGTsWPYIJ5Z82cfdJw+4pMGchU50adfmGRlIsNoAPV8RiA7
OT/GENxCMMU6JnV9nkQzM0G9j09KTVGLD/aRYrNQC3SrwYPvZddjSucLNEKCDNp7
nK6Qh2l0MvadpN8qCtAANoSXaj6aYxUQqd8C1tcmPOj3oXCetI9LpmM4W7Gj5uMF
4jWQ0FcdBb21luekYv1qGDy467v/bQRqvqcs8U1CmWFSc8UtzNBxilPC75gwrxNP
JS5YTEb7QiqAYQMv0xA6CRFRypZ+oYnXVj6H5hMmp5qB2pIGxs6x5dIxXdt0zxJ6
/FJWuq2u97AAaxrYdRSGTwAX4meJ+YIGAllkMWR59gs=
`protect END_PROTECTED
