`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cPOgsGpJf/fI35gVM72H7Zh2JvRDy1K0BoPD26Vmq6UN5cvYwmXyFVVNy0meu9j
96Zb4ETlR8WjoTp7BDblR7TsiWkqp2mLFT1TwY/I04mjWHOqaf2e/RHk2ncZGrnN
Xkjaba4BsvysQ5KsfGIC2F/EsnYIsAJkKXLE+UGskiCpqV39E1O9Fl6P+Q1r8AUx
EVRcaJM60BuIMPJDZPUplayhh1cnGsQsBx6xVOhJMCB65nH74Rn1WwTw5Z/rpTqt
8bqaSqb7tK/xbyDnKDoRTbLh3SHAu9m9RdczhCK+bD+itwro0d4/O6PErzO0Ws4M
rxWBIXLoezjLaSiLULpxEhoezsmTyJMkyibNJep+7zJ5Ngt9oHeiN3L+/UrXkZ1+
JGsWVRNX4pqgoz4au7Kmwv5reLD61ij2EIz5EmlIwPGlYyJ0NyOAmoU0PsuoQS1V
Cr9a9u5GcR7/Gu7B/RWUBMaF86pzhZpbuV+dLq409saJlwSoJO6ND1sfgk+K2LM2
BMgUKMt8DhivQdrx/bcn6Z4ro7h6OdtNZGhSlcJDQ7/QrZzxjIbFAfy/esJ6e+q7
on7h4FZWvw5Mscod0MpPdQ==
`protect END_PROTECTED
