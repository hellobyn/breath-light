`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xW/C9twMYn9tvqVQaE++ihzpUO5kUaKuB8rAvN4LGHncZOUdqQsZRo/EYUivUVZh
Lnc0V19Gv0b8b3b+nHR4EAJI/1fgYw2w2q/oGInDs6bsERUjgK9ZAta5LrhziVEH
+DzjvSk6cm0Id6GazLBXnN9hnRcYF06rpvX/gJNP7awWk5mpHE/p2zSgXQc5ObEM
yYphl7CR4YZJ+9GfTVRJaDZ5Ie6zOQ4zZD1HC+qeus8frA5tWlQZ0WGn3gt/yHrr
Pub3djLWySE/iidvpUaUb18gKRq1bok2JDe/PKvNlj5CCdvcbOVyB9VoYIl6v0dk
ILJrWQlmlNy3oSZoXb6av/13YQDNyeHgflK+mU8AXyaOO1hcDwv0FLq+rWyPRNed
l9PpOPFpxgZTlQbzT9DjWtsC8IaSuTPJR/d2zLjajoX7kYrKdWot5CWc9usndSY7
VEvbC4k+FqofGhVyuCh9Qfzfk8aQI1qPRwlQvPEcNGoRKb+4Q/Cwsd+AOgo/TVv3
uQ3CJAXR+AvwmTZ15cW5JtZCRudbkRGzzjpG0VKSrsujbssNeHA8CREm8wimo1U0
bCXYOOqLoQv/AeEIOwnO9itxSxlal4CaJ1WQweIcxJIBVNWAEpOr3sbv3ZpKXZok
QptKiy34j36Z/OVJr151we6tjT+KhBSCA7/huunEmIeZkTlzTpfkqwDTZequuXTt
CK/vxn01elPWyaPFRDUcoblCX1DrztHpB85iizvA89JhzpEK8AzhyrpDcI8ndwxq
ssxupDJqABeoQkmCLN10SXm02ZkoQlPFQmeJ5DdjpcfB385DPNP6h0lUi182D7Vs
/lxr8v2FjJWtAx6anbRWIw1kbpql/2+hE86TWNIrl6607vVKFXRU3TUbijfBWE/B
P3USFFgmPziJoW0DDqyMZHRyFmWr8pKNOnMBkFmO7LbaEhs+dOlQtVt+vIAPTF2a
70oXUQg8mqYkEi+fpj6t3Cy+zkC5JP8ETsV6qmXq2okWxdzBwhzUruA+zYhfsPYO
2paNHHaTbOhZryHu7zdFwxBzNlSzzcj3bZhdopEExYFGaUXJj6q4UCNzi/hrn6tm
TBwmXFHjsA/YCm+DC9+P9jf+TzqDHxhfoxsABZnhZs//Dehzua792vzL5adL77Ay
zuOn6XAkKVoE6TlxDruIu5aVA3Xi/GzyzfUmidp7cR9auNaT0WAiJ3gPmeag5Rin
gEyy1ki+aG+iUtbKlErrMjsO1m27i8ctmfcoCoLBui73WrpxqEQVwR18LjjDBqlZ
7gHwGD/nDhxrvPBiS4HXySpufmhL3H4ZqNbyHnHWd3qJCgre2ukbpte1rbPRVwue
zOULbRbRNHjrdmL56Mu2nCejky2ba6grYik/qOJ7X6X2X9McFWPSb4xUAbo47K9X
BzxgMi0DdZHc+Ei4pSvLweKg3i1Y2O7fURmuWrFIp9g0fhuE1GO5hWejobE1jPba
L0rUcleKyjpSrVmkB5n2tMI0ieLGS8MghYKeIloKxF5TNbfmfDMnE82RbiCZlJOF
cyqUDzfBshwIUK+Adic8IP7W20e6Mu8MiFqDenwM0ucS7JNi/IoigcqiCgzxJj2/
/1T4FykeezUy+PpEEAlywQ7bT0gxFxvECkQagmrVHT09h8ar754BAkYkglj7Hj/z
AeeB0ChKc/GXl3l4abQBttWrJLLw7cmVYowfQKisEB1FSitUJdzGxTcvzXAlkeEN
eB5u0yS/4PDCDfLZuS3U9qNszx/8I9+5NWaSHAJl7VgKJQ+hEKcpwuLaBPGhbHvy
MV13t/ahRXMEyleI4CeGXi/SUhoDHzABAWh2f/si0Kv9PltdXAc6J1E4sxGmeXUT
jWpGxyN7gLLcTyhj5RPIgyoa/ad/jKTbz2IOG5lUqsv1qpSbDhbLAo1t7LU/bcnI
kJMJRhYwBQ9xyig5hRoXpRwwlQ4duWS7Q0VN12eQvr149WbswaKW0KBumpst2jhq
qRXIzzxSlbnCe6SfU61j3Tiu99qcMWYkpUL8A6Qza+//sr1ahEWKyYiWJJBG3bI7
OAuUWO9G3aeDDIE6euGMbVqJZRqfPULYJ6auCjqsCtR3ewcvXJqzoP91b9+XhB8X
+0xoADUzpdO1Ere54nhxS9/3nseAQZNXRzJpugD+YJNE4enFQt7XqjnxcbZ4xr2/
yiM2kf/K0+++8z2xKimJS9OJu91HWPaO8U+lfz5WFNyi3wTfOEQDOYmNpbpdvtpS
i1H2+2uy6D+/6yUNPZ8fh5foNSzQMugLi4FpKpsO8Dkn6mRYespv9tlIZu3ohakz
Mahh9ZimhbwuaC7pL1EstN6Fe5g9MLUOWffCCt+BNSliW9OmVJDvin5dhZu1nufp
jtECCbiDisIZ9SVCgIrX4gt6YCr6efr2JfdheNDHkYXYB4X2v3Z7E7MgLnQ6mbFJ
LVh8ybBzioOAsBVfGWk68pOq/Jv+StTgq0xnJEQnNuLwcqNuVKtl/gJqAO4TCXEK
dzV2vsn+neFtcE+0SsO1BuQosuO3HyVrR5vA+19waRGD89qvm7jWpQa8Rh2mSpbH
hjC9IA3hGzYVxmeHxi5CkMsl0kev89bJt8I+azofcg45myRgUiD7lcbRSVuX8WIk
lGODss+it/cuS26xIHy9WeDiMEt7nblS0Hp94l4kw9EaWK3q8Kw3yfXtqY4q5yz7
B1Sy3fFRlcIhD/TLSpE0QDmBfQ92dkAoWPvngdSbhtCvMizLjktdIqR7BeRJZaYE
uQ2UI/z3pDMwItuCmTyjLfI7l3DH5oaZEwmeskv1bTuLP1dndPmGjlbvjtIy3tSS
N4F9bVaDLqSRNpbIZwrV/GeNpW2GOANrz5OBBpmy3Tq1ttCtOg26DV0nqqC7e9H5
7Hj0qsfkAi1d9X3CHLXpw3YvJmVGAyh3V6zHaNgXbALMKcIefm5JXtjqAmQFweMg
/WNW9UORaaubmyQRd9+o6Ydh/vlTOjAMIEPpK58RHcBedKxpdleo8Tf6/KtI7gpZ
0A1VpIKYrg9blRZp5DHz4HeCDAZMuQOgR6SAF5Yoba9y5xDFAp/wHluH74zubZvq
SjRVgIQOTaK3C9CHZONhBgI/vNn6HTH5KE20CUun8U8cAWidVC6fRiXBFXcNiqFK
fQmStZIBVZ93Iu3HnyLLwvlNAGVTU6zhZ1+4DEazvA7/pUFK2+2hOcoHJ5mP0L+i
vC/ET8hwAGXxVA5Lt/KYprOZ7NC/hSP2CRl7S46ER2mY8Fw20b41h4dGQ7YEg5H8
ADsNzwR6dfw+p5I8WPRswzNDyvWH2SGUXmO4a0zQnhCFQzPF6rIerSRVIgrgOb4C
AZK0aZFBbuPlsDmrh40XGIIQndnlfEbs6Ecbfj4/x1j5A/v8P2ZymsyQ6CMhxKii
nbznGRg2u0x+1C5QoCxbopOTFHQLHseRB0RGLfPc9QpdjqDqjPThJt97IGMQy517
p6lStPKr2k4KIpPe06dECELL0KIbPlCIdwCNUz+HXfXUfNSa2a0fYvcSdjpJnSuL
+++hs7FlRkkWer9XROAQuxIKG5m3Z9rB4JZZAOMV+f6/S2WdDYdECh5I0RKYOo/Q
hSkc8PYOLhxZhwrmr3zREtXy6ad8EFgDXnK0PsqPt2+ZQ0ysEgKa8OazFmzGo6qm
oUZE/o//p9flzSKO1GDaVZxgELTxhBh9wBffHkaaJvQDmU2IOaBNEuLYLW+GRkmM
S2x0GP4QjgqHYrjmOeXwDYduKDQxqENoGRPIGx+J3zYjwI9ZrbeE/vmLnDkLC0Yp
vsYQHpvW5buDWg8zdpD8bJXDHEKTxSyfk1mPQVt3evtv5Seo26+2pEvFfVRGVxjO
LkQbE66T1NnE6cJ6gDrKa9F7GCGAmMUPqkqAXNMzELEzHsn4/E3mpHudUWDuiHjz
m55FmuQvglbGhlLAszu6+WesApYAAFAUhcuuJSdBr4ohOZHw9She8H/boJt8Wdxn
l8NAbDX6t+QAndHUTj82Nh3WXLNAtviYGAHYEeoeCZ1XX7f8MpjyeQgN2Pf3XMvL
EDAhwigW7xxhIIrISadEuQ6NKWWWnMgTexIme6SVOOrwIMNVRc1uB7qwZxnXWror
fZWxTHdRufWada40zoM2oQzrQepu0Ly3WPh0JJQAXiaaYEgmIF6JbwrDC3rr8oNU
u5/e3GsmiQZ7zQyxHUW38tBiKlinpFp8Z7kzaU+4SsdaSODGMKEvaId2rhhBh9Tl
ms/g+vIwVq+2+EFIGszp6tE19WhCCedd1df5w/apIf+FTuDWGPLOR+zHAY2G+J+W
hB0bvih4SfP+mlZGsiHv2GDMsT1WW7ie4wcT92Zx7CpR/jBqKlC/LeKBDRRJG8vG
2oNdkfYjjAyJo1ncoUrIIjNI98fYG79WBAUJrHD/tlE=
`protect END_PROTECTED
