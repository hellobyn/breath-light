`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHfkgFrf3o0kMcXvGjA63IIK/8nNGp3F/q4/AlN8gQYkPt1bqfenBqOJt05I9Cq5
GHaxOHSaE8x7wN0e/y6T5vrN44NEXmiR7Mag0CPJJdA8prxKWx8n85aa8nfPNixb
6rYu5DKxXQlfqJ84WNDaL99xT2VoCqHF7s1FRZpgKxLpTf9YJiBFB3fIyz7QnddF
gkepHCcOP/wajjv6G/aOXo3rqF3FnWCs8JbJQIhU4n5+BD+qDfJkQY6Vcba8MYx3
TutEKwCoAlfH2R43myy3Yd2UPajfo/JIHRVP3T70yxUggRJK9qqVb94gbXtSor89
yrf8nEtzQCPuOcHe5lXcQrbHYDqA5vMRuHKgK0nt/EH8pdwT2CcWTZfJWmFM/xBi
y2t+N4kAmDAhx1+eDi6mnZLM7yPIWCsb03HEpIOb4gxxqomxSUo+iMhb1W9s3hHn
S14tWAgMUNaUNGhnLFpvC+zWL8YNscYsbCQclzAG62WwHSYqnkKbHBuMuR5Gig9U
3cuJuwuN9yqYL67AxKpOBMMIpzNUHJDS6XS8zwKEyb8Sgj01GeFYwgxe2WEseFga
MJkt0XXlZE5jxqrarnZXtn8e8cKc4Uih71Evkq3Eq97gANtE0OScThiJ0wYg/N1E
RtyeH1cn6lZvWklysTDmWIagu90CVldC3J7DQYfkBIhMBRmRa0IaMIQ+PGpUhzF7
CVSsYpWMy0juS9q8Wl5mJVcv7QfZ61u9ZH2+qYFuDkc=
`protect END_PROTECTED
