`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mySnnA+EZg3yYs6zpqRSklG/4ThxeIPr2Cch7b8mYwP2G9Qak4QZ0HS0KDwwlzzw
vk8xjV51i6iVn6TlIyX2I32p+caT/+MdkUQ1fJpv/Jcm0eAVYKh/wGFvySlOGx/Y
wFFDJTi+MjvryeIV802VGXhbI3mjNJX9EGmHWR9NpE3X/AXfkSxok1Khw+nz4YVO
s/iP4ofS05LOpih0F/RIUF5WefrSLwAypBubyWQtOM6APTSDgCn0JXJYZblJTNFP
azlwbg4oC0/hrxa+o8QkBn7QFh2IbP8RE4B0gHHCJ1z4EOHS2PumbwqCckMkhe4F
xo1c6Os1JnUsv1Q9D7AtY1Zg1w7e//YOhbOvXGI9OXuskjv4NpEeTZPBjOqzKg6s
x01FdkQcXCiFzDWUDTpxu0EfQ5FnSVKp41I3goI1g6Urv1SfSlwP6kAI6iJbn5V7
Tb5ZyAiT8lSxaWTtWi+Fj+HZrZGqNYkwn1h0my9qIJe3pAk3k1BhjTsf06a8EZ0M
EuH0Jp+gKMEkj/3efLzazM38O5H+fWFETQhz5fV1XMvl9frAX6m5izqLq4oSOp2G
Jbv7TC0AwPNs8/Gtzz+U2yJCi3bEkDBHf525JPKWxrJKdrDOnFGUwGWwCAIH+X8E
tC8h37aIdzIORg723Y+XGMAMU9jGxSgD600+Xz0y41AYPrIcnNQXqiMNZIxumpgK
e8F/krt0SC4wXRD8JUO+7WdKzqMhIeRpiZqqGMLw9OJxQOvrnk+QbJq9WT4/22bS
0hROJ+GC8o56p533g8fNSVfaBJN7AtdHuvratflx2twjIodloTUV6oGieKjpYVRt
TeEGOaCF7c3leWl5JhDjrFQ01WE2IVoBw9CbQAgouMckhBCGlyn8MrXElQBVeMWT
pTovFvNIPboq/UtTqfQrElvkWMBCfyGQk1NNwJSxrDz1uxWU47qMcLkVz9JVEUra
tVItFS5LTseEDLHBMbz3E8NuyIDnpDqpdPssqUN1Rzi4sD/9lDi5EJndgY3Ct7Uj
lN56as/WeulaXGuPqFncKAkAdQ+fw4ua1/wMbfDCBsCVJcQtO85v/1uwPvT2iHAn
0VS3Bc0kfRpPCh1ek25r/f9VeXG8VoeQ3ZScSSCFuSNlrEKaQ3q9IwrwD5/UsHxn
U7fIjR8lItgfqWfTuEkxCXQF4Sks47VCnGaDHJnY8I7WPtzZwODRePa1g0oTL8DM
X0oZzfcGll5cFT40un3VLncQ9m3S/5ZSQeHNIPYNFWpKyDSpD3ikVWpOfttb3Yyk
XNfbYSMlfri/xEV2sBRwgtknvOALlOfevVANkxBHvUoUcNjgH+pTU9/sHOuvE1PO
RUtn7/PAv96PM29vkYo6wqKjMI/Gca7ker1f/Cq7wEbAN7LCI1v0H7+rcPfl4IV4
+8GMI66BbR4U8qsKLMJ93gJzAVVCQXXA/S8ZMGKhmj62xJcZeIDaCRetXolfQedC
y5tKbCt9foivuYqAljFj9hEFxElmGm8AmMFKrqKrfRM16tLd9SQ0lQxZngfEwi3X
e/lbhWhD2UAxGthxD3hsCqta7J9+z9zFt60Yj4OjROh/cfxbuTQzUUfUwpgxpH9O
`protect END_PROTECTED
