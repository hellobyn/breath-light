`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDuQ57/wL837XZ1w6JzwkyWI8RLjOr+jQHb1hfAZj6a0/9GVhFyYdayS7WIBvzsQ
XucWV8WRdCf2basL7rZ/18tSA1My4ddczl7vnvOf83k6yWr85Y92ds6iRInnnwKo
hAocawrh9Wk6GFYledBVUqXYBuEc4+QTsa9FBSHI9yPFYEvmXZAz6gNzWhZ7UTYI
j9Zr6Wb/lBUNl71UUzF2YeTXApMS5scNMdHhlw3ca0UdbTzj9jX4jhDZKCDBPpNz
pGt08gScKywnn3yfLn0/M8LhDxd2deHqN719ztjjxZpByY2y0iaU9tpOYCUMrVAS
DqCiBVtbE1Tfkre82hque8yB+k/8UN9vdfVbNeT1pLEoUGAgxVi18fUHNN82vqTS
Fr/EpWDSlVHLB/COuuHDyrp8dKtwZV7vCr1D0f7ffluIomuLiFBjXJOMTP5uWCzJ
v3FrZaeurh7gsxoSZExWbD4MYZ9DiR0K3RGTfO8p2+LiOckLuAouTStCbfkEvzij
gaOi3DiNoYjyLIkJuAdUyifBR5O7qio6j1y8X9RWI2XiUJUnilov+95OuDF66LEj
3//+pEgdrqrGu73/F31Cnc9heZJC9gqJgN+pLY6OoRXuwJowz5kOTzXUBN0ezC/Y
`protect END_PROTECTED
