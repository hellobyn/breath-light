`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QF+HAZy1o/9JutvuT3q168572w8CtBd2EdhXV0R2e9M1I1GtYcBHD6XTqS+R0wuC
jpa75mY89FUX7/AdbuTl990QSB1BVsesMBNrCeVpUiAEh1xXH7yZx7oMzTalULzM
7qV7GpskQKJobIuWB5fKPdvh/8wC+IUJlGRkinYVrKY7pbC1A6T78hYO59gJmbER
cqrMvYDbWOOABQkk+ClDF77Y3BSeY3TQGrkRepa+pr4TPWhzR7pXOsUGD3SomWb6
JYHHe28yopXG3j+aZdKTpmlG1MAthBU32zPLHsLNLm9/TD7n3LhASm86vWqejTl2
oHScKPmdtYLsL0r6/iQXP3QaaXmHOjTnBkfrMeLpPLaCVYfj/jnsqCjyiLgwpZhF
crVXSExJ9cs45j5oA6nDc2RzzRx1wZfAHUzeUxZqR0YHBdY98MPP3K63UdMCgNb1
dhwpEUTA+uE7VzmMkDp4IokHcpWoLEES860pY/t2aL/rTwRKx/iyPYo2GeoRTkPE
wfOtDMbmhA6PS4peFIzB0WEfam7P9ZhcQ9eFJAWo1XqseviK19XXLEqD2l3yNSCy
1fejoX8lUzJLKYHCqOvTSpBc5LKnK+1muYXCnZ20MXB/8u5BlnoZ+38ACr8cGS30
2flOPIV4yVYqChI0+zjUTIA9U7NNybmNz1O8nvHGqtWKVaIJVHPuWC2PxsM7bekb
GYWaeJvA7Kszx9QBcKHymVIl4Z8Nlc+sPwZbo00sSC750JZZHi6Qu8W0Ne/AkGVb
Ypb6qYb+olzyRCf+J6wTVvUjtnA+3roZu7F4OMP4jH0YrgifoCAeZwuOMXtq21hK
d5F0/LRYpxA8WvvBu7eXD8DynaTrZdvdMcebYAFjmQcLVbC+EvjVgrLSf7f88nX3
hvLfKmoDOieJwq3ssdSU7r0zn66wwpWd59RRyp50gPBTFyyfXLS+klmL3rpIttYi
FehxsHr2RG4e3JqHdzpxjMQnBb0OUhhJYoWP5lUYLCyQvG9lJxPOoopSUpXtSfkI
a40EUl0Eid3+axM5nMT5v2SSqUxMR0nvaIxlW+LLztTximPJNb9KDF/tk7UVu3Lq
E1AIGCmOXEOLaT1Iz9v2JGGbXf1S//F17UQ+mAgphEGbVDzRO8qFH1PIwiNilxq/
mel3G4Nd7a3EFYv+rtSz36PyjdPzCFd2DfJvjPeJYD2MF7S0ILQXmEKlDbG7j2Yu
4qsEpUrH1x2GDxS+SHP/7LSADN2t3FP6Eup0pnUVjvT8cxQbKMs9Sj44xW3djN+a
xZKN7rGH/6AzbV7HcYMNzd5IFMScZFOqtb5A6ag3tdI5yclHcC6pbB4q5ekvYjbZ
Ln67EQwdx0rRSJyHa+wxP6T2Z0qL9hPu8xf3ENcLYpwDMCl1rCqYRDOyVSKxCKKC
CZC/Vcwu2DuJsBo4QUX4myh5+srcadvaIrpCH9eN3ymrI3BSeEfL7g5ejZZdKxpH
jsIe6i0fdz9fTEHt4BH5AO/CISU7JG3ixz8lafhpz1vSxapGI8vJyUB7LMymhk9L
7SFcpQWiCsGrjaCeiXyAVus7RdazEA5T3rHdERvOFbbQSBqmGpLbAkdCBj4pxYEC
MxcVpeE0FognQ5XCnVIXhpomo+fKHeqF8wRWIjWTl9WZ3lsQaynFtQQusT2E5zAX
0F2i/3hvBLj6oGkVfB3YSK3HmJwWtDQhT8fbTViPv+qqGgMAzaWs4GANXjN9X3bd
fX3eNGqqAh1L4N/L3i5pLtRPsiY3NmeDGHGQsnVZWpbwvzSGAqWnPZxgIHLdggEe
IcmCr9JuSLPGsSPrCMhmwRy45j5ylF5EZa1cnmy8uCZonUebFFJXvFjafkAuBqN4
`protect END_PROTECTED
