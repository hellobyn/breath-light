`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9Iy/MY537VFi0M7EZsVNS0vdTsx5LStAp58JjbNOSGC2ALHoyxDjtwxvNMDfPf2
bq1ulLlmxBSJKcTY+s9N3rYA1DFKVoS2bgN4xXaPpfMhPoBWgrGM0gjUksIvBbH+
2VBqDLmtP5B7VMDzPA06AoyAnWBMV9geN5ZNXWj7i7hBhShsWVQqcpP+4UCbLr2B
M3IAQydlqr1CcVhrvaL1ye64Y2ytMLatV06WFIKZC898l6hlWetj9EWcbh+kJRlN
y7X/ZMY+mldvLonCK3TvOkxJhY0YZbCB3H6eH2n5CFzZ0RFjbT5PBvEibj9KbFIR
U6LRZRCVQTbH4UzL9w3/UNdwshCHGeKrLZRlIcrQxWhlwBy/IzsnKCrdIfdREQwt
`protect END_PROTECTED
