`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
es5eFD3OONq0jomrg8jhWPLTylhlkODA3bYxJLaIo9p345Qp7MQr/cwVY1wb2UYL
uTPE8RGgd97DxEPyZNxN2Ohnf/O3K7WpnP18IJ+/ZcFHwP9DAz4pOzKu5B0OBuuk
yOW9yApa/FUth7wNauWOy0bswf5ajGVeo6x7UyBjbN/Dhvpp69i19iYjMh5v+ZGr
Nu2pwDn4aAuEql2v7qD2nRNzvv3lgHPYQ4YaOdLYjfk+eJDxaoX8QmlkmDRJP9X7
ow6RIKj40PX40yplxjOfZnwrhPwwn2OCVmLKNIBDYItQ+bsmt8HCUysUUQxonLjf
o8NhNG0qmZFCteyysbF3MqORE46DfKsAH4yrqXc/yAmJHZv9koB15f5D8UMx5Ih7
hYbPZyl/6kW0wVvUffdvI4IXkLgMaOWIe7Hm7Dcl368YIrwu3icyaYumwpSzYVy7
maytSnmGG2VaLKi9mC8Vtxp1NlbhTirsMPyJyWPVvxFfnUQEn1/XgSMf0r5CUNxO
/X2X6PVtIXwpauuXeqM46F7OYoRM0lQm6wSynptmiFNEAYzqDjv5ZZ32wvKIWKD3
qFXLlOZfrncwni69G2J42w4ggSE6SkNjvwA9Wpfe1KD3yFYO9pbIeaAYcut2Vq5Z
1YpuJE1E7hDtidvOrmj4pMPCZYuJ/hZBvgfjrPEgNgxPGMfC6P9HAn/hZm2eIx1k
PKrrg8AEHlbCUYKFCOrtzrWZaGYfD33ghTw/y0vQ6s+/Rf+ZK+jghLwv5Xl0zLM6
VzjyIZwqz1wi5AGCSPtGB88dnNlb41Z259bI11RnxGoGyAsF9IBmoQhguyXUQIXp
x8uZpn40UjK8BIs9C2BqyV3/SDV5nzGmv/qvY5zfm+wPDD38BTMPs9Pmc/4Fas+M
Bv2tPCKIPYB5NLegPYXX/e1ExEoRz1U7wZu96636LVyeqbytP3VgUeBaFRnIp9Ox
OpMjG7sr60PJsgS3uGTqFkPi9AmVL5E0Fz40XAvPDwrcD71mjQ2ZiA57/8+oZAUx
Bg4kLZGKY6UpTJEEtjlawtHzC6Un2d6Q6E/MSyS/oieLFy5Fqt2dEmeMzMQQxqLQ
KBZ8tBheOOLC3t6VWwFbe3KgIzgIGiGx/oArTvPTzhaBZq1BKEFGxdbX529fKL5o
4e40PmnXOxyvI0207niAoGVPfSTDQmjauPr8f0l6TKOMZV57o8/rzHX8xVfoExRs
J96DCfa1H+VV++AJ1e9ks1FUlgqQ293Ulbsk3SbcPnZcaY3GTTzfNbcgZkiFGO3R
wTMuIv+SeN+GxhSb75fRiF5lJdBAYe2QWWAwrWIiCsRsSzBkTUFPsQxwZnjjSH7e
m7kS5IqzdgSkk69gd2d5SKMoBtQk2l0cyS55IUZpdvwY3kAY0HLmT1wv0GeBW/cZ
NfVEkky3zdUb8uCKB6/enL8RFheqvIAqeMkXlap8e9k/+JRKKu6Q1XVuZL97Duqi
jDvm5nUpOt56mKhNKBuCcCgtLOgjUHqPDv+w1fh9ADbAqku1CI2fjk0FTPfQI+s+
tLP4rr3pICA2yNNQjcw+p2ZGDCjgAxZHdaUF/HA6cXFJnvvtM4FgPWAk2GrRZnAL
0Q7sLV/Y2pu0o1mPv8+Z6z2pPslBERVuRtu4eHec4pOXS68faEJDXdsXa40rXonj
7OmV/CjqUoe16X/EBq8yQ4TJYVJmXxgs+c3KhDI6JHlukcALuMyjo2ve1Pc1CiGC
AhIaICHRL3FwvSxLIrVXCQZdD3qFa78KhiXRM/GbbwuxEcv/hDl+x9DlQb7KGYhm
7IgICx71qTnOgfplPJumFMMGjbO1nBQDrFdB5+Tt2j5SiKPhLHRkTrmZN1Ba6lUv
o+X+TgvymxKnvU3SBh9AYXqjjSBW3UJxMXpAqfuLemX+VhcgnC5RfmJC3vyr+iFK
5dWZgXgMGPJsJKTqMZY51tR6HitY3UPSbO11zLISCF8wugE4hPLekIgjAY3CZoPQ
QhuS4oqGfTRVWtvXeapBzrtbieJmuSvkAOJQEfocbepA3edtvu/9j/kjFHAvJdfd
UHL1gZFXFXC5IVKBKoy2KIem1Z2X8zBTDgzYYTdvDvBTg6LnCqhEcyG3NoRKIeOh
esTZMQ4ZC2bBfD3ce1sNPXZxWGdJ+DWF1wcHDaqw9jfrW6Jg+DlFCBvD3bHSbbHu
l6AeCTZcs4PW6joRdqxYSNU4y/8wx5L6/kTuSckUbg/87d31QMo3ihAuIj35WV97
G7Qbnxj21ph83bcL01aB0y71TfYKLLkaHswD4jliAwdrtIrAOsDcCIWR65B+6Y/S
yMitNh6jeqdjY38uoJI/pdiWy2KQo/RfpHjdl6hzLcqQlkrqZieg3SH9pAray3Ot
mHW2n7FoXhktxotyHaB/LWYAuZO6NAlzfp8f32zRpvJkcBMjOzGYdRr857vcSiGe
F0s5CnXsCly8R0A99vvDVidpSN4/dn10bdNxlNM6qL4MDaa2s++eN06QGSicPSxV
pJiHPzADGtc+hVvWG4v2Al1VUTxVUbQAtD1v43TENH/Z7JggUTwKw0oxUx4OkK1p
4gGYZo88KdawxQQrfeNdxAJ5v+2zyqLwOFWXBwd2oguuawjZ+Hcf/lceHCGJArJF
4GyVkFygcM3DggF6JQDBfb6u+hxNrhYlNlq6P3+5Phd9gsV3//RM1HGJB0e6x9R2
IYo2PuzRoDdmc6goIp/FWGXxyP0gWGOfKL8r0EgCG5Y50Miqo6L381p7vWdL5JHu
hiHUY9gGKAPCVzrUhPQ+Mt6RqXbpxrFFV75ow5FUw5a76FzwUlY0ex5ODr8U0EZZ
rEWRBGJpdOCNOkWzXG9ibwMdoQCklJY+eZNCN1vzSAS5tr010pyUpyoEHF68HSjK
ojrKu5cPDuRJuBqfx6qh+a9iFT91s2vVdtt+fM701sJg6YxCD/z6bMBWEJgCWLIu
wpFnBwx6N5zcw8exz2iZPF1jCxrrFnKT6c3u7vQx2TZghmX+EAwz2u+TdJOI/laX
e4zLmHVAwMKJkTkrD/0rYUe3sCRt9RvBdli3UFxRn4pnuySXNjYrMlYANIjCaTCT
3tR37Pv8BN6lS9KcpV/sJBjU3Ec3sJHZ2Y04RCEvE3mKASghYAxPmpag37/wTWmM
Oqomcc5571AGG/nMww3xcQtR5MAUrXX5EDeHMTq/5h4vjh9mmzbUxdV8oQOSshdQ
J9Hg/ZmZjb0bc8auEEWCcuFUQdG/5QIn+CI0kDEt1xPFdSydkb/eMcwEes5Q2Aos
HqO6hNkUmnSFR1agCrdohPWTgbMzOQgCZDIEmBwwSlzRecd190mjmhkhCxudAcQa
4hJKIz5vMXQ5nCTGgnQLYnRrSFqfrv79jVycUI6ihLtonDeB7yhGLxWftFY8ZrJc
qfpzuhap0KswyS3jR05TqJTn6aX5eQnKGhE01kk46qEFPC4DTo7xV6Yxh7/BcXN+
ywfcGuUtVuanLWnBLCaaVguLAKhMoSYvuDVFIkbXLDp/xZ2NpptRI3ew35ckpRjy
8qUct1d39SyZ7ZprdmjR1uvERC9R96ZdNhCe+j03HS84HOpAL1GoqYpo3QKUnoIZ
EoSzRAyoFjq/NjlaUDyg4og8X0YQdccsdmyI3Sn8yqwgTx9N5ieMumOg71JtK4OA
DHYZGospc6Qzq/F1dqVs2Q+7U+8PvnGbpVdMIuLA0QPfW8adHW3IRe8WuLRHShF+
pyAssWBjWO8szKMv8s/DQtEloG+dmBLEOsxlwk3VBJTWulU5TRlwjDrZIsfBprI2
945s0U85x2yXnxk1p7XTfw==
`protect END_PROTECTED
