`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJ+c4j+mT7jcI9NpckMhPTU5AxmgQ/ffkiphVomOWb/L9e3vEufLu05o3NjyElL5
Whyq8ilP8eKe8Q+9d6g0EgjUxHa33m55FlrEQSbz+j9uAHkK53+oXoeYidVikbFx
fK4msAdcqZDMET6Zysl7rzzPDqj8zsg6VcXcjTAKM/cFvpRQtANWgli9D8GbYKtw
MlpkKdm6xe5rMzbmmj1S5r9jldpOljQIdX4N6s7H3CaM0EgUE2bWmihMRgt1kUC5
u6rza6lcsCZ1s9jbFVrQmgDo8xp9o5PXlRSvKLhjclZJVncY26Ugy8liUFuEOqhR
uSzDrc1zOnJyz7i+jqLlKTbGnm/2kS/5JD16yP+Z/qYlld+8g8/kZSm+YfAwojP4
MhIsLWtDJ/rRlP3PGVvypxonood3jnGMv8+8JZ+G0kSgdCc8ra6yidFPcOcToYy7
akbVz7rXJm2z4jIEjNEmHW2aAlVziikj3SFmoMXR9+w=
`protect END_PROTECTED
