`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nzFx0+lquSXk8kp7DfHt+TJGwR/HkcnVflYdv9h5Jto4E6ucL0EJTxF3keiX97nW
+NUYfIqH5McY1fkl0AzR1KR3AVXFCSMSslzzk5Tq609efdDWPzyb1UXWjrZ8RFET
BHVYaRh2XFnbwPAdUcJaNwtH7bwdShFkq5WyYDrT0+Pn6r1esSyyR9ZNwWh1Wfdo
7khQ+QnxNhGelIq3uxaVhSHP1YpDs3m87/YUro9sO91NJXPPugz9uMH5PRbmvSXN
jAfaRtg8cWgBarBP4vvNegxo+PUq0yrYSaJ09er3Ou2xfcsjmQeglEcs4c4OaYP0
HC/GKf/EcbkXz5MEWIPTemt8gsyjZlPL/CcC9SUltWxZ7OEVTcE/6GDGaKWIXV/n
/CVDUFGtJfZ92iUPatCtGsSLJmyu6D7KD9VIhCwzCkd5K/Ccp7GFUXHMcwKplgeZ
8RyJ5t4gJKou9/akjliaffOci53ZyjIOGvzEVjJ/dCAPmiZGAkp7F3Uxrd07RVZL
9RJZUbwxjy3ggsQeWAbxuAZ1Pr0wbSneo/F38HvDbxR6nhl0wZ/ZeUt2KHJSAiKw
5Tg0C6RFm7JtkmPbDkEpKkwliwtjcl54Rl44uZmL72COa+zO9EqJcrhlJ9oHLr7r
nhVWi6LGhsIb6aUV04HuemTzNHUc4qEfGG4Gwlsbc4EOg/2SqphE2/wPSyvXnEpB
HPpLM4h96FOnE96bJ7ezbjf0hw8VvrqrRKMOyPBGYmglcII8tnyTl6nn0/nM48Su
AUk28bNVUSJpYqv3VAJEXVeq8dLG1p7u32l7CevNZoPuntz00KmwX3qalVYyFcP7
1WN9qTfsza6/zPC4X/KtI0i/QkMkS4iO9nmt7PwJjg4hfrE3dDN06+3YX4thAJc0
LSDA3nL7xHLpsG10CyRdSFiEh+BhcpLVl/L+eJtDnfFqOeUNVT+wqAp7NzkAGgwr
Sk+u3mYKgV/HUwomiXcBMD3LveoUOy8K8xpgKScUOvEQatN4XIqEPeXBOIhNfm9+
D2r3UMcCRuYP7RKpMuM/iSiBUaz0HNV/Q8vqkaDrzGPM+OT6uRYuLqObrcC5s/dg
xDuco5xJYKdUCoABH3GZmIPTwXf8yzQOD8wafJdW3Xs7LYxUi/doaDEC9Gz+njLL
wqKTHl9BGhXZqP7BrAKF1wbRpu/lX8h186l3wQC+0URKM31Ch6wnEYQnC0bpOaB3
Jn9e+qmA7aH5/MeNXVDBJ7q/wNMJPfKP07VEL72p3A2QXrfdXLQiHrtoEPNwf/6q
e0s0D57kv/xSmaJ4/rBndP04LroDZgE5uXMRk1EMvm7n5oYtMIYefwOIrrTmh/1l
dVepmIJ82QTTjks4zn2/cCBc4OhxeF6hV/DitcXbCFZdN641WrTv9iuTPSw0BQ9O
Da44jJmI+6H2F9PwiAfoqxDzb7IIk0pQzuh6bVCXX+2rc6EZAeLP5woN+WNxyaf+
fKWsxJ6rjYH303ki/cbl0HE9RPrF5s5rRPzg8A1z16E/OxEIENYRLEemHB7VIpfm
Ot/hWdMT33vPpO0Q2uMlxDl92VAAIvGxKr0Vfe/vJov+QHKZh5LrGmVBmFtfOMR4
rLjXCF73XID7RK6LuTlg9OuDSUdgTACdO4MyE5UF6gFdE4oSogmckSAPxgh1FKxT
mSlDakAMrO/QCG4yJ6FfsCl/sS+daJNtCFPkFr5/bhyo/f/l04yh7KRjH16WiIuL
YYoE2bv1T3Ksnv5t4CXGEg==
`protect END_PROTECTED
