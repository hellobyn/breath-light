`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeyVB+c0Vyh+acWLFVcM0sAqxUlBXOHGJH8G8U110hXiR7xDg7ThBNxK8zDZFiZf
uPDhnYoBca90RaAxh3yC/gtQYx13CWCu8eig6TNnfzFRI1QMGeftqxzActqn1af/
AKaBszNkon8gv8NrM7K97yb+3Jr0K8ss2757dYWQtBW7flTDIV8YLtPjeKNYKorJ
tiQ/JBYOoXKgOuN/jUWZRh1Y0F5ooUU0YLNQBClGlIrJKfbVV+WTSkW6YsK9w+cj
Oo4SKv8AluQpr39q+1nA7dHiGbxVTnCIXueLYGWSuZidYOJWnJj1wFuoKSO1Vr79
OWf66OhemNj6xDaCaOsnqMP7IteKeYydIsCR4tVkXPMZqz3WzzZN15WbxN0IKHNk
bUfskP5qhlZN2L4AcfuMPa+nVvLvzCNClRBHpCkKZLFoFy0+pqVzQq9DI0i6FHiJ
Pn85C/kgJCtQy23T158CdjiifJRX5eVtF4DFMg+J4UZXip8YdxZRPayNyIvyvz/z
F0+EYCulL+OSI6yLcbWYHix7aCpV34JSuB/o4wK2w+PwjSyzIt1jmIg/KMShYbZ0
gXBOEK324KDdwDsaawGtpnLhcF1jvFr/Oqr79EgaCNdPC2v3rvtljpIo+eJOiFcD
Yn5GVDR+xUdp6dKOmxEG2eSxb2UAafOuFxRMP3rkTTLrrHJ6P51+4vXoblgSNA2U
EYRWTZUQ7wXLN05tm9niYd7XtMODkOehVxcNOqvfStrqzh7NUabhoMTDUB2P//Ox
TU1vOx3IxM82+S8JAOskbkexOBOfqla/f1JouyoEgDbLHOLqmmrhKAv+vorjM2m4
CPaKnsqKW66P8nA8r1zw6ILDPE/Ay2JlMhftTalJZ4GEaG9zqflGLNA71h4QdV2M
Cp3GYjDZZJvPp+syoElY3E6TV69il0lHEzkbySDJVKc=
`protect END_PROTECTED
