`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EhBdzoETS2tU81U7YRZKfCzAkX4A4k0rHb2JGD/lgIxlpRZCL9aJ7/vSIVEXeduN
ZobcBARlIplh5whEISUSkotO3vDmjRD3ldPP1PvRHlHGGSZ6x93MItzD1Aq85UMx
qPdCwjRgZ+9qzF00R7O5tcEiQ8aR0pHCkLVnmPTL9zG23/Q7x+2nNqdUluLsgVqv
94DPsb18LJn5vFyowoGhcE8ism7jvd5JBlwk3G/duq/uT/AENzAEVBG3Kl/Xn3ZB
sG+L/GgfDIKgTNO3V2tYqy/e0gPe/zeixiOeYjGTne9yWTTUTzZKajYZgPme/mAI
L2QvHepZM4bsddP0h51TgusQ6irvOBo9yIZW55JJ1ZSv5I99YLSJfOLQ9k2KMWbu
lOoSTAij/k3w9MDRdjgdCi/WiNTH1tQvm4pDM4aUv9kFpPIgUFQaNQtY67nopn4N
8DUYozi6piwYEXPAme2O+QI5JdF7rwPsQh0lybmAh+0kjC+5fNblVPCviSBPVZGz
RhfTlsuSygHQBDUg+758Dz2YtpydmLEaWTiOQvlLGCd21PVzVheZ/4Rcz8Hhx1Mx
ffTWDceUuVjE8p/7NwnVIaGVZf5fei5SDaypEdUwGyyKEmvKoSYX5mT0qhnMDKh9
c8GaFsYjbSOke/ue4eVj51u9KMtlgVjY0NGakJD520kPtOmQOvswbJxpA0qyN+K3
m5/Slsgs4dbTNDmwcD0t749wlIWHx9rWFiFaupHIRQx3Lft6OS3741LvBLp97Jev
zGYReQKnmmp0/Kti3rjmCF5vDxqNgEd+D4kgj09X/JwyHlxzFW6ReOq6FHYo0HDd
5iEUffq7RoZQQ/fl4Zv9A8WytsF6mGPicBDeP6OWkzIVVLof0jbXP1yNMmwAwd92
xjCNqptelce+12bEdtwlB1a9u4Axu3BI4h88LcHGb/jnrEKy/UrDOhrCz7Lds6+0
WBUFiNrC2H11w0jLCVTsrCU/ZAluKzt2nw93rFKQsIerlEw5eV/8DR3Fh+oWGzaF
q5xHGuocyo78u1fkxZPRoOqV6AYB5+VM13oEgrl9qZlm+mVHsWrKcRsbuIiP+y6L
VhwIlK4tDcvSFnIB67tFvRh2ZqhGOjexZeR7JsxkF4V5bE/2VQEUNugNXfwrXu+5
Y2i1+bGM+kzBfx7W0revEt6icH/YpODBe/ACYeGTRNPmzxyIwULGh5ONLKkUwsuL
4lmtRFxnkc68oTisueC6bpMjyvSdEeosBncgIfrewChFAj8oukxg+Ldw0aJqtT+m
34qPNFz0fyH2anjxyl3+vwyBG5BpIcwTBA1lNAGc61HrMzg/VtUxCrPwtHwqqkn+
93EospNpRtbH2dZL03KOD/lF/ZefV11eGkcL1mtWDhBdi0rAoRpN+VLKrs/HvSrK
44lSLtdIkY/dn5CWVGkopOKaXCelym8zQ/vIUAMIo/4Ox7yPiE5fIaXtwc/O1c9B
rF5x+VRsbDAGf1oLDeMBBvMwhtjxyoKfuJ4gVn+/iz4=
`protect END_PROTECTED
