`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s28x5zPSiH9DkXAzVsiNx/qNAz7j35py7vvyVtGCHroUVzC5Mg63TZ8bVgNI7Rf3
pYujSoG/jhPMSVjH9yi3EXElkax/QiPcuidARfbtY6wVoj/gaafREJxLlwNJm0Av
EcwUfWoqaHgofLfhBaPujX2FW6C3+72l5p3oA2o0fbV/xoPDrephklVJLd9W75K5
AW5g2695sBMZ64BL9lf8GYq/F0IkLEmrIgH+l0bg5eilm5H4iphpzXXDKlSOMwlN
zRX86Wcl9qr7f3MvwLBKn1V+nPi+UWwokp0NeIJS/qXDSQe+64k79c4r36uCMOPE
Oz9c8krHCYvEDsau8AEvJOykjFY4gXaQ5V/7QUY+iq9bMQJztDA5Dr8X4P5uOZ7f
J0fqpeNLs/ZJb70UyarXa8E5s1Wl30PWZHYuDU91J4HymySvYJyOogR21c6qX/do
hbCm+Rc6P9JUTjxdlorf8magowSE95olzt6UzEbcDrCyPheRXpk4axV4MpjDvQfW
tNjBU6UZc+stnj5jYGfYlheIvbSAKL+qFtTlTbY81AdGqawWIWrR8LCiNhiIg60f
tRYG2t6E5G9zXB7y6/8RojkwjI9RN5Y6w/fIwvEMj00DVE1FJkUcUXZUTWcHPVdR
ZNC64LwkAN/RgC8EWnWPZuUcFuCffZ3ZuMZ9QibFi/TL2UQ4L9tmSgrrRNZ7DyHA
j/Wl+j7nqoitfsNQw5jhJ+tyDCwASr+YFyApKUq00fJ5uYxf2eBGNlrQYbEPjwNa
`protect END_PROTECTED
