`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZxo8w77CHnR+OFjFuZOIgJGe0T8gDbae2M6bZUtuPMF9shwHTSuG7PQ6s0slKP0
lQOzBsVX8dJwAYD91I4eZodj+gfKn0/zLyRUl399ZuZNHXoifPtwDzcWHirkXJES
QlzVqxqDvm7Zityx5AodHqIhzcCuSjDWde/yjef58AoQa9/bhO8qY5CS1CKPUCrS
/wR6v7c0ky/aqR+MptZ6tzgaIaULEyq46vQ5eEOHI7SdFIm1ppqJs2q1XcyVsAk+
9nk+TrIPugq1VFrK0HUjPyK+r6iBZDvFTjicLKlQoYjykA+8FYKeqben/SuriEWY
7eDSGe3ISkM5OWYy2pqT356VOhz7X+dPX+6EajrtNIZIPhMcuGhJeiBYOjlS+LRB
1tymZA4mOsmVQSE+taG0xv2lT2xZ+2t3/6W3YAPan+0OOLczQJ4N3f9S3W/P6YXn
7cRre+wD4VBPV/5UEevLKIrhkbqJCmEomNsBd2oo4S5NikLotQf/NSKK4LACEZGB
d4q9JB+mgIpszxBLc2Ea6ssEZaFU0Seep7qOQZi9Qc7k2Payuikhn+cHxUFN1USk
yAwVqN4lf3Sjs9g2Xn8N0OVIKTI+AEn7tB+isN09a5NZcr54T0GBUNbAF7ViejlO
refHvxQ3QZ0MqCW3zL4GKYdtXFziqI5gAVwvIYTLwYFHyJNiPziriibk6irg0EFT
R+zsiSQpoTs3cPbvgt8ih3braSQAyo7PpR9cAOaXtyg7BKODqAAvXsNn0zKfUbJO
JV1Zju11yClgy13JM9nJy75lKM3W8ENQ9lJJ/oObTQA=
`protect END_PROTECTED
