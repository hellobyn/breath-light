`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTaRe8lNZQbZkSbO8z4ulfyje1pqBVhQuEOMOQTeU4XnGuushtC9QI1Tm9S9drtr
hwl5RSsq8MeT86mConEGiUbPa6p2PIgP4qxdSC5cSm3riV3PKFxHPMYNgxQ+ovZS
uJtBEr8dtxbp9hMo4QXSHXvzAv8XHMix2nE37bS0Px0bhZM9QzuTpAwilWt3D7e/
0EnfNbQHEGYv3ogSrabnVD+0gn3AV7zxYfcQMotN0gbJX8LTVgNwa/+O/RKre6u5
F/fJXv1cKzBThD/MhRONaYPejj2CcyfEi5DnJa/34lLppQuC7aN3X+NOi371HDnl
VlCfGti5ptkgBCcGSOAnz61CE98su7/YzC2TACJ9lvij21OMrAUuLq42HCLKy+Xd
LnS47AkJqzhb//Igc/DJvcyrCBk0rwkX+6CDdbIO64rSWAfNt0UIdIWGw/9w/Fn0
Guy95c81U/UDR7F4lHPCQ7devJ7MwednVnQDWcwg5g0tYwhG42Nq4ubiKNtoGsTO
8Hk78/0sHPek7ASonupVXh1vkxyKEllEihjziMVwHtNApPzeQBqZGwO7kjBFla/A
qlW9Y8rJfICcVPeGK7B66wgLwensjHmpzGY7O5E+elqaaXIU0FA/24Ki6H6r1E5K
1OlDGrw7kwBRdEKSS77SahSbp1Ty0mHbaQFxk8+gC/MbZXcdF6jOntrvEa6vtfRQ
voYtakS3efR/ANxKbTnJLJYVCFtZ86hH5sqh88Pa0/mpYKtJuHpHRCX3+rgB5Bzb
fDg3vsv+v7YHiVw/O+7WxEenPxguZn6VLXaIn5fVZQ9prpbsERk9OUy4XWAH0aVR
gvVKL7MEDnxzm1SNyuB3YEKFRm9iuS3vAchQaD8MCFT76g++190XUak+ysW+NkAZ
Qev1WEixyW6GoqBsFXUZPMGK0UR67Rh6aV8WFIpGOg4haAjLIrwVBuZ6uIpDAN1U
2Fhwzp69m9kKcYu/f4do/XZvyHDYie20WS9UgmQtgOb8PGuZZ/ILYnlgCiYlg4ew
xuhafzhHtXb1Ea7c8cSy5wsy//t9JtoQUwCgCC6CzLopolgJ8fStSZxDCg3f1HTw
oDhIrPtGwsGIMeEAOBsS71zgZVZVEFSOwYrQUun0INu11alSrVGwSAKuUzPiXe1U
hvCmwDNylrjFuwpalqn3KyliEVQg5OEYG1t56CXofgPeuz685uW3M14LR40aulIl
QxGu0KKXmU0acyLMZ/z7/Edvtrd7ExqtD9IdAlxN42NqAocDisglbbh6Txna5ewK
jNHDtebNfTQX2VGM4LNP/RqsCtVUovth2/41snCgBMq3ThY6MClroezLUOt/OobE
4ipv/oBGbjyTKsLA9c20xe4M5M0OWqeUZ1W9/g4P0/cymdnzaDwQgL4gz3H8Uzbn
gJZyXYvdYHYB9kJeThlv/KxAfOs0XGebRxQ+cciNmASFuo8CfM29ecxEDLgHD/sm
BoCizvip1KsstWCshUhOJttSkc2ZxUBvgvJo/zhJW70f0f0PF0PA6jSvgWtVhThO
0XkqE5uEYbRi1rdGK/m0qeelRwHnMgmN9JitRT/kvdzzIgpbCDIVPKrHpE5flz8N
IpK5Q8ZnzDQV+lh9e9hMvn5kBthUHllxi4nOL+4FPUO8N3pyz/yl54GwhfMVTfcn
OC1OecdUA932dybWuV65zPsxk+6X4GoWnoL9XjPKvEN2Ws2MimqXVS/cviuT+0Du
MHHzMpEQLBTthkgwtaw8waJgmlTyaTlfs3mG9OOKVQmiWMFQjBHiozk8w3DNh++H
Tdv+knw3M2Qh2psASCs7BfJawUIiBunCBRrlncatCPjjOAssRYlE7iOf6FfKbCbA
XPv3OK8CFvYCqImDXOOPOOcYEOnCpt8IYiCQY21g9b23tfbcbm5CTcMWMV8BV1GJ
+H7ht/tm6XdZSIBXVA/FxAp9dTBAVvzPPqbGsR5FLfrilDeLfUaSkY7g0VfE85+k
TNUy1H5QaKLi4+thjkMsYLlwFipcFepGdxPJM+p3O/sauLVqaE/XLnVyGR8IzF9x
g6YHlVZ4jr38x0gfvJrIrvQirJG5MHSNd3v8ucWnMEL+Jx+qHVD/+X9IsFXZlCBI
rA1aze+CWtDY7OuvyuUxUz3yDCeolphAjTTQ3NXy5NYeOkeXr5IWszbgam6kGDry
2GBQSUJkOrAjYy3gixii7Ir4ItbsduQcs3uKmXnGKhXrz4nv5Ar+PIWOEU+w3EqP
0+o07iGIFbOP1GoVsmiBtduomc3Yl9JMc6EMsCp+1CE9zPvxm7i8InQHkkQJXy1t
V/3zvJC7qC9qicwhl0Kal6FFpxMX+GFyfnWZd7LlK46F4wXD4vAuuw7HP2lK5KSn
g1jEAQ+VBMuethd7ZegsdBLe1wGt0+rJ5mwTy1U6buXIhiG/yMq8FVqpX8DSVOHI
4rL8LDy15VHGkYw91GtHcclI3t0m3w4v1wfhJE8JGi0CV63Ix8hJocxeFZBh3FCW
pK3jiQ9PngVtz4lmqnJWzVFkEwa/gyo8L5eQtqmvwz/2AxL96yAvNhmeGcnJAvEv
bZwURhGHoIRBf4IW/SMxRRi7/XxgmOnkbT/y0Un8MQIeI/l6khOij0g88xC6pwmV
Jhhj89oHKZev7O2xQ6egU6TvBUAdvGUgj3XcqeRDJLCeAmVNwiBCOcNbphuqbRhk
Hv457MRJ3VTWvLtPFAbdA+qLukBohUPowAnOQkyl18JxF68/BY9woBeVbtuJH/BJ
xAIYCCU3B+ilz8pLCDKZbpqNWCPt/fFNIyo92aRaIMTLCJTiAD1jn9t9tCjw2Z9Q
dDm6WH05StSxUAwzqlejURwkiHaFbJq5wp7cjJ/7/vuBeH/INdUAMZf7YUpowdcg
oEZCQ2+gyAzeNLbQBtOhpf9LRNkhLVkE4+L6ueIh19lLO7Z8VHT6umMwz+TBXBOm
xdqxdJdF558aU92/x2LPgtOip6ScszOazZOTboiMJPJJzFcwfxs37Xdk75rAp1hR
U+ilGnB1wO4AILTorjUrG7mZQnuwX/Tv53sUCwrrlHngu0Bu0+oFyOrBMJE8rgDH
Vf9twnxTq2jHW9XvcAT83XVUA/td5D6j0HbXGJTA+C2syOzMIeA5rpZVjfO8bDF9
T0QjW/l4DRQc8r2Gh1B6dCSJjFwXXYM+pDT2PtU2ICE049RyM31eioJrwwaBXjkw
KUlQRjBDg8z/CM6qmVuAv7x2xZKZBfSAhZB06URQRNDXWzvrM9jlcI5hH+3PP4P0
/cBdxStkJZ9PdT3Mt1U6QH53nXAA1eUqtHPjaLRxW5Cy/uaUdwjYfzeV2HsL6rGq
KJRnYa2kaiUfZBhYv/6ogrhIMyxdA+jyNkbtKn0sfsn7c66/jqK25apuEUYM1FzY
X19aZaARTDF69L9lTlSTqxI/PzrxjIzUpZZQXJpsjbEiOtGSJDTqy6ockkHtrN4b
nKA5EGwY7SZfAkMw/fphCeNrnXuzBcqyxdAcFtloKY7EXA2HgHmwiRxsANUP7VGC
my1SDfNuMJZQBZRsMJkc4CQ7buEGLlX9+YEt7EkCxeh5DvRDoErJ3OhAxGPA1Qq7
93dlYDFT+3DD9t7vDCQasUzBYJERroCdMQ4E1MFozJy80fTKGVxhkBBkZ0vrR5C/
x++Llkll6VzvRhHb70kmJI2slYzbRSGxrRcg+6shPPakpDG0GE2Wa04HP6VbORho
UllTYWRAZEqyTd/cOupOeqO1kOWDr1Rgzi4wtSs351hdkzLOXaGZgPNX2zOag3Ub
vF+GSUhN/7K8YMb+a3R3VgndmZCd1Peel/4TRvUkTJfo0CGKi3Y4bG3E03a3xMwr
6Pq4NZWja6BRihtCZ68xIQlx3zTOPy51FMJplW4/vOY=
`protect END_PROTECTED
