`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyyl1pq47I9hCd7Zk3biI5wZ2yUUvns7ARXHj9ft+SAqRgYVyGK13/Hc2BQ45mI1
G9pv0GNUMpO3Gpz0G7D4YqjAMi8i5+6zUZ+7+0NkFuoneuF7FYjzYBdOSjvgxp4y
DK0ETidRf2LyyuA4YP4VLrQ0KR3ueQUE59aQ9UY5iJEklkBo3RvL7NKvyIX6ZmOa
YjeFS+eEziYbgIBiwqEHZRG5rGKxFlVDTZh8Z7r23A5+ZRnGroryguXvgQsDuiJA
Jr0YS5kz+T+xtop2EaGpUa60W7G+o9l7q2L6kJzDtJb4sgM8+V8wWKWprZgw51uZ
t0XbXPGshLbszuSr3Hh1D4uS2Fnz/g9tYC6KxWn3sRObWKisDfZHQ+96MKlUhJZj
qYv9grS2j8t8uhfd9B4AbvKqWQoXnXdmtnl3GYvECb4Jh0l1COpLwOQblZKd5bZQ
MdRrVN1AaSYE2HSu0pTml35Z0pvrgrT512A48C6EKMgy3OqOykEbiMuuFPN2z25A
7ByOdk5aSNveUn+N+X7acPoc8J7wAtik8yA491G6DAh9mHXzsDciKSQMAR2KUYyq
3OUtvxXgJ1qCI/SMDibHYvdTzVYYJ1oleDwqixwYPPdTkmlH99nVbIVtyrE4RYgy
1TO3OwIExTtQwHz61GoFSFaOOewELXl6/p0ErZaGzB+tiKzxdNGHIEFWSZx7xyyY
y3BwvTaRxIQ3Q2lbIjtRkPFnBUKDj/Vbc64ip5eT99bnrwd+UPhT9o3ggpWoqMXE
TTYVnRc0+Wd05qvmSyTCAN+TUwPZfRJ9AeHT0AZcqqpDM9BNX9TV8Fg4O3kOyUaV
`protect END_PROTECTED
