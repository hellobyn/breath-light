`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fonZ3ZzKs8Ar2pmNBus5gQSPLmKxwdHS/cSRscLRxq2enerOrmV0EgnNJAzcFO7P
Jt4w2MpUypqYBfSRZ1uWanRWQyDUhXBsz/XwgzLvTFAn5NeIlPiHgDOVl4NqxDJe
ZvLZsczqJPzrn6OAC5SWDNuuR7RxWHymdh7/PYOBYE9SCcN0ZTWiNnUuciVOGPys
PQSM2qUgXXrKLsxvnOYQuFRxWTiOmq6Vn9dTTlhOcRf/853cMpNExbQhmA+2XdIr
2wTgrG+XC4S1go+7aoa7k0NtYgpikE18rNcSAQdrIPNhe0cnoxR+dmBhWk/gqAnk
zFsurj2356r0YcTh0Sof/DyswaLKhqDvx4waADTPMAX/yU8duQcm/hewEdXuzU/8
Ot6nytNfv170kNUaU4YLCoyt4GoP7biBN3rFd/+gPF4w+8flEMlWohMhcSb/uFoD
qKMKzxrzPnLjua5Gbhk4343vpo8yTQdbXLnsWu/DTbtLkzODEiTGn/F3/V9BKq1J
ofJHwCZFmyaBO7p/5f7oPLUnT3wwhypdat1mQLZx2J7f2BwcdUtM+qC3IPWS4e2x
E/AUbd3tRI9tojC8wPW2AVGBbOnvDPEqp3jN8V41ODC+E2NCMkB39t7lKTvNJ6Ca
S9esTQXU5v76ZcQEVXYmkRMzKfe7TO3fecCrVDG9nDk/Xpp1c0fIFazPTvry/Cmt
t+fKG/rsHbddOmeSZk/c0SYd+LpfHD93NBpI2wIMtL0=
`protect END_PROTECTED
