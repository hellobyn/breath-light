`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7ZwNqyioxJzIq9v1P+QS/XGcNHBGelOZnDVF2sxli6jz6k9ZvkK7W/FMpbztrl8
Cz+mVD8GHsJvXDvrfr6CsCKcGVgtrRzLA/v8cJ9+2+QBZK6SOb/CdU8BwPAHOHq4
FSLdR4xQIcS+svMO51cp3acnAfpqg1MtW14PjCX6+3vfXqVWV7nimrM943ocfdXr
5B5v31JHJek9bz8AMwTCyKeJzE7xnNKqW19vCzdUOxb5Cc/RFKumyYExiWd6E96A
fr9UeYp19MGTjLxbvx8xNFAB47GDqvb8O38AKMTqW9eIygccpaFA6v2L2IrIGw3D
g5rSyT6+ZREJY0r3SSNIqNFVaHJqAVfUCGofM4E5Jxraz/wR6ehVFxfDpeB+S2tr
EhhFDNhYUWCYh758qZIImu0u42o8jkNZc/rEPArYZN5TNMp9mnly9BU4KmHlqOhZ
tP9vvWUZjBOdQ87R4tfpgqGQq2q1DmFJZ1W8W1xHAXLSt25AlNR8qxf/NBE0eDYj
aldIw83g2B6Xq4h6hIPRskVIgZjMnzS/Jl6NnMhim6BflgqJSvYqQ1UCP+TlDBrH
hDtCrAzFOUl8p7jR1/fDWXs+hnbhVEFt6wzW5AKnliZnSVgOMn/4SCs3BvVkj4Sd
5o5QPqu3V7U3gbAG/sxSY7d0OPIM3FFoHr6EBxDuG20FCfp5PP1JnAOy40bMwznj
8qFWlSNKW7VIP+yQG3Qwcmd3UxQEFM27ERCEdaSC37dVOavbqeEOt1IM0z6+KeyA
7lYym/05nVAej81ss8wU7epB/Y5lkpXCME9RdVBo0zD4VkE21Tm+ad2S6YaMLnIO
AVQE48w9gM89MyIS57OPFzK+6XxBCPes27Xv2Lnjst0MgVjQY81XD6bUoC0OStI4
N0tkWYIZ9i4TImo39+U3S/Qs3zO0ZZDm3mcR0wRwQ7ObGEXPpvm849QHR63ZwW5c
dvkwpWpBlfjBIzUSqriLFEtZYg74QD5fPZcHAyfjLOtJPFeZ/1ZjV1D2iYXnDTkl
57AKJNPaQZLUv50uHliBAjKjE13Bt6J6WzN6YFKBtPF5mavyj1xZ3TfNh7zg55SK
uXz1uzRYLP20kPhXllsLp/YMjOvppDGGxkjAsVxL3HNG5VK9NjM1NNzKXSsD1rv2
E6kNvTwrCJAxsjboZTeoMSmf1q9yzQUFZP81ybD1urd3eaaUAyX0K5l7BId7vWTP
Ys56jPcx+PlxIUhbt4qwreeM29YEGhOVulDtTxQFW5fUD+U4QNQugD4S36l4vX7V
UWg5Fw7fZWiWbCflixcT2/knU+bIbgYN4WXPHB4xuUtTanqbpzpA1DykvilzhQxv
TWqxsUZo8ROItMx92Mi2ApbjSKa8s5+hjpVlcG4JHgmewdH/pqnkbDvRNzqe+hex
mNmoVDcFTwUBMa3iwLhMf9bCGS3UVnGgXSXMkdYATGttMYPVwvxSvnlht176F94w
BoeXJfo1b2lFKO7KfK42FkjR4pPP1DU6hCkanuZpjjmnjLijSVRchhVcA1Rw78FU
5LVhdsBXVbMGzbiJboDewMQHfuiOjMxVkBiMI96+xHRSiAXd7GGt2eJ3h3E3jhcQ
EKgElaXdP1WTJ3Njr6hZqxw7Gy5AYkzZoq6vHTUhLoTbir7up4vCRjErFlWJ32HJ
cdt0wcEEvG+vQ3ooeIOLgUGVyZprkSzgYYtpuFrhk6TMWjR8Pk8gDHrH5AA0mCaF
ZGgBWxi4eVyv6hlHEVmV4gOGanaAug7QKwHR8xBl6WS0HB7vxK02ubLQ+2TQBdOS
/j54y0F3bBrXPBzcT8tEFn1wewnOYx8nAEEOSwP9tTLM4apsNGRhvTeMrzuMEvsO
ej0XxzJR6t6aIn73S/+TgG/IH5+9/+ydDtWZcJpjsLWefvOiEEuvqIxrmY9f4eQH
FlWxMMpsQfpHExtGVMb4HtqoLjcP/u7FZv4Nmnc1O8lthx/05PREqsrYe/L6kXqU
Rozj2anKIOnzRiF8C6xJbsXYRfudywD/g07zje2a3zEqXOYZLLpWG1r8x85UfMiA
a/laSgPXHVbtG6ZQ4KwVAFlYnYfdhF/dxwkLR27cBQozXOczQaGLnslSV1R1p/0Z
h88+9E40cK5jpLczYpGbI2Wohu7PlvNxwDJ9RZi+s9CTkPSGmJV6F/ikUhxYOTW3
cKVsm91MGTkBsIY5ccJ/U/0P1u/1bDAJJ4DW0RdLCcTX5G3Bi+soW0sjj2nWYIV2
fl0CBFkoC3DvSO56eQ8/F5vAcCIljScsXgY9dIWjXwniRc6ynlMxcMMNERLf0iAI
zrlmtCvL1jWX5RURM+En2or+hKqnePrAylUY/6yEi+Twy6I8az9Wg9IdSE9XloT7
sU7z4sJcHk4yQZrGYTbL3EO8CpZWUU7lXgm9YOnictxNpCUERsj+dma9qcJNArmv
zis264ZMvTb4CWklcsPaR1C3HyAOjohO0O8b40CbHBFj6zkvZ0+pVRjR4TYlhvyO
V1rPcKRQYZYmrOduAB3KYydPrd4JIsntsJ485rFJxTrwVAfaN7KmvI3dKxP4oHn1
y2B/Ep3UYwL7yAJodFPKzQANZBWpVmyfFZqXUB2Set05jrBTdjNZDxWSuLnaIoV5
Rql4rkf3qopR4k22p7iObxoXvNutuwOpb3EvY47+E5ZXK9kKMFJqHPTk5jth4hbk
y7UdVhAuxztJXOgrEJ8SMgZ6NLsE1KSr82xnd5BYfRFmGm4e2Kd9ZcBXIkuHQ3gG
KgP81uHFA0X1XPOu1BwjdcMKu9cE4vplsO5ngxlGXJJGmtZdFatjzHEBFMyPwRDV
xW9KWUNllFY6sasN64UVRzW+nmXqfsa42rU19V1IpNjH9FTycPtz0ULy23PeS0+E
v+cOMzyhBX2VB+WuZoa9gNI61azHSk893uQLjWOUA3p1fB2bHYAfCw/SHgMEBB+M
B1wwDbvqVTya5PQcz/VmT/BmyEiCEgYc/CUgJKQ75OfK9EsIPPkvbaCKtaoVLBdC
H2aRTND5pV91UHRymOtyzYVnmF71j8GsP1qr9xOMZTZjtLvaGB5STO4tsJ0CbC6H
lA/FcaduwTC8X54625KXPlyEfPRgtiWMMEOKeqanILNgG0H2qkpV+RLu5V4Gmk9H
7z3mcI54u5JdY0+7aNduq9D0F3FNHyPVXThqr0ohfHs9n3KtpbKkPWnGRbKii/Es
buQDPtv3ta1+fRNdh8Y8L/HHfNXP1DBBvWK6Et2KrzK5gPmIBFiNxxmjJJJ6N1QI
s+d4UoWQ8izTGYKwKcDz2ccawEAAFF1sBbLLI4lxE41+up9kWngrqJK1lZTLRvsA
b/whJIlC/XckETs0Uz3PeItOAInink3Tf5DNv69kDd1d791bEOB7iDbsZOPEPhVC
+4CguxVjnmDXHUDE8EfKiN2HrHBasOzFF9qgAyE2QF/KQrWacYscQoL7ADB2IDrY
ssFcHOG5nvvrBG6Vrg1vHH+BKz1eEonnhUAtuCOzsQzi5xVFHEEjcryW+FeA7dVW
fRwcIyHisfaa+mOUaDXFtvatXsR0E/teit0ABHtf3uQPbkH2nkJzRYDVvZMclXpD
q3FJ91EkzlaV+Ndu4xL2FZlhBb7iZ3KdwtMpKnmJBr1nHS/j8yly2/9s7h6ePC8A
oAMcUA+CANvXaJcJIp7EjhQJgdJdu9otT30OIdYElEDNgJGqBGvjINfJeNN8gmbU
+gNr5XZOj7Do0UZwTU5mxKgViQtWaqw3FpMEantFDUX4OuA1vnEJAexnZjJz+27O
CRGnXsSLOrotJqUhWBchAoQ2MpaJRIa6j1MQaVg/MYdI0LOJqF+24Io15DOn2gvR
45yUjRHqonQI8t4m5r4PMPJyXdH39/TWEejc1+V+oNvmXYKIwM+tsH3vhoX+V3vB
NDeF/7U1hGayXC9ZM09jxLwegFX0OmxvOJ4NakCtxtIV1mru7gvRA2XapwqHTEub
o13vmDYz7hh5HmZ+YTcW2GbX5ijPiVKqEfvWFbej6TTFRtiQ22rSmgIfGZ6YFt5o
jMhQSQ1Z8BUX5Q8K6nFcl5H6qHhd0JvMaKENeGm3yGXXaUids5yp9ULOklg42yG8
aGtq5G5P8bla2plWxL5hBsIIUWBtm4PDpWagbdyHn0AoOgFMpVz6ugmzzoJ3BHAe
QpWYYy1Uo3oHR3OaG20qZAyomaL6pkpTVcyYyAVeIihZoGUOcwDqJwnY4r/SQs3h
YKVSLXG1YxnIVaCiE3wlO8K0Jma8aZbZHLjA3wbZnCTwt12FmH72U5XBLu0XJcdc
SsNVU6Z/nBXRyiZS5oxabWIE/OXKzQN0mJIf0Tjx6toNDZzroyZSsiXRo/v2ch9W
NOU3DWUtMXq5QQZT9V2KfhMUGbDfsQTiYyL7bOsm3TltWGFcRAwb+BUJuQS1AXIY
kdWx/sn7nQjpVt0UBkph1d/01cH+eSgmSEO0m+zLLr16UuhOBLjJcoatWukiR4G3
GyfNcRKxUULkOFLvlaAps0B7K+0N9jEZoPi6wgLtjEnzGufFmB5muLLP0xT7/wEo
joBm8exEdBPVHQHv7aXC+LTUH3DCYyquWNUCClAAW6qZSth38kvpNA/CEUt4CJHk
GTVxNpMSU+UJt4GgF/dFHjFvb+BMCXwaqUcWlfVTKIch8cYEPkVCBJO8wW8PVsXl
sZ4m0xprI8Sdfwgn1a0XG5PWF/TcX8M8phlAXcGqUkPlfgb2bfMV6O5hipfLYT1s
AHf0Xz2Joi1j3gsX2zzg1IDKdASPMaIDDl5gwQ1KsZdjLKq19KVEp9sT5cw+8hDN
7rCXT0f8HZ+N+oWdBrAtcDlQGCPVj3XXcgJrsrDPs2ryayrNKeWWRby7SjL3H+2t
tdgq2aZHw9ehS9yY6ea9gBRFRuGFdZlEprvM1DHA+bWqzJQ3EscGl8HzyKglFdBx
56Ef1s/S/+XSklzBASxHmm5L8o4SjAP/KK99i9pkNmqcLjPmsMtBS1EG7yLG+x1d
35DX4oFgS1Nn2ZiPrqWva8zbnmSIDfUEpULyXrfbLzGCGd7bBys62JxvCnW4s23e
7nSMPiFEdws9MbUqfNU9kwKIxoQGapaVOwCEJMajNDc/sn2FdILHq2m6mBEx4m8o
3gkLe7RyWbHaJRAy20oTMiWGvFZNk/J6LWHrN6S/gJvL4A1pHNuq0OD4+Td1O8OQ
2lZJD4+yRgLCUM30YARlk1ip1xDii1rm0blPjqmj1I7k55hWH9R9kPzb7d+6sVFi
czp6nR05SmKVGTTb91/8xtVvi6H5uSHxqVgrUTdnhc4rV0yCJqCk2J0kwiTiupJX
HZQj2RkOXpjJTo7kPYG4J5tdpWQ4BvZet7pzqQATE6cSldVcI4T1fQGmgWAb0sOp
lZYJEeaELmk9yHcNA1HNGd+IqWh6vhFBO6rC7cAtr73OtgUnzBVHScScq05utuL5
wjLlyZTvKwpsr9LpL77QQQ==
`protect END_PROTECTED
