`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qb6mW6Q44RM+oCCSii6yoLvb325mipTYFsdt8nZAB8OAhxrexsQ98uJLcXWjV/C
p7Tnz0RfgI59UMk4e+rkh4gO0yArkjQA7ReuJ3SEHq8UeR2DILW+BAwqed59gEl7
J1Plg+76iPrt6m3e6pKsRVofMS1EExhFjNkvH/fX4v587ygfN3+4+1id4/ztmuRI
tW/Cqh2FcNqQ5diAzWdTo4uO79C4gadhiY5vWd5nHDbpPxHO7pZ/GgcVQ9Yp+Ody
0pykyfi7EwmyjGPiI/k1LNdCe3IJaajQTreoERs+kSrsGGhHRLW4O/umtpuJuUKJ
z+V/H6H0x0hgcO9xEYFQu8WDfuPCPg9cMaPbSVhP+8DaZLJSa5cKularjBjcTV49
pnw9lhr7JfVXhnSktC/dkfLK+6xKK0dgLI3lxsdnoBp0ZI0UcKFOlKlGjyNqkG/v
y3wjyfSwtt2huOJcw9oO0ostKoGUEejMmGSrWjzkd0UaDL9qZp1R7ch7gxVoEVmu
zqflbYwpGuyrSDzq6SpVXxJcNSfQUXuAgwO09D9q2PeaPQgrGeA5HNhaXaVLKbTM
EBFZAUB2svG8XOZuIiurrm39/8QzvrfEQ9elfjRfD05RGtCkZhpy00BPjlwjwaEE
Kt4jF7JvxMOekdVPndwO4bFUryGkNSk2C3uQYNgKj5iMxCbQRpoayL7s1qXotWEK
8Lyqjw8iAnFmpOPS8CjcnRtlCdhBoSF680LFeJi6q4k=
`protect END_PROTECTED
