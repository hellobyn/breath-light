`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccfkEX1TlB49TJuj+FqDF/ivYLlFIb0jwreb7D88U411mWp82n9Bq+Z3FjUDFe4U
/DGkxKOn/xa9pIUzElUCV7glPDmJFfW9OyHKtUqZuGo/dGf42Disp8rdvplZJx23
FLku3ycA3Jpo6s9rWZMoOP85+IDMBk21Hcjn3F/R98VCsuFajALBYNJjeyeZOXsz
OKvZZI16H1Rx+FJdJFVOzxRbfBrpXPAzME1X2/+lQoH7zkd1kzy0o31hObUxxWWe
X+b1SUHpXuDtUQlCkgtNgdWnJoKmzCl9QQd2OnL0z/y4It+/QQQQQrBpaeNF3bWY
FIk3xuXND43+Is5IHeyArvkNEHWgbkts3RJnNTwEfbKlejPBrGtPJR24TusA/Lrn
0X6oNZNyNtlzUrj2ZnBSYYSc+qf77u1dTuMMEpBK9/602ERPu0hrqCRiYE6Wu8Lk
hICBmFEGMkFyXNdJqBQ+qeX9v+hfTKDZq3wrKcE4UzfGTQUm9k/BsdSTHxsSj2NG
OKaL5ZjQtPrmqeFQaZgaXGQFNAwewjLvLXq+7IrGbjyuqcsBNpG0x5jVll9mQ0uA
z0jNbO//HYokIV9MxHmaUbbTBYqRJ6PZHB3OClcP55GFO9m/N4+L4uwqxPKGQfp+
N6FZs+S3A6TIyXZBq3A31neWv63t6jie65AnY3EzQ+DACxEtzVsD0X4kg2Itq7+r
SICc6bXIoQMYce5c+OgoIEtdaym7M7fLChLMmljipumBZPrnRLBi7K9BtBjoSR+f
m1D9j6iB5DY1bqK9tOL0w6virRIvzqmAqXGQlfc8EyJQSBw0AO3XXkRGk0zWyim5
oXXnEYXOAn8bNA0BMH74mosJ1pbPDOLs+wepN5c4Obk2kN3wbYrgP5gfaD0q+SMO
awJAMb0sUfbZBZLkXrJZwFKm7CJbCrKr93HYXVNNsnkRZMVT8z+l2X8WD/Da1svo
WmR3rw2A+HnIxm8JqMhCasbAvzvd/ipdAmS9RpwFRP6yvBzeSegOOe6kVwDdkMom
pSQB/btEKQplXXXrmI2TSGsYr9rDQfwl0AdAYb8CCmakQ4L2sM0wYcv6IQ463p6R
qPmiCE/WFwW2Q+q75Uh9JgfZHyKF73Ig8CONZK7aK5mw7plrbWRwtkhjL34tsZiG
Bx54U8ixSDo0Te4Xvg22C7pyx7sWcXJg5J/EpnbyX11Vfb4VRafI1nQmZzVL22Li
B+FG8umHIW6xCAzvE5pOX09vbT0zggJ5sNF4iEI855w=
`protect END_PROTECTED
