`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+/l4jpL1OKXBuWOQ3/K5Fk7uT5ZUZ5Iqez0SHDowokBMTtiP31CDJaRGTUweg/G
BWYEeDL+35bUtDbBQBTeXWtxsGwLa86HvPlQg58qdwdhuzOhzR9tfiSyPYQZnt0L
KrgDpp3KRxwJQM7IH+z9RbA/kG1iwMlpDPhLfDMx4IXYgv62V8I5NxTzsUvyeAvb
SJRZjeN9aiDqdp/T49wTTMTyx2hfkzR5wbdHMg03ol9rZvBqmkR/jsrDGj7T+3es
q9XXO+GbkNIXkY7aAQlEEQ6an+dMY5WXTeUpUQPiu2yUcJQlDTVlEPcRF914AY2q
y80tQgVB0WJ2yJ5wpGOg6N58Z8h8Xs4YXvhxOqHiGdQ66XeDq5X/tX2zs3z1d/nN
rTgIKzd7P96gWssE+FD9+LQHpHHRNsbYpRnbLUwHmmKa71JJvlzk+n13IskjVhYM
TYGsoZ2T8Z6lX5he8d77gAxF1syF4YU3Qc5ZlyHpGeOt36Z/EkxPtaaBgjmE/2EK
RvzsLK+H0jyUmpbxsbycLllWtIx4AqJ3Z3MogYLMTMCFDdYLmZfMyuRNpA/xYLcC
pW4GUGx04EWd6qPXhUHvnd9HjEwDrc7YeM3RQHynsdOYFJdAntgcHi6s0ZhquF21
t05yiTaCObtUNJTUdXb2ntGYM9wyNWILY91F0O6ueVaKuI/krRnOjFMovcQxwrU8
7yev/y3OiWOCJenqolP1kAD3ACmxyWLs8E4LOP6Vyq8CB1Z9AaDWs0mDw2COsXYs
ZLzk1xG6ob1VZeNc7FxTa5Gyj2YejdVHXHVrL2eiysXjH0Eq9KPKvqvzjSAa0Jvx
W6B0pJpgnWWQ3FcVnr9VwGyJ+9YmXHiTBVsIGmklyJO9xIEiRf8dZCOnww/12++i
H5SWMdGqr1CE+P2iLS36JmdnisG8nfhVkfr1Y5iba7g+F2zDtP/ZX+w75mALRDFa
2X7PBHWa8D217GbHF/13ZZWnbHGO0DDjD4jyjgoXP6t5Ti7DkWoyLf0HkM1xuT0x
+FJqLTZO5LHbzbi/y1g0HVxbPF1hn/nwrbmROtdarePpBrABghqg80p+lQXNmS/l
B+G55fvCCMkUKG2zAUXlI/27qasC2QSUVuM3RLhZt/qbVejrSOVx0+646djgrhdh
cw8fL0bNQ/KMse2HXtHZaXACEMbs3YvMPCmqdXAH0rHsf9q33cgCCJA2/CSS5+FZ
zkCj0Q07OWHVVXc/8F/oedNCLQdRUneEii21YKTteD/2UT/agKIJyd8688zgnbEf
Ko6pUgUSgU+76AGtXGKw4aNbqMi2N5FoiueCrQFNEo/7I2+H6favJogGtYitkFAN
N5o9S4aKKWeh7ypa3vmEjuzhM1uVmpqk4apFNMVtH0LGZYKe7EQL67MX4Koe/CVf
zgjXZ/J3fdtEuFIVqlO/OleUKXxGW6AxriDtGf6eTSkpmCkO+4kUEN2RrkCWalUL
2oMpM4qe7cnNysikh2pRtkpD2kam1eGaVZv7ekS27M1NOOLmJftSSYASF8gdGyh1
FcUZRV/TbiGos8o5yQjYOxQKLjxgM8g9gS4hZD4Y7/mPcgS+ek09fXJiEL34RdIL
8qrpIiYHrJWWfNLYk6I2Mex3qXrv3vSoo9np9RxPGi19+glVwjSjQWzTVs8Hx8bK
Hugw07/7Ns3WrItEZiY3ANkao51xBDPGCa50DEV60Hxf7yL4UNbWfYxMgNG2yFE6
pLpkMUV7lHjNehjUd73yWh+4hDPVeYNFFCmGZdfFqgvFub4xOtgeFZ0tQQwYbVIF
cMzyU9LCI9ok65f+BVBQl9KGWoN61MYi738Ejw0M2ou7+3EWiUQyd5ZYpqeiqpbs
96oQdrjgmbYkLFH+5wOA84bOW1b2roy/lQDZ6kWqo5Gqlr9znS2LXksXAXCK4Tj/
6xQ9I2yxAGlUKVtbbpRFc8k94Zy2zoJrv/UUfyfKgT4iOSzGazNMaoJ851p4jDXq
RSUiOmu9WDB5oz8K+qIvTkuBHLt5umpbU55raoyO1b12ei98KwDEYdQTPx7kmSAm
uz8u3z/9bdA+HqB2SGIAJfJkjKyffJGBGrVYZUuoFExy96oXzGDLgwoTop/FvII7
EIML4ylg14GmtAZo8caoHWVvcOAetzBHGKmD9OZiUQmJWe4EeapumFlUPLCBxa+P
rvly9QCHOGbPnBukuo25EZzxBObUeMyQMMwERQVIMeG1SnW5VQqyhebo2lOKia/o
9WpCyqMOWYYIVDJk1pFybcampwBi5Gkz0um1aim5YKiggRnKIZtlwY+1/dJfptyj
hnjOwXl+aXm9f3fYG7IlALBej9o7oVmhFw7C1+EQT3kcJ2CNPWaISAZV2JUOC66G
AmFtHrPmj2e0Piv4os8QpMS44nWVSvB0jcRufk50i5rZmBa8n6vgMmae2lyCR5vw
hykCJ3m6GKtjy09ByaX43Bo0VRhJ9ddq8rE/w42iER0MOYVoNl/HmEegOgQyw1Do
sdrUPgAnPC/NsjtDx+Pv3G6ikgWCiqTluJQ1Zsb+nqPPCKL749dK+LIRI/cTN7kS
dB6HLqrRAWWZwCOrhAS+S2U1hypgoRK946nSAPpKaXl4sW6UDp3MUV/icxiiLv81
e1kpOMndyGIsu+cWVSrqJzYtRM4Cf/r9HVpff9+IHsXuDbPlRXVB5KUSDk6w8gpE
5Qx497d0BsUvHAwIkF/krgMCsVu5EKaQhnBW8BoWQu5TYrD2p5Uk2ZXrrEQqEMVI
LrnsBjOhZvryfT4QYIXGXh//wKUTl6yLjp7u/BXvH+YdnNRQ4VYEPslXPo4NihhD
6K26ot3zxIs5zCLbfkhXXBjLKp6FEMCLF5eKa7mlb7OisbAC2suVCk4zaYxSBXAD
KI6wJddwVrzTFwZA0xiI/rnd8553AGk5AEj7JDo0lhpFLKr+Aso450kM7T0NAESg
ZaeZ2vQsocDG4rV00UVjrJdAscn3ny1OOVZ2szxuvIdWt3WlnF+YzhQjc2SQjJm+
JFPf0A23MCI8vcY5zXv7VWzFmIzPzI9vkwVNm5xddfP1RVU2nNqwHs4a4jurNDAL
HJH4KbRNUZ3Z6jlUYNbAuu3dg3/3QoLYBUScfe+o1eKTa5eqt2UksqKOGmUliDMj
2Ceukvx+IWBnYKAo3pYX+M3ccyIRluOBKmMgPbt0aKffsQTupndTOTXLkctrmRvw
NkRr4e1g/bpxxUggZFTZEtrORWwOmkNr0Gdue19GabBlYMCsvBJgkwrj7FtX2dN1
GZGtT7e/bs3zTpvfHsdaPCjGGEGUKZV+tD6tPa76d7Uv55xC5YbesogzQdJv43T9
HvbYKd4iSjLNRSBjCByx6Sxg7+v37PYX5gOI7duEdai8rQbBVYx5OkMD1vq4VpiR
eYVtQUEONrYNuCg+/Ay8meYTh0qhBKxhLwAT0gr7Xdkm0qYVrS7ks8WzWnpxxqrd
6Qei/QQGS0qjbszmsj4UYXDOnqppbzKJ7kW4tyd7uyEP4AfXVbvvznk7ZH+2EuLg
XJ8RNi5F1NcZlABpy+ho7ZOaAx/F1NmWk0q0AcOQ6Pb+Oqvg3ArkRWBbJ8y9ZdD0
gDtfv4YvuIvdQDKaJ3uwqsr0lE19Hv6OhYvJ+5OJwMvwb18JvTCGrGKojyXoa9BJ
ODBabYEwuQ3UQw8ps+QhMDyVU6MS5MlRO5WoYY4CLVw+sEdBVY+NXGj16hHJpmik
APlZnph0O+rDwO7LdhlwF1cw6NVMrDmQ3HzKZw1CKXCYsyiK0+qUa85nX+Ne+lun
8XRv0oO4uEzOHx0Kiscysh/epERugLVx4tKTDxA77XQaScHaEk4CZX02DZeD4OLV
VltDmbuNvHxF4UepH417ng==
`protect END_PROTECTED
