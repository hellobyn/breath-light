`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vOKN9FevBABNweLWaMcOyZnQoJxGIFIXwzhB32Gh5RWKOiu09jqWPt8wyOcHIcz
3Ref+xOnhEECbnr3zo0XRDtJNHrg7H1WiypRDXqZUYiLu5Ics7eu+9OvvfsaMXIC
HdmfWey3MgykqE/OLQL3r3+jmDd/6qb0leRSrvA8tPpzzQgTfO2Jb+qpyb/rKBYr
mwLjwlo0S8izjpS3uYMMoZsPyN9GZUvbDPHdYDomG16bp/qnWUWuHG2uppnnfKx3
UEH04uK5wTxeENHJkh+ZMotIGlYxGeJ8+RlpLfsLfCM0b0i57M4e0+P1ROwzdH2J
oBrEB/8SO4z3ZclDipFU4lkULObuyLnVib6llW95jZuNWZwCkdTIPrZ/iYVmw3KL
MpGL8GrFcMmdnnk7QKKrsGNRsjRxZXbI9oKbYCaRwuzAwd+r2O9UbbdQi398TG10
HQ4AsBfuV6j/jr+96TZyUUIEZe5eRXSl7FiY3ejL0KL1CbdIfEf78EtFy45d4QzX
Eq38bx+mIzBnCpqOV+/QQhLMgFAkAcyfUGGKdKPP3ZZactvSCouPmKM19Qse3+bP
W5P8zpUTZi80CC/kTsjqIAI56JreOfqqL8xrsh6vwjoMUNDcxtixJ0fBp7EnvTx8
I4RGGLHPxa/SYmLey+M2SsKg9CusoUyfrsG+RbwSKbh0uQQYELlIxW2X55lxSY4J
K2Jps/IXZmu72PnWCqo4HMYrod8ccukHRMQSQoiAlWL3nDDM+TKEnZEqzxHSi7vp
r/x3lDcwxhcop1rKbNgNUWM7HvRSt8bixg5dSQjWIHlBwBYD4bDcDDqYzt/SmcqB
xOgOPSUgcxfV2oqhLHE2DwHSw+8YamhFr+UNy9g/23NEbZFAx5upqZh3WWqvlFDq
rDKhOdqOBVtSXDnP1yAttBm8VC21LBEr1luj0is5/RVd+/W5Vr+2CJzFsTjPBRjz
4wzE2+kkZHd1NC1vN0XI3P32ZLQWzLVGMWYVLDUOwobVKXF33iXUsezh+AKF53RJ
pkE/6Cdp/tz5yK/m9OEUobkwYPqL8u0MS85Kw3+oxRnwQBmrV1giXH6KvqB5Hz7i
15Ixm7tWS8Xq475CsSTyz/8SHSaDaAqdk14hVAC6JRCWURKSUHags7ac2LJ/3MAq
ekMXln7TAi4gGHFokg74/OSY2hU+W0I8iAbbXwrh7VVFvQJD0ru9CiRFY1mO6bEt
JRMBG+STNknIKpqZ/QVrexnNY42GWnZGsEyRD9rbf7XhANA12e69jQbJiIakVET8
beT8bCt6tyeU4J2sH19EYaXvYDszJfaPMWdcRM+VpRhdGBlU1PpJarFfEwRt7n75
xsb4xdFfd+AtTuTn6H7pJ0URwzzrG1ZviSYdf3tN05+ec8DeGWV5iq/VOSdxKPEo
wULmbBwEXowStJWuxYOr6MMndN6KhuSue2el4ZgTuTbmGAreXxJqGFUrRYVQUBmF
PuwL3Ef01ja67FWLq6kUS79LTczvGlCnDu0J3opKgavoJHPUKdaUMgex1nDmEA+M
WrLHGCzQXyU4MklrRFrWpp+2s/Dn+zQi7r9CyX21aJsoDVP60UxV6cSSTDHFOCcj
QIEiNMShRujiPHaG+RKP55wNjdyOoXqDU+gZcRt05WUrNA/Aum/eTOWPjI1eHSOh
UqCKBD4SmCnju+IIDuRl029wzOf53vOAC/wcp6VPfWsVSuBVQkMD1/ac9jGmURyP
soN21LgnXj32FpJnXnWBMYZTrOxneIQd4hIQGtbqj4NpWmuvSxyxe+Uqhhg3qtxm
MGo9QZHoMZ8A3RxWRYK1A3f0+YGT3yNUNXOip+jvQ6aGlgOQGMLBqSKJPNAmtjAB
GibBwbaBVJLerjvDgCJmq5QqwAtZ0os3vTxX/PNPEE3QujcJb8xhTF1zIAtCPVHY
xV+WiBWL82Uj0QG0Cap/teOsYwjgTv2ritC4q0WGvuaBv7v+wdh54MNIi5HsSn0U
A+wNa8fMCgW28ffJ4M6++yKZuSNM4+XptD0M1JMJ7c7KuCCQ8k5UpBwb4H89w7B2
KjBfLushHr7Bbc7zbj3VZ+OBr9uo6y9h5YgKYD7e8YBJumGMvNm2l1lbMepjF5r6
TNMrD3haDsVt6i6SVVw4qBykg13BAFpLG6u6duND7UozOec4BuGEzuJJMERIqiif
kuwZ23+Y1/JCsx0uQYMhuEVI6gLciOMlAcPEVsdS2V3UgiWc7Blzy2W9Qw8xXxgZ
JKfBrP3TMGgQFmfB2FA2gNqDUaTJSNzdO/x49Hm8u16K2VTCRYvSLPdHqn70i/YQ
1DFlDEXOr3H1zDrzDQfyJFwp/3O5vS20pb22a0Z/p5SJTmPQARcQz25HSVnAZe6g
CsmCK42oUWvHere1b8G/jnPl1KCOLtYhHoTVi7GLDDgy58pC9tCBUSURqm5X1L8a
TyQrjRpN37i6SXi9yRkLRw==
`protect END_PROTECTED
