`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhq1QFZlhcrgomlH94/Y+vKg99Wvy14HjDL/8kVSxF366iEOv9YQ7YatbQ6QT1X/
XkhSFndol2EtEi7p5+WYMClXuqvQ6ueJo0oKhhthxHGwytPYS8oswrALXmMrAPkQ
UGDJvCHWf/YyJ+ajqM4awP5Gg3MOXI0llng4xXWutTT2cVD4ULj1sVHWCZ3Q4GVH
/nU5oXfO4/3nBX6iOIrZ8lPvI6AGl2edroeMXH1Q7I/v/1zJ9iIRHL3aqH5HiE8x
tMBAConBQoZXXPqAk0pceWm+xuR8RGlVNuA/xnxQ3hSvr1PxgiyEwHkj7olPvgtZ
Es0b2hCSJh7aTaafMD82T5HrcmAl/1fok7sG1ZmH8vddXcpxkseCwT0M6df9a/iA
nuKMZjFmx9uW67GgmFAPSuM94/JB0ASAVYh4lrlPOJod2kf82zjFhTWMGk9COPLe
LmXLGsP2oVYrWi44kklSui71EoDN06pjve/pBsGXI6mkKIAn8xLpQgg6+mIZo38r
3tv0Ne7CpRtQMMZPiDvgo+c6kpV5sH212uXy1Le2jMIP+Y/6ucJok1Q2B3Yt99LC
F2HaoKexeEHAB/Xg6LZ49nlFCrbUm44L5Dde7uW5BQ7c7KcQ5c2TA/jyK5Gy/vtx
9WsL4J24YAGMEh5WWKpytdbZ4SxJ947t1CfnolD8A/L30z2DI4px7ww7TqJxZlq1
XZ4RPL4t47lZb/7eIOpLj7VCJ6bw6CS+lEtPfaqucHsWtDQJ9xOpsufWqxh3qPkq
V87YnRwitErGQ+x6aEib5u1yfqXZ5mSZ1cPfRbjbPWD5bD9/uE1mX0ykJNiuTxXU
RdkUN5tkux9sDvR9b2S66sJiRw/LboaaaoMWLyp5AYSeZixttUo6lVGAlGSPvlW+
0XB9GQLgItCvP6lRQZOyRRNkzE7pnA43JaTMtTxprs/9nJpwdSkM85MrBmp2sBDs
zjngkB94gbU45NP5WLP6Z29NxHdgifcQqGX0yjOhIctdGFaVHqDA+V6sw1qScJ2K
NMfMPKXcU5VMZS0EjwHr/500VI707aDYnyxvQ87QcISh5BVyCFJcodDdvlN2qUpA
Gq2dnNvKXvv0n3weoLWA7xFJJigoRg1RFDvYysI6qJl8F8dv7xlycdmaeKa/Ip37
ejaSSOG5uKqSN+Ztw2Y5okY+i0XRvwoAv7XX/KcSNxxHNnkLfh4JW2Tpt8VEONw2
KS2SzwL4lEV5uWvXrIv5VcE60ztUZ8xyNZie/d6BB8cx5muD+hjt3Q2zVYXJMJkL
bvMvpbb2mvvSVhSQ0r/G5Pu3ubwtoBercelY7W1tRFeHVQUPhXVNJFCybRBvfKN0
zqVzagMdw7nqwToL0G2RlLru1NfkQJKCjqpkeCt1wZXi7+BH3OI+pR7ylndi9iHN
4dUh6frM5g1X1WBBwF3OksCZ7EUX2h5//cQD6wNFL6u30Gb9u+X2E9Ievoao6mxV
krvAqdxwcmr2WMV9F0uo5nO53W+scenNrAIOlgDG5CSXj/JQmR7uKKFthgcMEiBf
TLMdxmnaEPPFKXcIV6Sai/8iKmuZbNjSBlQpj1y/nsKxIdaFwhBTLNFiWxMAWbxp
KT0PMIYUE087zckpOzYOdZiw2EJd7HUtSjfxIQ+T6wSwp1+Gg2t65+aYzgg8zqXL
amEZoxyVatSzwxK5JUyEno9Fp7daIn9lBLJG79F6goG87+ci9rETiiogN2qfmaIS
0CGlfJzycSXwibiQXSbj8caAMDQPrGqGExB7O3cGhS1rB2JX20PxJKkYYzJqO8pi
Uhq8eSerPeC/H4we1DiQr1xoMgchN9UujUsjPjzmGcelkmMYMQtOT2x+/g9WsV1b
L08BmeBsWsj9Wtls3HAs2Ibp0qllcp8CICEjpoNmh06pzEPWGtwuaZGYejrxmMsP
TUGY+bXY5z2u/7rVPD74/RTBoKOFdNl1l+3GwMBTXjOrIAJIrWj3f/+2j715aQf/
zC74tipfTYHl0JT5E/iq2DFHcsodeX2Sgt0V/9mz5d/YeEqbQSxRbVHaTTT6vVT/
j+Cf9uJI1VxuAW+86NxM5rYwOU/M5CqtUVPPAH68mQR903HYOkg1a1ATQo4Z5qSI
ianqGKw2bLUyAqMSxiK3DaQIaskrR3KCIKqZkc6kCQRcTjS/uww6IxlK+DY/6gv+
2WqbQqIZGu80kn1Cjm++I7yE7l5ljXiljIcPZm07DPdMi+HoMQ8KPPiOGODTEF3e
Uh1mZH9TNRW1Rf8EvMVeOgDzOuX/Oz8jXQxk8BTbmyMIRubtZpqPvPo6+8CXS7Do
/tlVAQPEhkK9a/XNsclVgQxTiJVF1PnfWcVY2iyNyAG1wGs5FxaZ4DGvlk5DRmBJ
y5Sa59eTlQHGFfJi4wlqP7JelOlG8x9svpEWX/hzD75pildJcULakV51SXHGtIQl
jnNV+AIYTm6FH1H9rbjik8YB0IRKbS1jSeN6VlXH7OLLPjilmj9OQcby3sCzCtBp
/TwksRV8ZC2MyOnIF+mCByzBfKcu4u39bEzVHn4oFsG0ihmEnx48Y65wNQZlcubi
UpolHEKsAFtsjmG1awwEvUpJhBqTHVntqjnUwpZSXZ1f0TM41BlmZTJa2oJaqdRq
mgk8dgsZ1o/tj9l+prg2GBnTkl+YyQ0bzqgQunQ0uFL9Ky2A4RXL4HTF5Kw4JnUF
`protect END_PROTECTED
