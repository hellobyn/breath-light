`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJdSqPTZBacQ9aN+q5EPxu94vrxneCNHy3fkEGSfkQR2h1K460Z/79mUp2/eF2Or
f/Ma9AWvq5qk4wZLdF7ibQ+OCJxyu3EeyNPKFuXIJIRrK0MCx5n9ufWsnccqjcRH
0XDvm1XsjrfUQQwp+dgCZ/og9um/SFpWzqqKadJpeRiORM+yAbDkTBfzzyT//INB
++VEVUBjdCAnpcxemyn+E2aGs41/DjlTHsneep0s92FbZvKoc7xjt+cYajB0IMUB
lEWT3xrlUKsK+2M5AaDygw0hoHyZc34+EuBeWI96ta7eZI40qxbnExrTRVvPYNxH
aLdDnB83pT3MgsARzX6fi/Az2pg8qEpnY4vtzdECqnL462X527rTNU3N++hix+XR
+YCKelrsHrveX0ZJg6UAaDMN325sf18BMwqg8Ou3SDB3E1ziwlN9aOjLwmLtlKlq
/EB7B6JWYDgzbaV1NiIbsnd2eLjzwfJbcw5NYCTU3X2LocF6y/XPhcI1n4JafvSi
kT19KLN9YUdfyPkb0mnV5+axIVfiHg01Ydpv8QVHtv9XpN3Lsp+yzd9x2g9qR7eu
cC31hp6zGoGcR2X4MrQNf5IoYfHTmMpv/YRX0PxTo4m9R8Asm+Voq+V7CJiqGoTP
F1i/YS1HFDW4HqtEkzHs+5F5wA/iYA0Mi1Z1hDFoT2PnjyMo5mLw+Bb9Nd06hJtd
zsY/mg+pOZK2/Xbh2tBFxIFMqwmGgkDHTO6JqYe6rHWHRHnLD8Ks1jBOqZzhW48F
rBxnfz7+rfRU6A+4KPnkhWPHf4UrtoCR3HMQ2LE9mR9Lv92rZWOVZvbjPfn4jhjw
/G0oiTkG7XRF8YZVlFGM3kO3dY63NVYIjRdcfK9bIGmF7yIA2eKZiovEljtdw2qE
E/A6L9Kw23JSUM11FZGxtlTeBmzgSYAzVuC5nIW3MlD3zl2BfUnJpYwqkc2ga8uq
17gRz8uVs1a3sDmGvXTN6UIMHghLcfGA4+NBo7nKWfd8LMPWGj3ugghyun2gHGkp
qStU++ZmNpSvfm2QI1T0b6tlk6ioaLacFeSbXqI6NNCE8maO/E5xtpKPPxk3rCgX
+XXaURs/34xn6t8zFhFtgvLQy+lCBTKSX3BEkT6vFr0rNvA0uM03il4aQiBchQyi
7mWFQvby3Oc34V1wl35RWsADuNdKhfY7L2EQLL4K7AFr7gMB0PxT2A5a9IH8Mp7j
4ZJUHL8Z6NbqceJoOd2CTVUHTHMkfDzsluDBlIhgKQx0f5tT5AG0hahmBtt/lbZL
WVfKQshiZpPdilSYqVxV8ei7hyt8/twUpJ7apnobVOa5sVbLwWCtUu0pXnZjfJme
C2WeAMNnEYZ4hFyYul+K70VXjMC/les1ODa0FkcfXnlDSN7weSf7rvQcK/kQ3j9z
LSkZ8z/mIqUujln8VEW45yAe+t/Pfa4F8oRlLkn3Ar5Hwo/OltDeUNfK5Fn04mcw
aoAbC7xSff2EUxiPmCCd2GYjYx8RZpFddK1XzKS6/hcsrRAL2Z5M4QD3uds29TFs
JaS0itnQg6LrriIPUnTC8jW9Qs2OEG7TVe1KPRkqytD3PC0uKsNw0yTmFirEetdE
AQk0v99HZPkLLZ7JWrrL9GkKU2Gwa1O6HfD7OXNPGozM++DaW2M5KJhEBLzYTh/C
mdULvGYaHDLGWK5Qy6amIpnZU24HBW422L2EhmbrTyUrlHk47RYXOm7GCU8RqsgF
jLTF38FAb0nQmZEK7LSMHzh810caCfwxXpkf3n1jj6Oz+y+uolozF9epucSKhqCW
f80VmIiA+ye+IwVKC8UH9ROg2oQflzRns8tgrBYcNHzxCoahxeSxgeDDZ25nStVR
njy/n/DKQdGGIs5V4KUeGUedHJk1Y4y4rL9DcshBRKlg/H+EfZAdFZL1HFB00D/t
Cms0Be/zowoLh3d1FMm3GnQeoTA/LsqPnYXhcC03o1x2sb9IW3diQklzNEtg/mUD
xjetYp5T9itMHGxDRBik3b4KUSmlA9riNQ9F+nyGurA3fFQIw4Pq/PstMoVgLchc
KchKj361B65IaktCME4j+D+WG9Ahilb0On8f3NgOuxlqGjHTOtF04g4M7elmi8od
XdUuDkvVFU+f0VxGkOYZpxev7EFD3DAl6df7xJcMICiRaa035cQcZi6AnE/watOb
08+N5LbjBrYZuw7yhgVapUMICX+S/qJ1h7DpMxD3rCa+EkPk665TMV2vmDXLMw2y
D+73PiUYTHVP9SCV1dqNJTNgZP0LAFaWn2xOjdcavd9ck9TSd9GIExP0KFTN7bCB
xxjyK/wOoi7Zbr3XAJphCNiStFwjBrZALymH+ZqYAlM1xMLfL4G/n7RByYZ3oQbK
0iouVxl4lk6GG7tezuMkLA0mXzCxTf8UCZUHUD7OTWAd4oiqX4FwaTYvyiPpmzll
9goyNIvi9R93VNRiab6CLom4ANIGOTOUeH3by0fmRTfRKv+qoxqyHtEisWpHdadL
CBtlFheJlcOGOMrO4d1jzgNCCTo1z3/nb1sp8JXcU40Vw/d8Uuep+556EYXPxVzu
0WW8fdO+Zg6vi0fTU47UOn27/pRhzv02QJHnKkUUW7Wry/VxzocwZ/pHXKl0JIas
jhnPDktEiNleUAm0s1O0E5xhkjOfwwM7EQn45fKZheZjB7DkWBZywqcqskyteeh6
7DIVLjwMVsKoGRBbXzI3Gi8KYssslKHFXPvTWVl8bfnL88mfuV+O6vxpqbP1aIdW
OItx0duvO5x/NTzxPZh5NOrnwOzHNoaZ8EYLlN0iUO11w0HHx0XRTo6gAb5Ylo45
KcTsIRIvQwd4Rqr/B+7Skjk+ipAO6My83NWa07Bket2mo0bh2/R5PYoXwR9KoFiw
kR6h9b1rPpS1197UlzKwOCLYU1JU4RPpa7+fhetVzbE=
`protect END_PROTECTED
