`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IF/+3hcfh40KQwZAe0JbxigRqhIL0pgE6viZVQVS4vYrGNr3+BcXTThBAO5IJC3E
MjPvrRyJK6Ux5qhFhhvIFqTqRJQemgnU0RFlrFBl9TOxrrmYx+lssloYhoJFLgEm
HkRzM5KEh/mkD0CZiqICmN6XWMUachYgSXKIABKOUV6XTbdDjpwli99l5rALtitU
djz59eD5ZnpKOyjW+mZMfFXO5YtuJoXJeU0byTRB00IrmbgN8JQruIcwtGqX9JtX
ATxDMLuo7WV9kKJVTiexkRqNcwdQxWJZ2bXFjymx3BRaVUHn+e7DIqmrly2jgxus
cofjOvRYvGg06W5PTP5E7hf1zRY83we8zBmbVpJtKD5ZgNLPXWn7sZfhzALT8yZk
hBcUgmau+hjsdGY2fEN40O+qmCJgZMSyJcCfz3eEjugGCbaI+JpJYNbO/Y5ZntGk
TKWHcxDAnV4vwOp+u8nJifepc4xPP4FsKarvbrP9JqHqpcUfsxwRCr9bPDvBgEss
o/C7Z1WDAVfxqjde6+dTG7OJ+jRhyM7vMOzQCN1UI6V3h+n5sXNtOjLHfD+aK/Gu
KXM4xgE/g8/6WZqeKYZCryG1W/T46WeeMkLLyGxqcYQt4j2BK07WdIQ+eLcsnpZs
IO6G9OGRtFUWGRic15M9saWLT4cG186UFDRygG7fhlYa6yinEql1U4ELcX9l+Z+D
X5FaBRa0vzBnf2+ApYhCrAHiZUiNauEeveB8oNOc3SeTYTL64yjUtVBR54u2k2al
v+Q/X8Jy5bfamNPtfgBMJRyMe0oTeZIg8BYi+HaxESZL0iQ/eexxgfESycV6pTFp
UsaGXxAN3zgATJa+YahxntXkEdVzX2TWYv5/Z8tFMd6jVWO4afYXzNOyxU8w35hg
x3gItZnaCj/0yQJn+nIuOnHTHc7cPx7/7cAi1NLBSDTyi3ui1+rRa/LB9ObGRkXh
9ko9yPFwujcae+U6eFUt/BmQozIc1gm+CiD3HqJ5+/Z6uqZoKIiN1J4doEQ0iIhQ
RyfZSIbIT1qUk1XQ8p6DuZ3nPlwbCemmAilloAFe/cdJ4V0rWtS8MOxNo2Rq5x9w
F3O+xNRFJtLKun4w4M9LWmJOy1qoEZHSABE5lSe6rb34ZPjIJOjdiRVPomyS/J0o
N/ljJkci///i323IyM3lFI1Xczj97b3HoQZRqlAC+DbeVlEj7FdmVNOxO+7WbmsX
SucN1GdZIfIdm8Xqh7M9lq3DprfR6dGfStBH2IDeFcDAxKpuQXYjkbNc42h2QhX1
2jrdbe8rF0+0/ePm4lGEZdAoAvIug4IKFmHLxNv9MP/Ql+jXXStwplThe0z1SS4Q
DpyuMGS7TUjZh4mbaFeNrOaEGh3xrGVWT0HMQRfT/Y2bJNtP11ysQXE0eWBa9Qez
nwJ2gfB8WJN7vla5U6OO2L43jPVF8hrXE9bpmOasQ/psKdYzcawj395NRToWVV8D
Q9rj0g6g2ZOSCDTG6ThGM09xm9aijrJ1AkLCylWD4+TgM2R4ne5zWUboQoGJCo2M
gO/p0r9lIgYfWMHBuo30XxoLMBxqDvCVftZO2E13pD3jDekXoBnGdlYigsJJrUZL
tGdf6yxu0yPfTVM0TmdBf/Xx+TAf5kTes8JD2MaUkvi9TAyNbFB95WyvcfjeIaB3
Fe7Rx7RwfhVu5NXkHN6geBSe7IVttP9u4WboXbFnPwuXmITdtbO8Al14iwuIUtZX
KOFquY7Mc/Js+rmF03YyShLVr9DzEi7QptltP55K126Ax9pMU8OZ+CMYysNOBtwV
qqaauFrxXlC3RGPodnvdcJVEKsj18g9IsfP6/82b9xwsUj3ybp2z1Ox+htdoD3cY
rxoWWCmVWxHHjag2xuJTDeMSAfC0YVIY1MmQfHxTpIgeVF1LdP4G7Qi6ADm0HwBb
FIgsTLccqqqav0389ahTiPj5rin0sEpgm8BIkzpRxu3jYcYJs/XaNty7KDzL+g9D
hxMJCBA2W2pJt3Dam8DC9+9XCN8uJLv3/TSTm1sJK+Q/W8otb3N8eSRI5sVS3AzM
W2MK/LlJmt1dmNm13P0dCpNfvC+89G7XOKwr1BiCfdsZI7P+N3cRY8qBsycMyIrF
YfCmnZ66+9h3gs8HuqhDUQveDblkRhuWOYPsYgfY3Iw20HlAZzRgogE62VKMwkxP
1gPdLfD4sBwuTi+9mYksyT6FDf0mpCQdI5xmGJ9Uv2vnfod0OcmSYknD8mDWnp0e
X+ldEIyB70gYP665LLux0Epi+4bhMoZtfX9LRvnWXlWq9yonZBbPhvcQFBXtEqyM
m/yYPHwbWse5RWsaSjs738aFjZG40PhhUgx687Iwq2UKg5o1lXKmSyXVMwu7i/Rs
yeoWMSQWV5sTODEsoSRlqRDFcnNuUJM0439ugm3ama8EZej9rrcD1xfcOUst27A0
uoQdMs9oaKRNGc+DKrRsZJ145gQMyTqM4pT9MlMhuxC/jQ0/UUJUKaqpsPk7bCO/
Oo0viRcbT7R2O1mTuNF2NaGSRMvGLpd7KPJw4z8Y37Iu8zPmippV9peI6wfFxcnx
dm5KTth+ALmiKhCMdCNcUWbtqcTSl4xyYy2gKIHqe1xJL22VZP75+LYvbyFCZG5r
Tx1OZLS4NjGHPSi7Xna4pf9gJHcJTfBMAtiZKUEtkDUX9PM5sZFkpHVz2aTcNEBM
jkdfwNddCfq308ZV85jdelptheAIS092A+y4UPxMBPct/LGn+Q1bI0h3fXloTJbL
wBHzLwMc3uZXdC32u/AAhz+QzjNPPS4MW6lnigdqJhS+8PmKqF/yJU9UukKmH/u8
zcVJi0blQelex6WpOHIQGNJid/mydx6XX+JqyTg/po7oz3fUpOXoLyyBZtK23HcY
poeSR03jWUxszYiGWBq3WI5G9D9HLv4VNwnMld/Togxj7clLRvEmGqfSTQg73BXt
ijvZCyyGNcoFEB0jiaD9+RfHMrmWKsayKYE5W/MIjiVZUr+83VaxJY/iwzREDCYB
iwMtusI+jUypDZa01uHxjrdyJtgIZZvIr9WI9varhv+8Cv8DR+HU86dKvHuDWsvL
PPYGJ4Yc0TsC/rOADVMzuUAUmBGrWleFW6Kx7HdSTfE+QdUtZHevXo8Oaa7IpNHF
jOoNgnv9c6jUpWy6DVYEj8k1gHBBbyid2gVRynOlr2sVeEu+ee5U3KzT1LAAvEMF
DGBWTbp6d6l8tTRz7ugzBWgE5sNCVMGfumIiEJ6nuJ0kg1cOviQ2yC0xFba1BK5N
yQoUowIEdlJWcIiDQOMbPRwU8Cz99quo1+P3Cl4aAYehUt0xMVdnjR8V3LQPdk4x
doKzUT6/zZm7m7z9xz99rLdCEGGRnbp1D6uNPPoCpGM=
`protect END_PROTECTED
