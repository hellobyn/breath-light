`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMnVEHdd/13l1TXLjWehB11g4xOpQdoKkabysxHkNL0oLk1B1d3ZXmT9FavqzOqa
Cfr93RjJUfaqC5+p2IfPybyiFx333bIGAaO9e1K5hwrZ7qVF7j9oEKbTmo//JoCZ
MjO7U+nGS1iKXfkXyc1kx6R6ILFBzQtX2mNv1e64NSz9W/JtTo1Q9eJI4ZBh7hc9
nlb+s0HcPORUju8bfn4uB8tDwkhYHhjWLbxwY3/eKVKFfRWNt6UnWi3Vri8Pzjc5
7Kf+1UZ73Enh1XTAV9hSIQOlpdXvLDaehI/EV0ezWOUMDpWq+Q3x40+w02kIKrjN
qvOqa0pQ7LhOGOOfxttCCn7gxTzExpZsjpPp1aK4h4DA2YnPWphL39W1+Pe+5GLF
fQ6Be2gBoaH5FT0BjkNyrVtAQGyZTpi+N1mmDSqqIUswcbgZMiBFZHyJisXkuKtf
4Wd+qbyszyrPgXHsoR8IyyiwSW82jeBY5d8k/Farcv5kC+BIoacwbs446SUFGzyk
TsT8YO7cfasMwmOyAtOvwRiIn0WGx+fICMuZakZqdsu27Bzv98wD4yopcChSLOxV
zNuwwy+WaZyT5nhteCFUM7Mm/DTUpc8h+lEhgS6M61fXNt9frk/0aFigGUVXp1Wf
KV+yiXPfGrjzko1R7H5pd2qR4MNUjeSQnQKSetBwt/8jBt1pfJC0qWKjDlxPFXqW
DKwSIrBr+0dpybA4EIJKmeNUtdnNi/lWPQW3L23BPfEeQjAOXNIoc2pcF/0nkyKp
3OAgvvPzKZTKBxW8CFptEqQ4YYL+w8yP/T5iQnmxW9mByJjniK9QRYPob+z+OoKD
y2+7mKgMhYmusMvP2GTZ3ql9i09SkKDyhsIqiPFrsXvsR7Kvm5mkh8COdHYSSAvy
DQYAlgSZZvWhP2YySAyra5bGvada8VNUqsCg0QF3GT8S7tC51AaKgqgQvYuXaVXA
fOECZtKkBsK7oU93XUIu2HYLdN+YrFgeLxcnX96rUMnVtvwiKO93u36yXFqZVm7Y
TjrQKOvmRy6jInryEQMLOvWApy5lFesfgPwuzXvhwpGQ0eVBpqHzY0/bRd2yK3Sn
upzoGYyVndnv/tCl0QQQpTOwiJqADGirntJY8am/cW51ojHncXq58JBbEhoKL6ep
N7pT9vW0SI7QCr/Wshe84BpsEVkkHXxH8c2SZp9TonA7xa5lZPTgR/1MBB37joAc
SdII6sK5LGkTJ5uNjtNQKMGQEcZWvO0yvuFALabfOfc4BTAhPrCHtN8PfEllstD/
22Te9R88rLKyKcZ7WyY1Q0LSbRZ1ecqD7kuamGQoGjauvYJ3CyF1zheQCi020DJV
zUsqLq2mS2emUbaNlzhKf9SRSVmamLNFQbLw9S6T5TEo0uXLZzSMVVrFdI3mrvmQ
MPT2SW95x7Ip96/yvoykWw==
`protect END_PROTECTED
