`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGL6ddGQF8H1tMPo5ks58jpf53kJpehLa06TnSrH/t8oiB6sgW4Y71tIv37CROrL
8ux0rKGfKKnhfanhlin6vJGfxpy7JH6AKyX4ql9X8sojlfAmq4lw/gQ1TTtS72WX
xB6Mckn0etiiXxtRVVnmgK6uiuxaBL/InjUa1EEunp/c79ea+ANwxx/4y3fZjIL1
GPAmO4GImWuTZNzgJGrL4e3s+4063yOS2zCbWVLusJBMoNxURTcbTAL04UkQJC1b
nWDVeStXlkDggUePTx6mXuiWWT9xJE6G8TFpxXo6zxG2daY3xT9qTLTepJo8bWIu
m3Ll+f8kQ+Y4ehD9PQr/p/LiKdwstXRGTNf0vjXuy2BPCDqbM2ysAm+QvF++VJfZ
cxsEU5eyaDa+4E1dhe+e4Qma6jhtoW//qhNjTAteQPV/im8PqkxZo12E5ofBCKoY
l87pQg1dm4926fCcXMlb/UzrcQgXYqo3qMjgzBLrNEyUV9QJn3WyefdFMyNlITvp
qA7Z9gpIXpHS2LSB7WeGPJnR3M2X2VJQ5BJkhTXypyjnuF5Mt48ls95w7NlMo7PW
JX2Q4MKIMhVxFVCDlleuxL2YDNxGCQSm8WKSIxxT1uDFSepTGlTVxwKTNYrpTms4
8Wo8O4lB7d7QAYpax8fd1tr10bmVF81gnzUPzOBP4TAjCp2aRcwk3umQ6XoKsTWM
STC7VZXeerpO810Fr4Xjq7kEMEAPCkA7jynntJnKKkcpk2wstyCFIQAFtJzoD5GJ
j8VnCAmSC3fkurO9df/QH6eDqInpRFqjLissrO96/4m9LsaGFjXCjTVv6TtccYwN
+7X6dFuZr6k8jx5y9v0kAMpykPuUV3IzfbuhxHmI9eSoyiYrXEc3ybaYWAkfIbmL
JDGIp78OgzJ/qKKPd6Xtbwkh093oKp1htbuR+0g2vTBEiSpWk5bDaJiSIZ8iwvYc
sYX8q+FMFmcjMDhaj7y84NDoReFLxAp29ZHN93Hk37xKFtJSajblP7U/QHKSfzqE
b78/Wo4pa2rfhlALeOdJPVKVXJJE5jEh9W0f0+w78Z7HGSAzXAm2IO5zNN7ktwOi
udt0DpOlTfWAR5FKhRm8FLNc7tCrPyDyAdIE8emaaqE6g5n0naLhKGvBCSywQMAl
ZOedSubIyRmibc9pF/qkEI4hP18vx7IefVFAoXu1lMa/dpsNPYC92FUkqB5qAnor
qm8MdlifWSDf2mZRDlEJH4EbCn1bk4SRCk9SL0km1/IKlkpA+7umEH7ZK2JZVqjK
auw6IcwrMAN076Y0SlTXcaLixG+oJEPZ4brcVQH9Z+2LymPWvLXQdyc5KQs4FNOR
riolCnW3IE1HmKf9xdMyrIOzF6wIuVaGYeu0dY8B1jQ+dq1nTTZdo/vtWfr9R0jQ
`protect END_PROTECTED
