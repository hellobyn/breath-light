`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9r8gBGDod1i8xzWHFC1fKjCjro0finU4ZFQmE4FLKfb2urtV0BRyT+U4aaFGN2j4
qH1JdH3WXDrskJYCgFrlNcL8QNlHK7nu5G/RWd45LXCuVaxuJmlTHEhZPdwEKOJt
ls++vpjSRm5hXkuopgjaZ/90gSgrn8uKqCtuDO3uNTzuVleOL3K5rvtpZFwxCiJr
0Iqtv446uiUP26UGQtGXWlrKRzQBrjiMWEIFLaaVWrYRgTTNCWNUEqAPA1RkM3Q8
gfjRZSJPzNPgWNlp1ye6VNv4Sdtf4toiwDfPF7IzarEhbHyE3mLit6JpvoW2sau1
HQhaoN4ykPSfsiyIl0gZp1maXWOUrx9tISf+V3h9Y+m25/GvSMjdLCywrOWZCXAD
IMeO0iGoZCa7QchIWxuaac48hyy4Ch+OBU/AmZUdV7nDntIxw05bquiYxFgLUHL9
5L1vINe21RDkNG8jjHf2pP/vPYhlnyZRKevEKS/vKa72hKvIUaArnk0dUUlAStng
6mY+13mMHXSHJFqL1EEVRoIxKOLXwIPDqbwSmxvO4mAiRs91R72zaIVlywjMlYeo
CSNOlnFds1wkYRB4zm3Fo5uL0vAv1MEB0b7PsU8AE/bhkdY0NMjDHaiy3h/8cGgm
XoAF31UidOE4OQKHz1p7ngc5pPm2wPh1hWVN3bLf5d3pAficInwdfMk2kYF/TYch
dOSOiJc8QgMPap6JLTU54wbovZhPvatyuE497aj/jQ/bdWjwm46TfpfBCcs6iRfN
gz7FmIvYMyIsmy1ihL6f00lvf9qgHyeL0bmY1sqLRMclDJZXtWh8Fn7e0ZPubqAQ
VDWz2eqPL1VbxGqwpcq03tOtvfddepl+7qnjQ1xBGyBi+8UhAqu6HFjabs8pgS9N
ltCk+faUX6D/JnrP3mOz0AR7yFXOayTUXPMExCyGeUO512taiTMKKVLhfBwvZa0i
HuJzHUT2QFGEcAA9dAD3Hbpv8pNw3pSANRc8SfiRTTQ1Nt58vnP9Nc/B2WivQDqP
jtsIHMgKWB9tImz+2NLIAhki9WyW6aXmNFxz5vwKzmErUoncyLdBRMduiXWY3H2n
K5bxjVjxIQS8TLqFRPzZ7/dSYyJd0jlzFsimBrHtbmc9qUlx+kKVouHrhXsNxmUL
6XdJztXE/pk3o+3IbeR0RvR3qUazUE+NU3qD5m/BbkVrPk3OK+R4ZbRrRiLGpLCI
EgpJjTOq922OVxZLXWu7OlN2jcOIOoQLZtfLAyFmBrmotC9FEtGcW5fx3RxVWT7a
gF5iStlIFMp5ZGWLKEJFb5e8uD7U85GH3+q2/TJyIacUdS6gR/HsJjiR2117l4t+
KctD5/+PkXVrKefAGkrNLjQJFgg+vUuEB/UO3NneE84OW1VGwC/oYhM6mVfjSdyy
XUGleGhY88KcA9lYwI3vpX1NCY7SSCZy66pDf47AVRKZropjaoZrv9YwuxdSYjME
qTW5IFlETOYDZk2DSBtHuo0B7goJwJYhxzzljnL2dcG3Go2sSJ+giyNEJ4COt+mi
cUKLdT3eRei0NQzAkWQqirWTNStaMrNs0uzyRoxBYcMKZP94DWQc6+gB9D8JeDg6
pynDFthSinYXhVP0i6v7A3Axh6qwcOsadT9Co4fAL8uFxqp3gSjTX9GJpKTRZMEN
QyRZWBfH/wdTTx6LTYoQ2tshnV7kCm8cyHajX7v3luHUBIehVgQaZ0zlepPgAKmu
8qEmPAgKevO2KS2oMJSxYALRKTo3oWTPttW8gYUgVIeW2DhJCvlQWK/WwR/YYNPt
/xS7rJSod2ljQ54w/1C1suIBoJvf5PmIwHtI6qRxqlqzUj7jdHfIi20gygKosx7U
0GXoUWo/vfKEdMAuCmz2tsyMn0LGTDLjVdSfCACn6nKkO/Pr6dmxkMN96QbnR6jl
wzuYPwZBexcKger9poZnIg==
`protect END_PROTECTED
