`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRlAXpAg0zaK9DoCH96VHBlB3fZY0QHr231UlFvuBar8jPfnLma73WMgkLDIf/41
tp6o2z/hlmPyNAGsTESqH3JCkq3K8BjYsWs8Q4AKbwn4oertYRqDNoTPwFNnR/j9
y93QhmZTZDPM3UHiIEfNRVujnCyAvN8bytNOJZ/u8KDbteSIaY5HI5PU4yan4pZA
m+L3BJ6v4hy62VbNxLVjD0wV1KXbJ5ofbeGv5LSXR3ZNE8lCMlxiEOeQ9bQJF5fh
Rbt/l9jwXOHCLJp3lFLPZjI4zoqt46N/l36vVEA7IRVTYSEQ/qFFibgMww2sSpnP
bpj8I93TzIwAj6dBKPRyfg0cNa4rvrSFe8rGMjRHlifJw8k7nxxZzN3Dx3mdSXSY
cClmVFPMDBh6KKdRMrp8XqswT9BIlQUOQ8TGfBApbuSJlg/sX94Vp5X+91qmoYbq
XN2dhOEeBXx3qgxG38mCEX2Xz6RkV6nAaipSvcpj0fqU8Chs4GwstuvKiAduYVLl
70vXiCGulsJaxg+yiJLmwA==
`protect END_PROTECTED
