`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOQbOT3vaP+k8V2eI0EJ7Qbn0duzxTJkemiRGpJ5O4BGk65rlA/RtAMQllO4rSwe
yVEnlP+QYdX7+1AQUWvav/dqkwbkFeC+NJHuqYy3FhOiRv2AQaf8CQIWtGxenpjj
hyRSHZ5N+2Ow0/Pn3jQGcEs6RiPmyGEFjv3JuIFPmONMB26c04nrWKaHqedN3rRF
rXoAwAy1mYhr/ktiw+/wyolKBHMbdQJrPmcXmgHVWB4WKA7SxfhRdHBaMNwHOZHD
GpWZd9agVObgpU5kMlAc+SBtVqupCgWWZiLr0gZiSMvzltXrhOBVI2nru7D4XR9r
rOYBpgCwXLChXQ0coknTJduelC57rzGIAalgot/tI1WA/EUF0jZ3CSCWvXdRf/NS
o4K8etkBXmq3HwP7coT0Z2NHR2b+z7FFoMK9HgHHOP1ia7ClcQ9z3/ZCTKiMCn4E
L5oGO0hTdyAzbBivMgGn4zuIGGGbGY6w49ZQ1w3gpcsT0q22K/658ypCE6xbuHg/
Rrawztquk+8EgNa5ASwoMWnEgLaMwJuaHmLd1t8qEi1HY7gqsSKEqq6csCvRAuF5
`protect END_PROTECTED
