`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rK3tYftoZddshrHFOpgBg4dBvtcaDqXLnpNnm9BVeuS2u1l4QkurB529L4TFSHHh
Ch4Icct7tAyGSyQl015nBgXQleVOfI1gHwSFM33fYASdEaaRlFcYQrMFiUnrpbZx
EI7yfU7DFiP3tkBaNMaLNKfoVgrNNt4WDMXvLuyS6Okk1RgUz6xafofS2T6J4E3H
OYtjl/z/gH0BAPcMtcMpA2cJ3NkChKB6eh0lDiZQF3KPFo/dowdCwP84RKhIUnKy
bTxGhTf3uUEbE7rYX1/5zv0eqOt5xhCP8LtWmoyebIrkmwIDGXXoFqbd9wlPz1S7
6dybMPLySUX/9fQqId5C5AYJs4Y7kh3vJ3QvYu7XovlbYPI20+AJ/7BmkCsgu2Jw
oPWzSFpdFjGTWwUaD43SxCbVdsL4RErCGb/1eJE4CkhzP55w7qG58kgANlhFAzet
e6TQyytSuH0odBlypAAlV5f4ZPB9ah6w7EZz9kAVEVgM5hYUt1vVdX4vl5As2sPe
gyq8iz0qScB2VKmf3xktMw8okpTWpYccvH35t608zXorVmGsw4p2l0eNXX4DcR0g
kNevQJOFqNj/fsK+dgXDVEtzw9Y7NqyOrShEyvkRtBqVafmLtpuQEsROgUoiNDxf
`protect END_PROTECTED
