`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8yUs7yA3lV4JqjXoonW9QqUdsZGMIqjzlmdbTucovtWugvPkLIVkBdyFz28B4E5
T4+jlC5X8DCwyHMfSZZf38PHiNNOE4mw1+YZtLvZHQVes0QQ0WAPi3h4QS8rie7Q
aquL8cKtmdL+Dih5RAPfgvzz/5xdLxMY74m9vnPORk/x3kuJydFbd0gW6XCJ2WL8
zamDv31Cd51h1I+fcskG5cqCGv4XGGGSN5XahlBAm8AYKlDUz71jejcG5UjvlSlf
wrOuVcf+N4QuSE7GoLaynw9roc8vtoI8Qy0YRzWHWqCqeIIXtsotzU8sCMXxkn6B
x/iUd7OLchmQNU9gmzKbbn4kKieF0SrGDIbxhapkqtNg/zx84lAg+CrbycCR4YTq
9hsUgD/tMmHA5kkfH28U9HX5CZP/abwpGt9oWL1k3bDXrxFMKTd3SkOL0Q8JhUcW
x1LDkJwijwSuh/SA4d3UXkz/HywKnSlQKBu3HQBCNLwF4Up3NHcaSiw2vTs1RmxB
qDwJ2pFaiIPsV+ZabkSywcEJaq/r8qDKZHkQtEdsLhmI4AvKDKMwNTIiSpiALHQr
YFt41lbwh15vP5NDIocNsuZXLvKNX25M9VqA4ubLNa4cNxpL+W/dS26oucIndD6c
8+/Anrk5dJ3yxbVhNlVfN3dN9azNdynO1icNrffliCuF6LnIWbQTLU0cOGtbHjlp
g6TjyQ+yDksQk7mi05gXA3BfovNGSO+7N7ZR3fYRf/PZNElrJdF3NccM2LdAH57+
ZPgOkrLX4aR2St11WTfGzhf4xi32fHQ29cjwij38Om21x3lOpV16iNrRZLWNIyeU
7U+mpM/IheyofedoSIuabNsoaKacyUhCh4kBO0nBHNmW1ZZHKiJ9I5Ih5i1oHc1o
0/GeJoyiiHutoen9Xs4tu69dLosaou+JvPWoCBu5yxHUzZa861ai8Yi8Uo+phhjK
mTPpybltV97AUbv5oj6kThjsjUfV8yoiquv9LSYFCqY1I602Ub68k/zqEOyW5loY
COkqyXIYXbh643nkiYbXoqcOj3MxTuLjxXZg26U4Q4ud/UD+MpApaDDoNxnzNj5Z
`protect END_PROTECTED
