`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfYVc9XxeGvMcRWBj8nAy175/6rHcu2Q5QoI6k4Rz3IlqR5mMMNJvFPltAXUVGmW
ilxim0gzYHoCAtWmi5abGyfrCTqWyWGyUT1jXgcEifvT1C8LFXKIuqbFJO3tO9jE
mZx7YOmUdH7M6Clv4/rehYQ8Ay0MnJ7/l4xexh64BH7UkJ61ZKGHmhN0hbHQcWZd
BiQAxar1XV9r/29WdJxGZs21Ctz16sNRcNd/jMDSILNTYoCh6cn+j82TRCM31i6A
VDejsWS5er8NIrDoj3AbfKG8VWKqfgOj0rNKgMHKX7AXyKwrHgLkjCnrorlB8yE3
tipFxKlif4ZkilJQQfiI7eAUTiuAvY4ioxipq8WkVhpvD4mI3xKcADIKY5MuR7P5
KSx4LDg534tX42g//ht++OtCeCBQAoG7buTY1BdjsEgAiTmxc4iIbSvD8niFWu70
9cy+Uyk3nnoZetbvg9vPK/d1iiAAjtsqZ/g/IvzvIkFCltXg16onhyXXomNRZ8QT
2PMkooNUzYo2/fJoJSUyNA==
`protect END_PROTECTED
