`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYTWiTjvS4fpFAElsUwARWRkuFGs84kesgm1xjLlpjrSCCEspKQVuRI7zcSZsrUy
F9C2o8cb9wBk2m+Dy9PHnAGsJp5MxpyVxlyeJFb7zcKgX26MJ90G++QmIzHi61gQ
yuRS+hIfyDUcmHudosq3wvNg5x1pWTVCUxDCLoXC1Zd1tUavFVpWLHBRmrNiisz9
RsxbIWackOh3AqatiGY8dc22Rr1IZkWTZFNd+4YEonylyrE36TSnCkrAKmIf6S0f
yxXRJuUbPL5RiOnIY+ELpiFBeUwgyN9kM9ggWMahdwBNFACv6C5GW7qesAUD6WC0
egqxUDaJiX0Z38ONpeDZScYL13eSn5BU7TO+dQyHMIa+GcSSjoIeS3qx8EF6ZNK8
yQN1isl7NILkfrc9igPmTqEe5A13DaN+PGP9jJWXLeIAOWLYkXDsuw7qbfce0Web
q+Pw3GHozRCnLC+S0GC8GUuW3V1cGTolFnz+a/EmQRE0ocP9NWuCsIGJzsM629k2
JQq0r25JHqB65gqnrWLyZn/kJmIgfyNWg6vVElt8izFsHVEN/LCO2CcewcQVdQrB
zWXuMaAwl2QZ6/8y5xNCtWzjn1D7/RBDGiB8Vw6NNsNaVTp/+2MHaHpKBgC3rjX2
rwcOYnJgJ52+I5vpxC16zDuD9JEUzcHqNGzu0z4W4b1M2io9VhNqzmnHabxVYc2a
fbF6ok7rgmB0wi9hGxzLQJLcTQJbNLWAuRKjx/MM1QE5YALDZmpqvQV4PpeR3Vc2
I2b2PSGd1wWashJ5KCD+CxpJ9jYY+T1f7oWDkxWeCb1KhVfnLgMiEz+oAgGT2/RK
7zY3dR6mWCwcxqsMgFbrhiA9oQHWQY0VYITQnF32bSaF7Hu+QFUeSDe0InBXnnyd
4+HBdh8yNqnAXSiKBEVSXqDdOpfWfaIMxjAVt4Lz5LO8yLmCJq58Zb/GWtiQ5d0L
TorYk41wC0MBWgTLvc4p0Y6OAsjQm/OzADWp1bvWm3GhAWBbKMpByTnSMKTZ7D4I
if10NRU7xFa+HH/M22f4KVwoF7qU0DNMI5kYecJDL8S8ijprBy3QmlvCsnnxG87l
UArAL7Qd7z13JayqWoJQEK503fkiZJuD6LUWRNn19uK/rokc9DonEsAgfFB7fXGI
e3QNo2tPjgp2FGoO9+T77jk75Gb6Q0k4ofHc0/5HGDtsgc3ag5ctouah2aCWgMjO
k9IE4F+ZtezwfEwsIAO2Xy5546YD1Gy51UsfH6fBoYP/+GfuoBuLBA6eoG1CRvUo
v5HV5AS7kQxCxbdSloKzxMgGd+Jm6n1HzC42tmA5CeHG8fKNyQafVB4i/+07bk2W
Rp4t3MehlOZNCV15ZnXWh3GyA2D8cXk0uG7p2AG3m0nesFHhvefPJXa5oGgGIJJ2
HEWvnJyaOFzuJ5KoBavSaNdIWCccHs9WNJaJ5JdGVQX6ZqlZD5agFMfvOpHbIRBF
`protect END_PROTECTED
