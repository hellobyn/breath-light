`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10GsKAJcaPNunXe2VmORmQYjFZ0REELZUoGSp0/JWnEsnTWbTizOO6PlikScPpil
X0sJjOl6kcKp28fYzkD7qqeqd8Wk4hRKdxR9MP0QskKYHbvNv4/kGAW3qCuYxZPI
x9Yw1J+XrdKNhNAUSqRJF/XjABzdqeTMypu7YNMTYl5UOe+0a/K/gduL+kGnEQfT
vaIIewyCNOUgCCIk+ns0MAGmSoWCZaPHQjf4bvA+VFanS3aGueiLdJXFDJN1yyXN
d/LmWVbtWueHlphQuaBGvjD7GWHT74hd1/liRnpfMtoJq20umzAULYnzg2r6ikmv
c6+LnqVCah5KmOKxx4e+9qTMVnhytHwnb4ljumAksU4ttqQuOpqnYa6QRblYZXtD
rivXGyo29DVSRPBU56+/UvDAccHY7lAV4CKn7ssyQiyHF6iiL7bZ12m9UXMoOPX3
A5BYlTZAnJFWW3xZxGQoZjTPKr0MUefa23iiR9miCzBhx1JGYRGuyU/gN3/XZiKa
TASYU+4rjcRb4HwZLAYNjNu7h0vfajEPPvGhK5eW80TPRy1LILYRHrVeL+/ebyf2
mAIUbdMbLteJrLG+eLdpdr0ytnDn3uw4CV9VxryVYZirgqpvPX+D2uJAYDOKtb55
jfJq6AiyVeAEOSsFACBMuCin7aQtZd+lIDm9g4wbnwFz7jn+pjRxfmKWcLVAPG2S
xxo50GlLDxWwlROvXZJqudC59ArgrstXJ8GCwljCLqj1z+lRi3HdozvSr/efGS6c
R/KwUPn/3qIps/fb+qkKBaZomtyJzSamUzvhpCDtmaQPQJgz5V7i8nYilEiqAWqT
EeOLAujyqoLgc63fUwanjKQAEK1kWShcBPlACFs4MpHt6f0MoqC09sn4QcVKP0rQ
xXyOjFtCWRA5roHA/yfPLF3/RO0n7miaQHBr4aeDURrNYsY/mJyDNk4QtW0EJaLB
4plD9MpO11f+AKfr+G94TJKbQyYkNrvcHdPqaDbmsScUYVq3ZDJZp3Wl/h0HO+EL
mKZMyUJJTss7eV91mu9Cj5vXl0bTaqgI98mUTutPEbwSCvWuinwLEj5xaCXgQMB9
xyh7VWlXI0EZslVpqLibohYgY0UFybf0rwbbIU0U8/b9pAep2UOxaDOAOXVzJbI7
dN5IZrnywyIH5sNbdhjQ9ugVTt0PDIfT1OqpeblxHHEUkwnaX27woV2AaNxbiKsM
p2aJhmp7/f6JIo/ApQj7FKZFeS0HXe6aNtM/w9+EamyElgssbg77OQSeMqONupn0
Eul16Gq1q5yrfNwC89DIGR3XGWmkSjcnB2ndz8WUYdb3Y7Eer/8LlFnRPALEAAcN
ecnd2034rPqpbMpusHFDx2UD4BqU81LuBRm5I7GHEtqi8BcJj3zxC9SVTRM3owIE
VouVNvCs9M03EO8n57Og9hgRLbar9vVdXLfQNuNvyVDnqLGOqTqzR+doUd0Gexjq
egXKspQoWS3zKknLVPi8B80jdYZhdSJvizceW6HmSYQKUJFvxo5mRJ9NIWT0q/Zz
LJfysq41RnkvjNbz33tBf3Lhdlx89O5tUdimbnYnOUyvJPpc4By0W3G2ZXV+eP5g
vZUvy2tMMvP6a5e9pQwwrHOpt8xjuZjCtFFza1MG2E7vf75Fe5p3Q6uZSe+lsn/Z
phdFRfUnSAp7oUkb20JQjX2zhx0ug9RAgqQaE3N+PPMGFpkqKNNSPkt6tQaR7drA
J+i3zdwB3SjYlAma2GrswTnrwMPnX9WjSvRdc+DB1zc7E5DVC2e4CRqKwHb3W9Sw
Ky7E6tYs7wwA1zbSwv6UgjV2X0NilHqN4cNRdErG1oMDb4KONoMAUSo0UHXcgqLB
bsWECoJL1sJu59NFZFcS+BSrHb9+m0ys1zGTTjoQzg9ajTGegkD0nT2J3MrCLO+Z
h2HSt9wAzvqW2yZUPN2NbOf1tqp6GoqibHUplLRSgci4m/09FWRGw+GoBc+p83rn
KCiFZFvfW+EXQUkq8DX4zKVgoSC11Zoko1AtWc/vyRgVQjwESoOeJFE1QzBnORpZ
1ekWw+sS35GUxXaFbsuqi0OKWBst9qDc1UyvYif+p3bGypvabqA0L88FXobFV3bZ
NAmEkYM7vw3gj5KLJVgXR7iiJZjrAEkT0wvs8RMELSfSLbe2U8KbWUC7aT8shSRv
Yg1izo0P1AoCv3xBRvIQTDbmCAnxroWaZFFRsIIMYl/qiDa6ot8vhQIzk/97jazc
po00/yXxv2wsHGONOEa5vMDAPAjIo26++r/d5x4qvruiEqY5bg3XD+u8uAWr1In3
RpKEEMagEAsG3uIfKl276fF09vH1HYQAZzYEf3MYCirDHrsSRpbXkeG2XjAXr+Qz
ThnL6o86LMpRINLhjBqkBFxGRsj/DFE51jF0q8ROFGYO7p5yXHkCwJUw+7YT4NXs
obv+Hl1ai9aSSIgUf8BCbuAcw8HTmpJfse8eTSRToQT31G3ixhsr/C/sN+xQnh74
I2Kpd3BKw7vRu4ZYNqHzfyNOZUGorpAodJSbw7kaoZ/3YezWvye/sKmP/BEbOMkl
FDsVbyO6eANcybK2F7ONtw917VzvPK1DdUEA5/jkoEMfmVu/mnq/irmVKQJ6qgqX
StFN0AZUuq9tBI16M8BRLBe6JhVRd9MsYkFAbX3ACpabVHqszQVS29Yop3pb1fZu
PpGSyjdhjhld6FZmI+jB2c9OHAvIuD3fLEqAET0e1AU88kcWJZ5+6H1WYvYVtDci
l9AXirIGAnRhUMph+oaLXQinIOcxoYMtnDLCFtijOoqcamjkW4hLxw0iQbVyhiSS
5jEhmcxriGjnYsiZpwkDpsBCVLdI//tQdGP4+dzE7Kb+IGs5HT46d7zFE0UpffLN
VUVzdkcpqxRLXfk/FGjbCwlTuIahFRNF0GRH0PFcHUXTXsm4b6b5kaoCM5jkwSiR
CpFOeh/MKbrtvt5TtZZ5wC24Of5y2lYNH4V8aa/fwB+keEDrewT9c1879/E4hpyZ
JlBjsbFbaM2ryTzzSv7bQrn9GexABzjlifBUaNSEuZJ5NRLjMIpEmpJ5UdQZFcC0
GDvq8zINVaeKERFbhAn0xu/poIrYdbPQtkZ1NdTPWC3EFmhd/glDXt4l6EsL+HqZ
gpHxa20eUhgYj6v7G72S6oidonEy8ItIeQkJs0I1sEavUMqIVyHKN6wE+t4E+FT3
34Y4Xujk5u0emNBi5PbJw72WqJjyNI/EXDBNoTtjeLFqV9mmjXWS6ERF8xTnnUQA
nhIfw7Dl1Y4ZSvOk9W10yQ2L/X7dWlP+UsLFEVIjiLarpOQVDidWkjvCJkNl5nFp
AR7OOWw3mcr8ZZUcyscrZZ2hb5nfwvfLZftcMRhttNPj1lRdLMgqM25C7/iEVPm/
T1tEOoti2OQEpBAYHAFSDBYej1q0gx/xULs8SEpV0pc5+ft1OI8Ty0o68ujMHBs2
AEH7JwGh1RzDrLcyEgLw4GgucoQue8RR47lg2n07GmBUn/QdylIoOMmDnqU0k++W
X/yjhgXoxxsAe41zCVDX0GTAUFvKNWUvSiXFbkTjFC5QyE0UV8Z3Qszgf+RFPTsX
7jZzmfuQbM58uUibhnmPBOTBZ2kJ5NEprjDNCQWZzSxdOg++3vMyV+1LW1W26LFu
b/AAgMwj3O7sPjYZye8j78euc3yRwc/yb4LuhqAe0y41xMGLzcXexFq6BI4IRlPC
QihXrlXtDFhW0BrgbWaHBw==
`protect END_PROTECTED
