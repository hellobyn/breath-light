`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xm5VLBwgF7pD2ueDq7O+A2iFgPrdDX0SQGaXa1MscImq0O94nxIWJFOdQG5Ox4/m
BFX4vn3/sK/YuyXDSRri0HHTyA2hnZosHoGcdJz8dERgI5MqRl9dRyPxsLnEn2Hi
zGcBR+UnSb+egZR7WgAAVsEdEIGUOKealpghvlCGrjKdLuadU0pkCBNwLDxlOIDH
Jh+2ri2zmLbgnVr6xJcmpoyfRkPpKYzFzF1WiZZq3GEHQy2vQBh6QTYQ0s5LwGju
vQEaR5n9kLONIGU/Sc08X0JjiUTfLtKQAFeWHwnX0Z/ZIdZgoADne9cwR1tYfyF5
Kqwy+K5qEHH1qjbPlhH3lnJvHeoDUimxGX+H8w92pmhkuyfjBEZcPY3cIjhmTIcI
v5sMh0vuXH/IBwc+EdAveAEHqy7pH1et3NQNwm6kPQao3cLC4FQoXF2HmxFonsnF
FwYyIj3pCpF6hTpz/lS71lSH52SG6AlQIWGVXB4LmGGrv0+x61wT6BpLwnIOvD3I
e5RukH/3i78W+9a+LKbh+EY9a6rLvA3T8aB9sUFTYO70EcOTich/JoXMWSeek+vv
SaoPdwyu775QCS2rTj1R3IchTKwqydIaWWqqiqOcwUIu1cVoZih93xnDR+LqVXzL
gbaYe4+vEKYP0DnV+7f/g7Rh92CbIdg9moBHLHSsd1Etn2aR8+HLYPyuuzK2YXmU
T237mm1mB5/vQ7CtF0aMuxoKzTOSGGPsh7RjMfZr/IvBjASWbyVSRQgU/S18GdwG
80DiwrmkNo6iCsM5R9XK3FqfvNnQqcSP4XNelaxmMES357RlGyjWlKPVP54/3NP1
PKBIEuMwGATrW2seUjc3VizQc7Qnfq6bmrp3Gj2V2gjEIPGnEffPWem4VpDB5z/n
z27gQrbphte/vl4/zHZVNhP0nPK4ww21p3o8HWBoR8g88DcpB7mqomWUBmLqNYUl
w00cPJklQAvaq2p1zUJV1yBdD+puV2/GPPLzsRp6nZHM9wjYYdC7oe0Z5v9wDsn+
C7wUc//brON7HhjeDuXwGDRfoLB7J8qrgQmvJG/AzkHACbkGLd4jRlRxRplIjkO1
pPE6gM5ag3TjqpTCOrtzwmlxt2Tb5zx6EG8FYwlNm667l+MUCPeXlnPMsNF1nkby
AbF2DN6gThAU26zWtPsbiN3cipcx3ZZppYcYUW3q0u8X93EkumKtzK/vhB92l4hk
exKQtNj0Hu7NP1oq9OGaBCvvty0aJW21Eq0Jog8qshe5kdhIKjkHdrlLZqGWKPS3
wSHlsA6YejLZrIP42j952PEQ5/CMZ/WXjAddVrIHqkvPz7gaAWfCbFZrtgCQK/A4
xfUarudQhbH/uH8O920gGNm0bIJcwitZbzB3I6zdz7NV+gfgYgM5hHAqnnihW6xc
icqoJcppkzLnrUFcyMVECXuik98L8SBT8diTG3DQRnt0851CgFP+R/jKI85Fl2vr
GkbqnWUW1xDaKmmcmKH/bPAswBdehuL0n1IKqcn/gq91Yr+zYN8OiUtbJ9XPS9+U
u32Pauu1oqjST13KGaip3sTyRDrh/gikQ7N5Dza+QSHEByTT6Qme0Z8OKKGdBitR
K9Mic8gtoHelxc4WNbgHCdrVQQb4DEuAFSHGZ79AHyuZxbWIHjH6r6lkR8F5rTC2
H9WQY5o/x2T1+WebfuskOkBYWl/npoJ6TTYJ2b1H4jCpArVShGScKRxPY77d54zE
xasOMTmZJYTfcR0cQeXceiV0l2HdGT7EgT0KJ+bNEBrZSrZMssHUy2U/IccSYppk
zmoR39/KRK3OFlUmqbCfHP9s1wIbLY2fdNtqtC0Z0+CzcT5xPfdhTlF1Jkw0Ri8O
awlPf8ynAug3S7xUe5GfGiBSBESDbd/YwRfdsRmdntIMwWG/F8mZ5msjuW0IbTax
0hoFn389oK6DOCgwE6ozIsK96N6hTdjkTuff+QrhKfotVZiHc/Hgaf6niqywuD0N
QDLu+wAunwR1pHJ9+IdTTFIr9+GMTqb007iPc0AWzykwKB1E/42VSAJrx4ogY9xg
wjtCIHkODwhwWtrba2zG8o68XAWiPHGCAelXzPw9VDJPLXaS2E8p2aCWv5vR0RI3
mbVR77sJT4FmfQvtlUZrN7W0mLRvTRwORFIXKaYpKg9Bviv6ObQo0VIHypktWcA3
S8wJ8d0R/vfaA56mMFq/qnF55UKARhYz6kRozlcMiAe60am+B8KVpl8gdBew58S9
caG0EuOemIgmCAFqne/N23vxAp80UVNJkTsMx0Ee+umoZx8PgCUJrG4vzjWIiXIf
OUTkNKUB0GntdjgwrqZ0BHQIX1ZLHcAq86fh0zKlV28N0VDqssZynYZ1NqrseZaT
a750vhuOrvd/VDBesShyQWz/ckW18r/j8Il7bcuwiWD4k2N/25aWEr+F5XnTHAx0
iV1Sb0Vf7SdsU13VvkOIaGJQ+ZhbNwvVsFQLCsCmm2D3LyDOkxCJhMNnBKACBjNK
NdOpgo3xA8TDajYn8lMK55U5eLQo19+EyKKF+Ws4k0pnCvzjiUhlUSEh/CibD73o
DiLNaqWkAmP6euGFAJg/OBzQnC/+lNGmCEpwgTZfJCE4GEA/c9fovR6xS/oN9Yv7
ZX3pVxrs/tlNiUKEBPCjgNdOMB1f8ICwQibeEOj9fgMOKJO0cxP5XBOZ/IQu//O9
bNJGPW3eb6mX6s/5ekEtc1uKtJzAuTiCDudk47/XeiXraJncgSBLHC4g9DXs3jAp
iRNY1EjSRgnR0VrslvKHmNK7FTkEXcleeI/RKMOdEcN9kdbPQ9W6DecB6Lj85SFP
dz9k3vX29fO8Y5AT/WbMRJ7W7GMm1h5Ex365vauwwd6C6GtOZlG8dGFcDcSncMSP
b+pCqQFpzzWV0ygrDs+4m2HoKSoTpHyxZiIMCbhvUGKhj9H7pLokJvLubPu0csIF
u1JXo6nu/QYgdrCm+ch/j4MhJcjuQIhhIsekl1WC+BdM7LqJ9f0borbueU4xRWwf
6J3JLSLscc/Pv7OA1qh/eZgiwTskGq9dXgXexpjmuAyYks/I1MzNsmGnZ8B6eH2h
nPXOBoDKAkBXRt4kZNhOdDcA2tzMuZ02IAkYflqBgQHKEsH7PE74j1ApKILSQ62B
UxOVA0RpbqfSRyEExwjHbHth7edJH/QjIQPuQQQ9psvcLogBykGwMz6rALJubxC9
NSGebRGlFYa0uN/fQEg+yhpsZRZjKK3F8tMuYHsupRV/VdXPYLly+tQ+01kp6V94
W2sg2Z/tZ4SDR3DdsDN2jZfW6AmBkUd11dFb6cYZSvWM8Rb1DPLzGEl33Sp35+qx
`protect END_PROTECTED
