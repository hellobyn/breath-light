`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WvbUkbBP8lwUJzMP+SNl1pnvw4YV2xUmBSBKUdXrN222wl90HB0adethq+YC0OO
+mPn6B+SACAp2IlVtO9cnCe1rrZF5o5kQGmfio8DTMY2baMQuZIfcHSQ81VNsHlq
jw+4ov1DmokO+dD+x3TL4ijLW+zVjJ96HU8ltwwp4VlXEXMl1utlBwnje9jWBHMi
4AkZ753PYzsXJf/aJ3zld89frdf6wGZVvoxxIUciVKGzQ6wT/q68tlkynNldqpjx
leTUWHQ4d2NnEM65/jhcqrkb7xFgJ5KYczY6TG0d+WTbUPkdPBRCgw5nod/7kfGp
PGDL5NXwXZ06LoleRBQ96kTQYP2YcvEFYQPoA8xDnobtHXSK8DrwDRKRNR0p/ZKz
SsI2Zxn6Nv2UvZqWO4E3V4rgia0ncsRuVEjVZYl5+mwir0jvCSv0Khyft1XUkHMk
YHWEx0u5iLb48wCb1TbtOgbR1OxH3VF66h5jSzbkB/cAHhhvr/MDrP1KuLR+z5Mk
3TONzrH2OY3Hl+jp1WL0YFG4nP+ljfrJ1WzyiLzSwymEXLlz+grNwutWmqMAUp9s
0EQ+3ZPPD4C9Nae8hn07eL29urfzi7dDjq30pI2/U9k5Nz213sQVDyuYXg1j7W7+
D5ky4sgGOKexLFypfFSMftwGTQZ59aOJizO8SWOjkt6EDUvir4fXsZ8ezU07RoQC
aFsseMF5vfc29/faHKaUCqq6Z3kBYvjqZFZ/3VxO4s/D/+YMGiCFHcxPJFUzVuMY
4Jq4WzV1S27ZUFgpFtAhy0aw1D0uMErT5g85TBo6o6Hmazq2ozqooim2+1KFdtaa
W/5g9bxMX9IF6tRO0dnza47IjEnXDIbjVdiqai5R/Sv0KR5QKcolLEgiWcfYuhY4
rvpn+9T4jNMKKCJLhjNNKJiM4d3kXlZyM/9YBTi2BO7ByhSZLGkJOACuwiqk4bmY
1Ijvu93bh9ee4XfpKgKOleEYmugksrze1RxntHwSi9Su7uBoCtLNgiPosJtJKVnY
DlyAOKOFrOq6/FZ2Dmn4MPH5V/g/VXVgtRlUvenXJKcT2pyJL0kWRPiEg5WJYfSR
+s+xvUmH61/a0IsvVyIMwp7C27ap7tTr2cgR4jGm4AQ8cYtLMfb2NYE/EsbmtOP9
E6L1oQuj0/pXdH5XnE6QwYguKRlmtJ+46d0p7tm7nz4EItm227eT0iR3RoJtRuRy
PablgZ7KHy0YHBST+xe1Ei07PDyy45Dn6YCnEDMI6QLX284mHWpHj7OzgZ/FFZZ7
czOB0t158jgMcfj4/YXVq0HhHwdxeqXEngYEQqnyye3wK/jZWvXVXGigt195F67M
EUJYClQSsiBSp8/jUo8OSDG2cXGHPinUraMmzE68TNmVvpR+NOcSPIRBGXHae5B0
4XtjVhjmoIVumeuho+ejwpb2UvFl3Hol1DiE6uhHdEbOPoPDmRLjedDhuhH0giiK
1mGvoLw7io69ugostsbP5YWQ1NHKlAPdThaVNyJSxenY/d8StbA7atZkuiYYHHG/
OfFNFfvgTI+ijHt+4ICgUMr7UpxU8KOU6cy1v3gxBAWZKjR+LH2t6Ny0t0kGVp9o
38jd+8uYeD7HP+y6tuXPyoT80NWO+CAhd5egTIl2d5yANLt2b8487EPZZdr4cYhL
C9Kkj5iuJoI+MMEB5nvypWxWXbSsTUavhDx6gsMba8n8mMKw8vR/dN99j/Qe2rBl
SjVHvGccQBJr7Wt/awODD0a3Zjr+dLC03ndfboybf6meWFoIdkVUy99h8v9mX6G3
jGBg3X1xUuSOP7G7HLCnvzFhOcOWdchcieVNOImQRx9dQ+8m7TXzrf3YtfDy+Jt7
GJsX/YhPVh03Oqj34xmWH9lCaig45SErYZ9alsI0vMudpuYQ9E0sy5HqDb70bRmM
GSXBJy4WZe60ayQ6FsyDrUuYxd1191p5CnbGgApoqnUM/a8NC0RwYSNjRmRlUjy7
KLvqj6WI7/LE3czZc6jk4N8cB1t52S0bCyMa4HuLDiARFiAOMPxhIvtVXUnarKaN
/GjpxHGDyF+/wGlqN45jfUlOeXPi8jA2wgMSt47dyoKBj1zZt43kOeaHzJLLZxyA
hIqFAzCfWP07sxdZz8kPlIEIAznd6J+EpYxFlbUxP0xRagMOKJnx8roasCigtD2P
4M0U3bFR4yRrCMCnZWZjilr+V46Qryy9PN1zed7ew7LOIKIO06iJQrlDOK0D4Cei
JkU7lQzZ6hGf81FY5GUrU0e36Umq+SCd5sbnIsDCzF9IdNCpBnlSgF96FyhYdlWY
zvIeq2U+Q7tzq9spE6QZESEYkPYEp6NS2+keKYwjk0zqg88YaLTXfsYJmCV88GD9
gE5s9yADvnAJWcHAZCyyXTRqf+am1n/5Z3lZjVnADQYVTB0sTYtR2KAGIrNML0h3
dnLhfR4arMuJ+VFAU/uXdVf3SrbLT0sYvF5OKM5exavVqBR6EI7PVbuy2zrJOetP
LG/uJY6KKZgrh2e/jDERG88ismoZrhRtz1b1cdVbFwKmkDHaAx214oIMnzd/yKTx
CttYXeH1D7ddB1knbuqOaAu4DfwT2vZO0nGyy1LrRVJ501z6sYUCeQ2sOPZ+XXY6
lO4PMvK8lnogZ7jwPgTxju6CbdvebBQGg90JAj54MNUCpCLT3OmVrFi9bA1zoKN+
6LrcS68NkpL/nGkJd6iIyli7yC7Cth/Zw2MYoeHQC7kmDw1C83qNsbHhOZqNZ2xw
bzFDhbwIiGLU3BKyd/LpCvmKrMpyl3ttrfYfP59qsRxgHImNaM+ud2yjqHx/5wou
DsX2+oFNmhkhg8h5tWn2iQvmcLlGynF2OrulJ2h1z3XB9qWJNuzI4GbrSRu3xqNB
7bTuSQs/nK/fT023NpcqTzgko4zDRnZcU16nh2JbIMoi+GshpUM9FyVQIns6hOov
N7/xRHTGxRyGqB2tPRXqroyZBkTm5SeaIe+O6cd9iiJsIyv9DOQFwOJhSYsNhtKS
9pyCm1NWm2rU+RqkrL6DMz52AWMXIlBb+h39lFt0wD0pRfw1LRsw5Cx0QFJbyT2H
gJIpRvGGeuYkXE9wT85gL4u5MIsTHDuqnbqPNX7mQGM01sSrexQXMun7DGnacOxv
An1MPZIIIsffbjUXbegFQuQ9/v/jWnRpkPGrB78YJI9Msdg9/A2tbv9RMH4TMKyN
lycJjA25VAZX36ducDfOGHkxdIyoZn0F3I7Io74tFm8GrUewIb3qSTCTpfpw2BTW
5uXyiGYAA0FBqZw9xzjUBcNes13A4v98lsLPPvjx1SfiUd9NAXKp/4Cra85UrI7Z
UHyHanuvP/0QoxcZ7mBq8PP4lFuSMCY8QOJypbUXMoiqkCrDvvV3M3bH3jHIwJTe
dOjyW99aM4HV08ZCsdSmzWRni3ER0fgSLcYpFaC+7BvquPOtuxyG8J7mdNn6SD0x
kXRCBzaMYe2lUWTKg77UmTLmLgSrK538Pj6Pmz5RFcynM5QsHy8/DktOak4AIBMY
cXaE/DN57Z2fr7s20hck4+B1sR/qyjawtvOw+6ERG7UoSG05ltaRzjKpJue/3Pa0
IuqXqxez68UqxCwmZZnUPuADZy1cn6Z3AmPAbkF2FBcYajJzLZ4r1aHjBQQCFZLO
/I7WODAzaTWFdNM0+eflm8EKV+JM9InJXSEnJ5Zpz4eNdbgzEo8ObehKF95icUd8
BmXeW8KpEAgyy/h4hksOwIb/i5KMLESf1V1XTo8Y6d9qjnHjLfDUYw5SsfrpGrKr
UPOJymoiIbPiU6I6gNMPNYAwHXenYqEnyau/1BXu6+dzYEUVjkEYWd2s054pwcn5
+IWm0vj42L2OL+3Q0oCaaS+/vTH4X8SQSWHNpGgg8gf5PgEGci16i8sSI3YqTZ/S
m5cP8x7I8LwjZlt30K4KztUee6UOLJV79GDn1L6NAXKtwCVgxzyAsLSe/mE+6Yf2
OlDHCkyOKh8HeGoCP64Fiw/Lv4u49xdWylY6zgjGQ1SH4OQQNmYgILdARJBw8yhh
qoSz7mBT08PzY08WDPzfmpBWfD2decRidhy60cc/hRSatTmAO8Ozvne57QjyxTAr
oJ2XHkRK6tHI3yimMoEhZ6gltpzMDr1zuEMnFnpkPBsrN/B+n++H7/7jhjVlIyU+
ln74yHQW75o435CwMnLqL8FGwCtqegUaUQynHg6iYFroJSwXSruUDc5XEaDOf07l
DlXIAvUXSY1F7E4sYQ7rFkOBAATchgsUlUNMjgJ6+7T76lropr5DsEgZg+u5MB8j
vaf0OtClP3Y5gw9iQsmDRm/2qG9CKs6udINE/pt8kb/1EJo9gHb6hRVG3HmRBk2/
o0uHofYovKrGvBGjjnN3gsIJEq6sbdcLTgY+zokNdXiout3H34X+H2iC/Z3FZPhF
kQfw84hH84cPbBKWuF+Xg+yWhN+IgVZlasjMfX0GchLbhc/FYNIsalCaFsKpRXt+
NPq8wv8B1kUD8N1iM5ERg5906EXLvO/BaOpjP63pCvPk3VEtMt3Ca6APrebYeG9X
7t1kz/L8hLen0PAVc7vuH1omybro5F1Ce5QcnEo/z6aE1BspXCXi9pkIcwoUUntm
yPN8y0ltMhPpeeyXjKondZyHjZKnFmn/+N9nFq1oj7mNZB9NemfiUMJaVW9Byi1J
d7E3FkmIYaClPsNy54Yn6WWjeDoOBYzEyaO83FobaJDsmSp8P7HczeHzsox/zyaU
n9qsLacGuLaX8nROA3buudfWpVfG5QqoRg8GVibHBunWMhozOpOIy97hJa/XrH3w
lMsA+6SjDtMWQXQ5PE7THozyM15PykZQXnzVPcg/HWoKpkpwI3ihH1AtHyPU55b7
De3VXPnXKZ9nqycjqKJmK67dC3N3Ogby+NhfCnXzriXrtxRHLYN8JydNgHoscKiJ
NvrqAr1jFme98NcFIa+WVgYFQ0MeIXGD+qbcISotbIr7XDTBe286f9SHHW8deikH
eOJFGbGkwcJYachnpdNsvHeqp8F8HVuVySiSvCiZ9ufL+NFaFdm6m6LCJ6d/cKt1
VDfsfq3b/1mE7OxjC+Xg/Zbij8Reu0+DDJ7J2hoeyMLtmnndCqqbQuAa9JWsvwQ2
9mm2aIuYORGugWbsNwSgQTW+hH3mjaRzY98ijtPmYrc8itIspEe48zHEYApJ+X8n
o+pAtp8ftu1+OS8I7nd9wDLUcFKjjh/ZORgJW/5pCFkJSd6OwWzSvadidpf0/ORo
1pWXdcRvumvAcid8vwiTR2WNnHXrAfOXonP68XoappyHAStn69bjD9FcngxKvqK2
rDJsdT5BD96q+98cyylBNPrD7fk4BebpXOlSBeMlarlBUHuNMvP8ceZEhzf+33RZ
S67MQ7ZAreKUk87+h5T60TsAZ7U1KVRmswCGM67fw3El73+fPUURAzz8c9ooNCcf
S7SoK9ymMPNKndckpgcyB+pCvFfzSMMx3eGyOFC5NcZxWCSZn1Fy58E+818tn+YQ
30DbMPM9xwlHso0cSJt0OwId/uUZw3vlWUZlOqd7JVUhX4KGIT8GbWJ2gSQ75OQh
B2HXgOwK2CVEXM7+/qvheROSzdQ7M2WeetTKOFEW3XmdNctgNuy4upupJ5TZBw4V
v6zp4IsFQ25TDXWL1LESmKgnizgVGPe/EV9JFctoN6L4Rb89/VBxPqZbT5OFtPYh
Ru6EI1NnT3hfuRXjj9Ts7u+gu5pOrAZTCQZ9n6Jxs6wJOBRfTkCQ2liVZTsjy+mR
6qCnVTqqcmDaDYZXCY8GfFfo+JxsgkNITYXJdYoa/V8Yyco1s+/ZX1mNHlY0Q2HK
M+Mzu0MLyXvtGTM0rsKvaallPVtEga0yP4XuJDsvsnF1HYDSw9v+yJhpbw35nj3L
71YmoMIBOGGMEz+iKYoia1sNTYGcHwlcMksNRUw8hJIzcteEROcJywT0ecO9vlt/
tlq7L0cVVhNZiij1scgu+cH/nFqAZ5RghQ6yshXOyfmVpxLm5Ggz6ANm9h0ACXLH
Me8G4z5AwM+xHERuw5C6m9bGgcfvDhDCQV0Qp+jbu/FY7akcIkBeZGoou8Tm555K
uos8JVEaUMuBq9nq7GTyHenzFdwQqmGzSUoaKt4TWQDqrMGMm3BF/Xbr3zu2ppcM
KkaV/1XtE8bVQWblH/1gwRuvvOQmzjpTNe1Q3NvueHZTLMFhf8zPM0WWiok6/F1/
9AcnMMAtNne4e4PX0oa/JeuQlVCxuhjqoGM28ZEvmr03Y7RTl/QZLUdE3rCCKonm
rAZlOkmWf5GOruosKaVt3ZT4mBYkw7Ew/0VYKgXHAHsyn75x+VMqZn7H7NN/ZlDe
t8pXNRPB0fQKZLhKKuT5DT/NfBZxbY9uhdjoECIipAMve7rS/kf3OTPVVo57PmPP
0wfVtQzFgoufVbZikjLgUDMXyAi/yzcIZCuE5Wqjj4uoYjizHzcd9rNzmsMgcn1f
D0W1VvubNO9RpoHzk3i4g6+wS8cgUM8rQU+UlCDe2RCm737Wz1YV61lHhNktKdG2
QeFQnh5rRbw9nFM5YqEYbIQBqG65ZL/R1TLJ9sDqNxW9ZdESsiuydVXYUUlFIA3k
lykKqIPaO17aEGqvjW+3Dd3B/l+tXJsUk6aRL0w3JkirM1z6fcJHa6RmkMIrrOk8
ECQMuPOY2DcyAOdv0zBcwBoZKsi9T7DR0euld30WqhHajW2HScGwuV1UhpL746Zz
mqQHWZOQweiDT7py+uI+VZB14flmiMdjYUUJixCwYtj/Aw8C6We6iyPARv0WxIGh
mnk2OogIcLC/e6fQevHq38P8BYIL3d3VPm7g13TTgjuEsl+YqZnBtCBwosxMQQ+i
KAp3lNG87aXxKwqh/Juv+ShldZ7dHw/XyfZjD4/QCHl90UHTvoiHiljTBKu7iN54
KRFwFGjTSO591FE3nxuPVKJ+2uWXYxwkgDZRJ+te81Px0tUeBtUxGqJ1fWf58xWd
hOsp4OTr7efAUMFwPeJNDvkTTP+868sbxWzINqjQVqC5yWGvIzBEwTalgsQhmUYV
64rOYRM94vJyxLYT/p2rxIMnWoEWCXtj/WG8X5p6IRNTAxEhuKE0PsSKxM+0KKVX
8/MyWkaJN5QWf8s6KSNR6vQZDFImPPRHPYHWhZ0syVKyRonB4QM+H7OVycx0aYgq
qP3s0mN3ARqHFIl8/ooQtqqxrWYer7SoXrPF8NAtKY/1I7S1MQYRpmAcKCuXwqL+
SDSN8tf5o1gBlx5D+TCNrEMFJJ5AL0HcHoTf8+9m23jXIFMi+R6mPzwE4PZeU0VL
3005KgWJ5N8sCWA6RsWdwDzc36iCDr7viUCR/pI6OHUCcErKBgjxEzbJG4IRo5V7
hC4CGRhyvxWRbqF16Gros6D+ZN6eB8agCohmzlwOS/baAlP6pq8EFyYAcwCfucuA
D7PancvrYQw1Ewh88JaeAk51C/m1+iVD1dYxOsPFs/RBuPMqflkLh91PcUp8NQ7c
aj/sFd3m34Y3F70K2+wyERo4wPGPQ3hRdnkubYZw0lxFC8OkTvZr22iaMsKEpThO
u/N+0m0z0PW9yuFX/mqxWRMcj3c3wki6PbXnJHf0WuUVMDOHGP9rWqJMtpPgOmzq
jY3gzkvZw4aG9pyNPIPohhJDg05gCuYw1NFHWJ873W5cU6O2cveN1GsYIUohEx9p
VmLK7fx1rSFfK5qb2iiE7JecJ5M7aBi2ZrqkUE2Rb5xNEMGoh3aUIxmCMghVoL0g
Egr3yyQ3OmHmYNBOe/amrTQvKo2ygcExoasHFyvFqyvlKMCgh7WyqYoVHO+S75G2
wAaIDNQpqzPBR+rEFsfQAppO8RQ5MtvWi9lfM0rwgeNvXUtWPElevQ8tE8ygExbN
b2hOhw3q4ylSHqMlxCXQf4vufirBjlUOcuxlTolCiZKp3jyN9skJpY0ojR/gnAwp
SVipJsyLKk+p84ofo0/XWtMMUCLd9/yrXaEAo9+TASXOiPhrPuylWHvtS4mLH84f
KEgJCGCzgYSMqX8pb0X+NdBxE5duh7wayojkyGqoGUoj9TmD3CMk/jjgPUARAfuU
TvUMCSO0V0tWSJ21KKDkvJU6RFdZN/GyazsgnmNeO3lTuNWfFtpUfAedajOLm4mq
uEQFSrR4Pb6fA2w5wZoyFkHUp82qcD9CEeM2wDrN1smF4gaCVPMFJf8nHWcIjyal
31I1GO/EQtj/d+qTcniWxYEVkiApY5MHlECyJmcFc6y2Fm7IR+MsmK2EFERvYfsC
6bHGvsZWvPUGC9I89EVRDZlX17ta6GBPRdpAaLMLm1f824P6Y7uBZRPoKLLJHK1q
SSBd1ZevKcgPuEG/99lynvVGGqvyXSQvkxBzqhFFT/GDAEP5ZHTuHrGDZK92ferM
55qvlsw9gW0UrAxpnNG5OX6D3ojeukiRm5oJc8gZG5IGwoL0F1PMpbGS2VcCnHb+
Sqqx28zaWIzxL8KSBNBPmIxRRLSTqkjTxXzZDACCPwVu//sDgE72Ax2oFjBwZVaJ
a27+aSSbHRO+4hviw3oWIWumZSglpUBhdXpICq3/NeRk0bm7F6vhIo1q9KLwgxPR
aMA9YVn1pb/Zja/TmmcckBRtJI57muRlCK594bL4fSywTpvZW+/LtoAvxbmPrvyV
wvjnRLHbrDTrLFjnVYsnCV8adsVAWsiPHftKgNBMY1U074UHbDY/w+N98aTOrXxj
csfgILxNgI0wrQKid0Tqap8Uh+fn/yxn4QwCDtrq2E3wg5UNCFU9jooAYx7W78ku
aoNS+pPwm3u7rYqeBFGihAHNulCoP8vvmW5CENrCape2a7R8Kn6gOXhXnfmO5hdN
HfD0m5w2s3S+XbX3xIAUDwktgFBKhapBGCRCi8OyFDHdcyJ417oKN4FdIIQAuqzf
foUNmymxwcRU7N4I217gzF9XyuP+4GFCZxWqtp1BsatqdnfgNEtEEODJUei1tMAj
bJ5arkcISPaR8OcpUOAbHu2AvaQEu26lYGP6+J0a1r6YhKXWjMLKZPVny4+gzc3b
ZojJeiqIypqjBzMNJM1koyW8mASoCMr3WgMROgPxlyrJp0a5gR8FSqMTWimfT6bd
ZZFUQrGczMqDDwm+LQt9U2tQKfftRgVejB/iSbezX1abVZlaC37oO5ST8hiZrW2Z
emjORWMpy60N3mWRR5JM1qrZf7wmsF8YhhUtA2P4b46aRjfR0z/OidOgPEysHVe4
0wMw7X7bPJ6yISB94C5QRC8k0Y7hzuUVLN/X4dr+YUXVQnv82nFJMV+jZmNfH4eI
GC3TAIJKF+jPpmLgV3gBQVrN4jIDdIdsn+Ol/9YaKtn61XwFqQAfO+6sLod0YF3O
VR6b83qBMH1b3Mz2+O8qtZP40ZoC7n7eHmeB1xXu7dUMxXuyGcdYBY3X1dXFqb7V
hjVL9P/eKHfDo/U6MIwKiGLbsGAV+36bAejluwnbW+9o7YfZp7BDjaXgFKYOKojR
Cn80T7w8ZKjBhyatuSePF5/aICW0wxUE4elYnZQEnqZfkaPcr0432n9oHUGNkXw7
EMUdsEU7NOdD7+1UA4HhCh9kp4fgA61A9dRbtfZXpzUoO0qxwiKgIvZH5ZD/DihR
eVSrFrFzKnuyso5ZCY+sbMS95+wHYrmqP/yg7W+uxsp/I6LuPzB9po80nrFeEW6m
LY1XOirxSg2/6BQtRP/Ld9h8A7BiIWlUB37mo2qTjbIvoWCYiUYsdSsIjIHlkayt
7vcmayzjxQKLPTx1mmzozd7lCsG6VSG9UmixILEc1/8MXvR5QriyMiMV1+/PJuq2
7bD/bkdStRTAU695fd2jUlt/WOBoXcWqa8sVn2tMKI1t40V7BbMHCSbDK/obc+EU
hPr912g8PvLiKlrV0FKmfaRVK0QCOe00JPIykigBo9qM1E6k+xkZ/w5gRP/2ZsAm
3RgGADqVMcC1OSeF2018XLGTdzKhu+7I6Gq5uzb9Hljk3OOZfT6jkdrj3sr8+wED
edwdu4s9xeAYDpEM9cdTmnDoVkyCjgsSiBmtBPWpUDUxzTU9KaOs+sIUbIXklVKF
wJAvVVL7yEY3EzJffeCdr/kRgBSVRJK5Pfh2KKrTRkzTvRKROV6CtAXnfGtPDFX4
Nbf8MjdoLiVL14D+OdyfHhmaSeVkTRuPTBkS1ldog4cNvROOopYqThiBwt4JdzHb
hn59Y+g2IE2nT008ChSOZxHq7Yt8I69PRitpWa+0hDLRpunxWetqWRrphuB7OX2U
doyMwG+I+bto6kFBpp+roaV+aH/jrWUbQ84YRXbsK6mw5FSUzzYXQA5dKj+T09ka
AX3UWCAV17TGDEeN2JO3AyL42LhWyPWH3NTmAHJfZixxi1n3hV3AZZN+vW5QpehE
ZFu9pVdOraylc8mZWOdsGnI2o8DAMhiDCPADtOnXaWQN1LgTqUsGYBGUAw9jLm0U
Y5evInbbBZR2WyHOyr1wr+MhdIEpEd8pH4KH5NY2xxskYClin9s0899M6dZJ/Q3R
Fo23qYDNEB8231zZgplfMzvoYqHq1X0WjrLrkManRUpiOwKhNR0hnGjQbgqCJkf2
otxmew46qh0PjRldkhKm475bb+vJsGK6UkwHj8ktBVLdR1Rte+nQ3x8NsoOFu8c/
m74URhgJ1h7/zCTh6e3+l12K3QDPm6XIPmVoBtPsncuuQnCcLq7h0wDsu/j9AVCb
cfDjin8deIsIqybQFt9vTKu4sNAnO3M2dF8hgXcGqNeLYiXiPrEG4DMDsdESrnQ8
WF88VP4ljUSyxrhGp1mS9nmAA7lXY+cwUuX33E7rmZM4wspXgYGFVG4hzFk04KRd
qoDxWU8fSknlDe4ZsEpjr3BALIIfJ6MMELOXEQfrWbVMfORxRAMuRVKDtokgMMN5
qYuU/TRTcXMYlSkDUpcBugNQGmyHVKRD4nEkf3QC6sVAfE7A6UAApd3QGUvi+5b4
Up/bVwICYM1A7TIrMQPFzemcse1yReoP7iA9spxtiR7mS3PhzuFyK9uFrUfUd0d1
0BXcghCAitdrwqfGf7xwMQIxqa3nKDHJEpNVpRiM9XRalHSvYBecQJrpFQiEoFE3
LS7dfpUWhokCNfPItdNQAdnEuUTpsz0zXIPslP/b+SxrQXk7jeCdE+1C+0ykASoh
GZayXowf1VcQLeom8gRAtbMi4ooIBz3uZuNdYurgT9c95PSBjyzjtGMocwsHxIED
NFRz1kbYsRtFD23Eiz25LwXggk93v/DkRPBbTwWOjYJI/N+87n/l+YK/iI9i9yno
F3YO25n9nVrASxqSh3r3Jijwu+wYWdG9nfnOzj57F3Lu6ZynBd8mMeYoc3+F2TIF
aDh3qkuQXE4UeelDTnzPL7HP98s29unN4XaHdbKhi/WoEaibp+gHgn6Avruw2WjB
vfSvH6aQzGlAdRsz8ubisME/5Ri/4sF58p5uHZCC3KgXJpTDc5LkmkExb98+CdMW
qbFyng6mpTxwDJZs7qzsxteedRbv6sblOAzMfQzxw7bNwQmyQfJgf85/cyNYJ/Ba
mMPDi/b2EG4YPHKIfN6hOH0E/LKWxHKU/e2Mj+rNaGKGz49wKQj5FbHslGHtukSC
kTuPMW05UY6q57mdg9TfcOoU8sScCeZa4ZKzZunrZKaZ8cUun6AtwIAt2GN4mj0d
VcDmcALyg8g3CGLypoDZPEgmrhOlXe/WAZGZZeTLgAjEi6Geblx3kI3BqKnUWcsC
9tN5yOHH5EpVaeNv0BpHOqzLgWi9yBXDbyXPjrLRR93KPRsJfN2zCNvNivTxgtdf
RXfUj4mcQxKRBAaKmecvd6jBR8FyEn6eChQisworKlbZU0xmD+3gr6aIkcoPi4hJ
FquvgatBceHSJij8WxbIhchqmjSIg3NeCEU8faNRxjlsLQJkQ66X8sI6AucMXlgr
+VJZ66k4i8lCofLXY1aBBe6dO4irsS9B0d35WzQGu1hRZmTvIjAiB59l0mpFUqrd
Y0sa175oaxuXGnWi20dcFmqalIybjrg/ZRPJhgelCDgpeGJBrkRLCiJd6LsQ78aJ
sjuVuzhxxyamsQy95zaCy8UIDvWELz1qvngEJWxgGPL9uVNRO8MTbqDYi+4mNjb8
RvKOYLoKLSNY1RVvUdod8OesEbpCWDLp7f2FH+FUzIfZ7FgAluJ5/5nlW9G3ZRwx
5C7CJfU77x+WGFrjUdyLFjeY+R1X0rzUwVZ/+/VYQZ2L8dpu0e+GdfKLOBox6aJ0
eQE7tVSZyZfmZ4u/rZU6ny/qmR71dok+otpv/s5RyMrKHH3XdInmzhYYyLYTX/08
thyYDyfwWwP3N84LuhuLIVRjPPj7z1sA8rDBpIlnSDiTzLPpWffa497V8i04H3U/
wHG9HvSW3HERbr1si+rNHuylzHiHBp3ghptddSWprKmAtpAiogE8EtCs7jUOUpTJ
ShTMeWAmuUfSn9D+A9TtglrZ6ZB4NlLolop+oA9i7rLYZX98EOnXO7SgSi+9YhUH
bQV0BwAmFfgYI3yb2VWqMYzwxbNyazbXVXE5C8HhHdi7XfQ9TwyKYsMlO3Y51Rpp
xwvEQaDld/snNMP4UvvuZeU1kZF7/FnkTqCqu/GxWeIakWEfk+mAUCWf+bJ7tBS7
OLh2bzrB4GJbdkoGyfOSmORj0DVkGyuB1pmLaEkP8JJcFWNM0FNcE0juBRhg/fux
HdMq2mTZt6LYEgi81KEt/g==
`protect END_PROTECTED
