`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
emVN/L6ngDBgDazVoFxfoYuP6fSuwhlFtx9DkLCRtoBLtB4IXJoZnaYEP/8Ljff8
SFG5XSrQaIiTmZYVR6gUrflDTMM1q9oKfOWo31llHxCbkF1h+KGJg7uNT0DwuA/g
haWnuZfynqyPBbauzb5XV2gKD5EzWCIgHficFb4L3QmOjLRXtwIA8eQmFdkuW074
U4RkZZ2bXwiVFCNkCTH84tyZH0QfRtw6anIlImlIcSgAwhiPnt96sA9tfRS8wMSQ
0PvbiomMpyrgI3EU+lovkUKA32tEHgTDBtllDLvIoH6SuE6o2Aw9RKq+lW1pYLCo
oGQJvtgWabZxwX5UkPVZ0Awhqkt5AryQ15CQpBGqFzJjKvwYcx6k0LRreUmsouv8
7rh5k3eCixly6Y8TSONJkcSL3P02W96loGHKKNchO/5vyJO5c3STwZnaK2yWne2p
cQoLreZL3Vvj2XrWYd5ZNg==
`protect END_PROTECTED
