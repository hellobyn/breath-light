`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFR39iT/jjuchoCoxOw2edyCKl6vPHujVpaTlm32MVkRGG2o8zy490DNcgn6EtUe
fe9DQXAVGV8sq9wWH3RsnFBxSDOEORTaymgDip3q5ki9B7iNc+1W3CR1+JWO0534
9XUR+iqtFjjplVgPGcuDLiyUBdKqGvmIpCVnbx7DhHx8DLn7qwEXpfmtSAc65R1p
rjXCUAGYhDd1W4LQ1/N+ZiLEo65uIfaz7xoQw0dH57svBVSIEXQ2cjbW3T86wMF3
sWDW8YkPyKg3fJQhIP+hmfvn7tpudEJ1crwPcH87dx3K0xRGWM6dGmrBrELNr2Sf
rn9UhfZ84Ygm1aRH9tJ3Rs1Fk7teDJuCHEN+LcKRUrahyxXGr8QEL25AyPvQqLeK
73MlV2tJhddUAaa+YMWnwJ4X5nk2bLS0bsTWgjJz3rmLDdGa15OcRhLzKc+esIRl
RqwyB5+CipsWL4zZss3rWfpk1wyeGIuTjOhidd/yJ023dFlxxeklFb6UXaI/H4eZ
i8hVcRnci12e1FYwvsxNR2Bt+7oCPs04LjmJ1fkBN2u/M5HJam+tl0MEHpj7jHSH
JOZqjMcmsUYkNn+zZ8RQ0CR0PnP0PuuoWjczzKMZ9Xm0Xzr1wiFvIiwqGEQWWssW
esSqxvZkdDsmR8BQ/nHV9FaSjYLzdu97UdWRiQeU2NGwovbuj/Rv5esDI+YdWWIB
Ev6ZDuqLDV+b6nsJGWk9P5C9+Eto/wIZNB9YPQC9tuEfJIviInYvSDNTkiVfaDXs
9RUdm8fWGwO6BDX8ydqwEaMWKqJ8wTj9hfvtcvCt+1+/uS0WM9P/6j/ggrXFrEt+
sxppyRq1z+rDuI+YhomU4u84+7PTPvVhLNZQbQCH47vu2Vgok3MmAJVZIMs53rMN
3PxmN6Xr/sfbJt39uV8aKifVaqIGIam00wNfkzkqT8O8xz83XHCZRZR2fTSsAR60
Y0A7TMIT4aCtjLx/Exnd0iRQQ9fzU2GVkkWXCfShky61pHZEXM6JY3sg8boAzITM
X04J371LoaQ+x1Y5e8N80fsUna1dqgM0SxTnd+4mWOPfoxR5V9AgjnbICqwOv87s
qyvGmEtk16FDX1At+CFaXSiumuNwtknGUyA4UFnXgpEnB4nYY2oMVeeo4IbUyjli
NvUyQ1e5eH/2kEXzdALjowHhfYfiQgRrzgLE1MZDNUPaVs9Pw8Vm6byLly6VrqVs
rAWbM2fBMeGBGARrnECkgOeWubsp7VyEnc0zZMHegd/rrrINlscb/WWRKFws/HYs
xMRb98MIvp4e+90SCsIk2cW9n+OAvkMMmjaO9bzMFk1mm8P8p6mbGGry3GPpyE1d
X6CAGzoJm75esZ7CdQMaHt1exOlVSbgsontdSvcAsgOKZXO0nJ45IDv2ps90KK44
rze71K8VgAtaALa7YIlOeHKcxETLVLdaYhxrhwg7aWoACFByBacyuc7QnNGoMdrU
QEFU3lkwT+R28+TBOg9ExsEqMcZ8nCyCrW21d8WNwI46MBty0IAwCpEaj0LkJ1mr
dAJ8qbmLmFIgJ1y9S71ZngZaePFXliZxrB1pyExDNoWqXiX2WEx7NJl4IwF2Tvtx
CwOPMMgwVWkhpVbufsy3UYtGwppAOxoX8w6nyooskYdU9ExmTM/fI6A2XyKtvh9I
BxNFG5jCCiPbHP6JfRpFU1ytegEVQkecZVmiZJNAkPchQEIl/9frO1if7xvTKN7P
itMA4il1ZTFzgnLsOPLjTM/QGpjG/Z4yZmZcg9efwLQigc6Ajxei2V1mPI/7K2Af
2jgZ5/8zwCSn1gC8wZApSyJu5n47J2NKZKB3VwPvwAsnC5VbO/cmeP4GzDHxy0or
hnDWRsHV7ciNeLhEenL9sVqn+uq7GJexhK4gr/TsTQlJRYpiZ4r8jgWTjBz6oykl
Y/ZUClPR+mHGZKE1GuVoUds33oODdWm/3nvjrU7lAvzqRcXQydX0Ny5a8qUIo2KX
8CnMlRYL3XByw8i1RYo3PlieHgB4adjqR8n2/KbGIw9Za9Ml5SBV8A9czvzKwThV
RhjST4tno8mXVpx0CmH6Xx5w2qSQRALcRr56Gtt/tpPLvICCOyi4baVm66mbwT6u
ULdpGRec5ItHN5WtbJ853+U1RJzr4h/FhVWdYCcUiOd+XfuiRyccNgAOJzRAaO95
vDpnR7HpfkJqArH4f7ZH4niQhEOg5NwnwDP9l3vSKSDcHuylzBRKEd0ke93/Yl1j
suVACfHRyuEtv2BEqiRNPOo/6TbQjb/VqbjXwfxwm84PVRfeBwQNxNtjUxDmvuD6
0e8PZ8cQ68zZazxui1Sdx0s9fP8D+r/KyDF5N1gkXKfMeEnVVXZaLTdSO9h0zF+A
cgAQyQJOPtIgqaMyhJjvIO4eMWOrtilucDFA2wt15eCK+lFrzOeEeWJk9+rQ0iTY
iDfqyziKRQ94JCHi3eKqF0bw/Sqrr6IMh4UpmbrifarlwTWrAKxa2EvlgN+IEGCm
jhmTgHg4UxNDzn6XHaVJhFhXGC4nbzxGj/ecvagb3Macssaim3zgrBsESzhsiXbA
XhBKNynS/AcHYmFDolyj5u1qRBWgNHEZ6/eK4OXCjirch0Q/q5Sn6QqRVvvfw9ny
yhydw053TRHI33IEW+IlF6RikXxZWxGhF9guKE02ferEc07MsHZeFLAndHf6ZZwU
u5r7ELAUJPgtn3rrIPSv9wBhi8jZrTQwfGImxqB7z+iRRNJxGkBIuu9RsEmE3d+y
9w8T5ZfZhQ6YLniMSALRq/+NeCW1STSy2mOT8K9z6Hn3nLcadkiu2vUGwBf2ent2
ZdcGTGpbZ2wPoCGbd0y2znjcZ1TqK/scUYDZAUIzj+kv2hgkAgGjeIQyZ6N53s+b
PW8rxjigoSCAL3Uo33i/6hgsvHo5yzrYUN7zWXOBI5N7fVRB+MZwOVX8qs7upvMt
mnYpWu2ujapLZwbrT67uIhWcZ+r80xoy3+bQ9GkhvUoe6f9QoyZndsXjiJ/ty6wP
dRRHCBj4d+izwc35OuPWcwVubKO6Tu8kzk66oEQQW4TCzR674QxEkyNGtkW0Fuey
Tufnmb+GYuye3p1sTa88qQJAXparXE6zxFpydiyl6meleVeoYPlTXsWmROfP6+Mh
qb2Jfu639cIkhGEZMOAw72J0RggmTjxHURpxR0pG4GFLSSQgwyCfmZ/xzeyeRwcu
VLPaB3fAWzA3EKe5nZzSUZUcECybnmpnzmfI3coDy9TF2LuRvbMjUAjNyT9XcWJs
WLegbuj51zyWw1/7ukikIBJm8RHvt+WpBZjSGBhYDuxqnhlzEJ0gfr15hw+eYAUu
rWAjbcCq6dMwe65QYowX/HjLDRdlNwsvEjLxBylOR1bNhquh/86iMnTJoLnH82s0
TW001Sx1sbKcWy0EIHUs4pf0EU1AE1Nkpql32/+ohixPhTxEQflEaFJDHY/suaZf
tApzjX9ueS1/o6yEdSwGt8mliB/ES6XmtLD37YKGxacWOwCz5G/y0JyZNyYjD6hJ
YcwL0kBPiNXgtXlzMp03/h8i5drE54yOghDTTIAZ9CN45lVx9iHVVnSaxVPI/QBu
h7TawqZoyzZ66hnEYKY80v+UXZaWyr+4k9zBs84gXxNYOAaRJCIokscQGVJ6jOV5
cj4mkoDcJ67Zt+eNN/a3v0F91yBRny9uY1zW51mqKmdCG/8QaSHPtwQNrpWxvtng
`protect END_PROTECTED
