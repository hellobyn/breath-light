`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73gwD63hTsd0KRBQDxNxIVVmWG2hGHaNepkMmhAp+wrJlrmKTuKRSq2Dar5KtAZ1
O/1TTowvuDXqE64mIKOC+ACaEdoy84Z767PyZMwPQtTHtAS0ZTEDnUBM4ucf1qwz
LcOGNNMM/tZldutWOOITEFuPtVA4Opy/npgi6030j6z3n8WexjugB9iR1MwrRYF7
1/I4UbxQnefy4ef2zNj0EiC8nJS9JVO7XlNBFeh8gjbEYFPweOvSq5VYSffxlgqn
qyWCl4dxdQCFqUKMir+f+bLmYzcU0AuNlCfwB7jOuHb0UrNGQY2zGfs27/QhyBAe
UtCuybyrpaOnVwxm9YHtNLTpfWlHdDcVVGdms77fOjTRxXKsdKc4I641Fd90ebNT
5J9FrLF7NLBdrYyRSwEpOb22cS6iMlKQXwz9z6Oa744mHbpuhFJyKEKF1OrCw2Sh
D/fuH53N/psX76cKA2AhcM4+RJ8VoTn7Z+D0vPaDa/0CewNtt71R4j7t1cwBcNPl
a9n0UlLTwYqarAyG2FQmMtTesA1FKEHucvu2KekqAhw0ENB01i8qqhYtZsbIsGsT
TWXvinPHGZsq/Gdcf4b0SSnOYNlkYQ7Eu6bWO5/KD3O4jGUeQyIBEzO8AUMMhpqC
b15ZrcRU1zRl+DTdiHjlcHo+P146FpoV6PzZo8QFxXX0mePe5vT7cYLwjEDY3aBR
cYXNEHWbJxzFtDSO5H3Ss9sPHMc868u0AXZTdeKhHIa14uQprwMvR/fCo8zQRDxU
1Lth2EiYbp3k4kaZtQN93cTh+dVevM1JWtlUEgG1bTHfB7mlQhbsnttifASqYYJE
bOUU83QYH0C5IpWLGi8gmlI+JJf+EEdWZTQzVL/sIhD91KQt1kUojvHfDo9o4Xjx
raMooYCaO4y2JcLTLBoQfvx9zRUDqBhJmgBA7acbdYZLWa0QTJ/W74nYMdez97ko
OEThAFkEMnWSqLP1kQIaQltClXMqbzQvBQB7RWdrXz+E4Umy2ScUf4b6vdV+OOVz
ZCLi40c2lL9lfTdQkS2KI+MKTiQuJrklitO2K3vit5wP136ENqncEjjGFxtOnAJh
P1I+l900w/OMIG+aCuBXEuH85nTDSBZcrCQn66pfqgyOPAodOIDIGKi8zfHjKMxg
xInmRk766BHEucZroF0b9I42NYpF2mmcKd0kze3lig5YXK50qzpS7kwm/g70OssI
RkUlmFSRJyUTDOlzwbvFMZBB+/+sx6RXawcGsy+ge3C4nckToabyl2LGmAPzrQjt
GCGFzFSeXdmZvJajDgeqP0kzHn+us245jAIphuvY4YIR+W1WXZAU8XHVvqAusrxR
TzORTsCaQCYEUkQj7M+JahbpiXUn+m+9ZSikEXPM4KpVP3Ibdx+4Y4Utz+E5fc9r
U4Q5fqpHRl6KUVT7A779vtnH9TRTgvjwS6sodfqG5r6r384gXNKgmsLOA24XZdIF
`protect END_PROTECTED
