`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qlC0sGZJrXnuSy3v11rnBTKXL5vHBtKQlLtgXBsNr+DOwv2k767b6R3Ml17x5nL
I2YgIgjdf7QpC8JY19VQQr2gzNq5pg4Tk9pVsKOjK3AQoJnMNGQw6oNjDYjjpmxY
j+3GlW5C7+2MnOIWlbSdWiRU+Gqp/ahtapcMvHpSA+g4U3EMnmiwd+mAQJTfGr9x
tFaUxq+h79BlyFWcPmecmdV+sc0fnmM/9Vya0NIso3ygwP6Ew0VFRpeZgvSe9exl
rLjqY+8Yx2seiEGSeiyGU/liiv0AqzWiqSEEmQbjNPM0TK0S8V5S3KgiUt+gltQY
B0tPF86gKgmrZkfKhlDE2LQfQIXLPMwVgtMpr3y2vAXmXZqWOePd+c4j3FN1Tx94
DqLNbtb6e758MRggX6TQiVT5iUojt+n+qLd4ZJtETH9k6u8CjhIl506ELrkUuxlY
ak4GTQQrmi6wVdQUGoXphWfV+zQzDI6uQE0jC4YSwhpZshDLqP05noa6fGKVs7xY
UWwPUzafEz12uoYejFcPuGX/ZNc/13ZgtXZT/ZDhJ6Bms8I7pBktGXuNzIkacOpC
aMN3pV3gDAyWYcHrWcb4wkOrJf7RShZqplktl2j1q7ncDw2rv2Vt2j4w9aQ2TRYv
M4++jdP1urnR/lJJe3k2hE/wrlndYemkGnbF+atWtYUBP4xLcB2r33joepYl5Aw+
1+/7TJGSEIJEfP3baOUWoXrz9RwLgE7oq7qKdKdmKaIFKZCINUGSSuzXV3O2dsma
ctSa5NPRZpSenYteM40A43YskP4VooAigjK3/KteQpnl3e/izJVQD0vhgD0+jaOT
OI+2Vn/BlA12B3EqoaCV4/yb+3RwSkVOp6kdLa81otQiB4Otzs5mFIAR2ID/wVXY
ukdQjjEzjxcOrpDiTnuYRSc2HStZznBb9ZAZE7/LpNND5o7hj+FDVkyghh2bF4GR
X1cDNC3+wLuYBICDXgvWYNMeOETAAkws2l9IvyxdVh5vshURBISS+kjZH5F7eCpO
mqH87Gw0eht+EjnN1DoKBBSV7CyK14Ahd9NtsU1v14nZ25ASWOI31bVW8xUiZW1w
uu5AjAjXwDEssOk3uLbdUTc4wNNPHVfipQxgXn3blpm+WhrlTomggu1p33I/8XPj
ngVPKt+2PY9t8/hZ1zBD8DR1X3eM0ugE+/v+TENgWU2TSHX5x5mqt05qnyfY7inG
RobeBTRurKlZ1m58dKf380Qvawi1BrIMWLs+SmzB7EuowJqi4pXD4gQu7wcNHUlo
fypCmH53w+Vicw892Kla40PlojNl92XnXi697Qa7lE57wxemUW5wbKWOxv3j/F3x
ZCMYsR+JAewcSMvuPXbLzS7XGcm3iIrGopoRJAIlVkBzzLwL1Y0GryMGbNvK+EiJ
H6JDM+zbdBbIlzS/p1ZWbXtFbZ9GOurr/QFtfiWqETi7VVO/qvybmg2Kn4yBQIy8
HUCRbjoIo830KfIe+hVkzbPtCLMeI6LBZ7sdpJ4bQjO8zxBn1Lj/99B0nY9kCHCo
kC/ONVQkLoBhuf7hk6lViRtMoTxyYKJfF6gFb03I8wTb0mCaxKUkHG++xmZkiyRE
rtMSCwSOHTeFwpMsyWD3ZGGs2kHdspvIcWLZkQSxTYd0y6h6gWMWyHdWGErfgNft
33kWdOer2kBOaYIX4KnUmx0Bta44+tRHExFBGTEVzmozPSUW5HfbkZPmBDTrK7ue
IOa4IWqkxYzC7+Ikv/+9oClS1bKhLX7jIj9adNM748iTAa7c6oSaviUeuKjPMsZF
/U164lGwkNUAlc71EDQ7qxKa+9TTXqsdPP4S7Qn8kX9Ak2UYAwBXX8qDWRPtfSFz
PWYwSGwibfS3ky/Ft17qXkzkaikO6K4DPCgOnmeLdcwsWkVDudD9qI8JyvsaCv8z
q2+nbIboRZVmXWmCHPaAcxKYrqnW6tK14O0ZI+ih8AKand9BaMlhsJtarAiLppkL
1NDVpossP01SPo/dvsl9N6b9xnOqgh8DAjxn7mVD4izjAXxUphlQKIi8fdNQV3+W
Rbd7HcJY+coUYE3tscurzR8tvJ3p2+RHRIPlRVYzp2vR6T3cqhQcxKws6CL3KhyT
2Ld+gkyYrS1SXgK/O3Vu8eiFYpEsFMroSVAeYs99BekBChoccrvDPbceXSTjR3vQ
G/tW2E60ukb/6sNNAmY26DpRKr4FBPcWMBpcnegSwTbJMtc8DZ6OpqgLl9pX3qxJ
zhospYWLGIrEci26CveuzkuCCNHikl7S1ge+wDKfH+I4K044vRYRIabkgDr2c8bw
qp0Q7+cmQ7m3xprpJRWfvpc5J+nd4Q7tQ3AAMi2210tq9ieC2BOSdXVjOJjTKR/q
9F+aRH8/lAtziL46NnizaJ6dCPM5EEBBsVpkWbXPGBGSGYvtZmf29fZSUoDlwCVS
cX+MAle3NfUm97TqeDIlLn7JnuyHHbcE8lli17ycd/CdFhws3enzVqUjlFEx0j30
7aZNK1vWdibGuzI7gvj0eVJUmg8X6JzLYehYL9XEV+dJCcmH4KRqrbwAN/pSlHz7
41OVRPAmoWZy8ysI/J9rl6umb7qKhh8AZAOIcoTJAJ+u6eyrhox75RX8p5cXDI9f
nBl6R2EIoHw6iQmhWQpPTbkKDGX/6i+NH6Mv2v8nXxLYYhBncKxuxzudmfKWVq78
UFeh96jyFRCbSNrzmYNk6+dg4Jvsf1mqIm49lbh+o98RGzTzwver2XbGzIoMTZyX
e/9iF3W2MZiGNYGz1lZQLad7Cie3IeIInEyatVc07wa2ndqLssemi8OJgPwi9YGT
yF4LyHuZiqvpTG9n4Fs7IRnI7oCWjpbkQf5fP650GrKfgRMuV0Ox++E138OKIgsC
ny/wUWq/UOaCFK1nfHB1pv2au+AgHVSJzKpmNfmX9K0kalOvT1BIx2exm7PxbMkU
4g1bh6yU5+LWLTZt9G99nlzqe9MZE0UTk6IaSkWrfNxh8WJDgPzSL2gS+lyhdk0y
t5CW8aAIfCJxTYLLnszWdq9xPKiDEFm0H58O/C4FodKXVaDCcFWi4RwBWagghD7u
j25CcO9Y4I5G6/Xx9CPPIOFVca26KsRoAqx1TnSb+5tDrhsh6WzeOoa3pAECOlSz
f1MZyaICQgA6iVVEEeYab0KTZWJQLI2ND+g8l6ahcoIPATrJ3YpLMofcSYPL8P0t
hPZaOxrKX2WPe1LDvWmY/i7O8u5cOPE2k1zds5MPTEywFKhalmqblc3af1qSewxU
RVd/HukzgpLN1JacpNS1QBMZiFSmWwd33PpMBWCtnxWpfdbG5Z9GDHRZ+FNUk1A5
6p9M53NY0Ncg64ua6uQxUYf/pie06S9S8pZj6wo4m/YzIoCf42bLBm88hMGaM38M
IIyrnqS+NHEqUiiNAqlIQbyd1cNyHUO8n4ozhtc3atH9Wxcow9C3wR4J6kyh2Lye
FaFDZbXXBhdmF58DIWHB6o5nlDb/GCCJYlPoreX4J477CzavSXeqsBbgIYqm+EuF
x1sDqmg/Y/MZTkaK/rEuhc+OlEWI8NpDDFl1lzxqE8Ojhr+buq8L349Weor6tcHJ
SUS2A8UON5yrBAOzbqNP30Qg341Eq+mwb71OMEG1G8noQ2XJPrP8uae9Bikv5pNZ
8VpM7xlO5pawErgfXn8AJ7Ho4BjkI8i+eJSnX9/lJDinpuzTOOycFn4bvi1tHjv+
jwOA0C1FWnfip+JPVHEQhoq4Jck1Hj441SxS8aYwGsLUgdv4mirCF/zTlg4i3whp
EZ5JUANVpPabcOsCt9RoOVJURV/gpVikXxPOBUqIRCId32SMJJajHqoOutJ8vt21
DDNGZkEEGJKnfJuuqPdCzVCap5frQHJXZCwc147Ov/h/RrLFPbpmrToUoZoLJSah
pv7aWXIDTR5TsC5nUFI7zvVUPIjimio1R926OeZuFODKuRBXXWYiT3DHVMs9smK7
TTmida6Aiyijk4QUM52BB90c0ud1YeA2rKvZuV2pUbGlXoaXQDyN2ifvULSv87mU
hUWfgW0uusaS8bxnJiLinYQmz/1lIKm3y1YwDtfj4n5uz0kd6rjcvOSOEZSqA4Vi
kjYu2ARPk3Dk+cE9q2EAeyh+TmHA64/GspYsc4IKrFBU+WKq9H744HzBKRdKxWDb
/dniQCQp/Mhm64G3vnuAnfsVkg2FVDsqlbg8TqC9eJlh3BgHIQD+vDN1VbziscaB
Ctp3DOAIt+sxqvts7ZYjqi3f8y5I+G0n66hzWMiy4OnEopo/zSDVJLel9SMvGmih
cj35kM4lhtdzniKdHmLsaESpabIG4eg+rb63fjF3VlvgM8ZcmgFxuoy0Rv/t2GW4
N07rV/tiuhidmVm9DPqvD37ON8z2eWgibFKUgoZe10NkTmlF4knFF/9UkHjx03tA
ewx3737WkTtgd8zmM7HJcYQ6wL+oF8gULz7HQl18WMTp+zCB6bRJ6xuhl/RmObAB
WaFwIbC6z/FSAvBv1edkSZ+FHRRRl906v2qWnq3rNg9/Hkbv1lENdPFaYy8r3/GU
BPaLOm9EQG8SCQDmynt/a92hcvTSypJj8xN/i4rInEv0L4w8gIAFwPPjlZyiv6cP
dkV+0uhPtBvVW1RQn9ZINZaqFr8fF0w0r3tVKSqz8e7UQ8NeJF8tvv3fKZ3pJfZq
GbLGcYjQ+scjBmwPkowxnlq+GZ1fJXAhhgnJYRa2hCrkciSRIabzacoUAummx55J
vThJx1hrnmiCH6OjXC1HO2Y9d9nGAxd3KJjzPeodjO9U462S1igXdSRbQ/uxr+58
QI7Yy/CrgaTJumNul27lQm7I06MJN1MmglHEQg/vguSaQdrFSHZ0ZoJ7nUn5UfzV
4NYJYbcVObxfZIk0AL+DM7nG7FytoXpyiT2jlosYUFr/9qt7a7KXiJKN0t70VQ01
MiXx3xd8lu+hoZRHh43mRK0TUzlDbsFE8EVSueKPAnz4/Rkt1t7n0zI4T6q2TJNP
ICjRSNFREl8rXhpDd8zLZxd5XJuFI7wKEXcQCrVV0gFYTXBaCAz7tFCHS44UW47P
q0f0nCD6XoaBdeh8PqnlBSXO3QqVm8rxpdh+GW9UjPNEgBsPyRqN7mVKS9XF8gDr
xxhds9t1KICHGiXW9+ygCL8R1MohJWz9hjmzeL9zEaFIqBD1dwvZBcMlGH0t9pSm
QTJiMjlXEoEp/1nsRPq1arRP70Kae6HwfuOU5ZhFuaj0r+i3rxB/x6g1PsLwcNmG
uLg71TmFBYdSh8mL3T/kyQMARJBaNxXgZxLeqMU3SwR+UTenjl+A1SPLg4pppvK9
k72dpKcrOrACQPghhjpGRHFgTcQLlI4MVVds9+OPz5f/P4hHt46zLzU1bucMM9Hz
ITMH6WFng4Wmf0NCAjbXzv4jpOnm5ErFtbPx3mdQN2j66qxF2bkTwt7TzdRHaKhI
qhxm+4AWNmO0HCSpDgQ5smBMNDjcrNAo7Q/2hYig8K9P40b1j0IxVI9gVcFPVRon
r3Yg6q+qx11LIe5OA8umA86Y16CRMcwJZ626wvtfWRJENJc0UrCn0F6ritTH+LkJ
iUFzJSm/SBbD9qM79z9yPA6GGLUMH6QVJxeYgbkhqmfgoFHEzZRLhD9751dQWccF
4RhL1rcpyyQbHk2kO1KIkvh8Ww8pXln0XTtuRyGfhxR+0/CPXsCvt9TM7wgpfO/4
6OdUQCjHLN9ugS1UjdyMUHE2cK1gKjiR9qEJ5utZCPtX/udAyA1NIEiDyTpzNsLS
bujWV966ZCI/+ZsPoQGIcEqZfY/HquM5XeVF0I33OTg=
`protect END_PROTECTED
