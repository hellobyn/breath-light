`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seF3wnQuD4k/GxSl5jTBh+dcMCwTGBM+OOcmJbULdF2R3Im6GsKpnEymmih9YGa7
bj32pQCxYXm9g7cFo+eiJbqmgw/7G8EcjcaxKhadRkjvr5i6FCaPTFEaoCOBuIiI
2Z688bTsaHrs/MXzYbRoWWGDLwswZwksri6GHR2O9jSxwLy0U/nNCVPZ19bVzfLV
TrdqT0DQdDc9Sx495vZfGJJqhJCTQZenz/fBPN6FL5cCh+ZLxyKgvSWcYdDdlCdD
keWGka6Zd26+m3sF4KSAM4vEca63VTjB0kAdN88MXA26C6nYQoA3Gjg8nh7L06g6
EtVS7CWekILE0c96/wY0U7pvzOs/4yAgJINiPFXMCw22akhvOjSWMf5ujjL/dH8/
PLz8s5ZztemvbtdGcUTE+UDfCDbfa0e/6deXUWzncF85p7utw3y3YBv3LlAGKp+q
99oaF2h2oYvKpuC3ikfdjgEK/eCWNWg+MWtmp8cYeR7wq4bwVUSm4OceXQmSUmXA
mfUEipl0HCpZompxZRp4QjDxiPkcbPXiPMqAUkC7k+mAJNii6rYJTeCEzXeJSse7
54f/J2IWAjAt2+8RHSgY2Ujr2Rv1N/aw8wMYMWYUrhUydecQYdo/Yn2FxPHribzP
awlKdtsb3wJukcdQhaC8NCI48SatMdHSxkaITzg9vkHfrigttyOwjqv4jZbgLZ2t
ozAmno/TB7knwGermPELrF2+2g8MxBll504ocGML6O/V3Eofq3lIoiFEtUFq1NkO
DOHZuM3TwR/t6Q4+XDz5j2jpjPwXPovuovp+vDn/fX1dLvMCy4B9xlHFbTb8y64O
VTPZVstQb8hjyLIcQxrEhtBFWiAM5imjWPLD4Vxa+idnetYQWeT/CfZMhsKRbRsu
3vM0S1E+e3bCHTxIa+P6PfNUqTYKG+eSeEY5Olb0owMlbkv5Czi9Nptkbv+4rPRl
qVpSO5xUwiXlUzCPrWIi3KpDmypOKMw7Sx4DQL3XZGWfQrqOv2umDQHelDfMF6B0
vYvN0hngntG3oyGc8QbWiVdWOvRaRp1nLOj2ltV7k0EHaMxX/jE9VeO9xDkgd/tU
KuEtRl90CFetPaiQGHKi4lTpG5ZWAaJLrob8GULas6cK1AjxFkLZLfNBIVeLs/er
PMnMK7tTGAzhcdkbagZtaA==
`protect END_PROTECTED
