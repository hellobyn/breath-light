`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfF6BQwU1nQVWEmoY1PDBlTEliWRGoP9SDlvieSFIYXGgm7xfrYTuWftggg8wpcZ
0voZzTJcAdMjK0+lptqVPmt/ZTrMaq+MigAeZA20swFk+sqpqHxwCHVzEcjBVHvN
R7+oc4ti7iOsYEZgUmnJO4IqE+zTbrEzxhM5kD0bLPI5AhcJsyYzq0/PY/F9hEuS
6rAxLM/YXFSX1HU76ppVg2033i01HRikNhtCIp5Ejn3va9Ez7G4Jfu4m+ghKB66C
X0MsPJz1Cv0mLjd6yOiTOJCP0r478PYiUtteySnPkzj51NbbM/lHqzLg38R0Fs4y
KTvOtldStjok4zCr/LQNRhRRvrnrvC1Z/ttesl+as+/9bx+hS6Xi8BM8+fxYGykk
kifRNiJCROubrAplzjb5T1fKvMjy36Ioy9mG/z2MTSdzacyfUAKpUgIPi4O1K2lA
XLtVO9e2/AchWPIGEOnLQt69Akmv3lP/7NYz3ytOJuMk5CT0EOVUBg2cp5wqqrAK
nO/+qKrJZLgFBEOBO2pgGSj0UbzYPOuUf2dDVTRFtsFlow8Yv5kIEYy65ospA5t1
YLpuBj5fbaGQ6JS4ZhSd60m4IfVEQxVkGVDHHniyI6W7kYP9nszzGrq9lyHTnb+q
xSWxChL0xyb5xbGiU3fFsnooVB1qRzmahLev2qo4PGSQRTCHA4ECMgf2GCvme9hB
lT/kbp45SNUnwD4H7TXT+ko2G5X2/KNRxT455CAiLRBWjlhbYRg8qpvu+pgUmYu0
WaCJLdXmPBXmYuwui1xNDU5y/dxzy+VBnJTgUJkFTcZRlff3vzS1hbjbURaxnVn2
n27HZcX219QUH55d09C8YTg4WLgrqtfDAIn6fpfCYd6eqE0c99mmfyrp4hd0zM7m
8deGtjxLgEmSPZ3jAMqbUcieyE8FQP388gyhn+Rx+HqmO5qivhxBh6mJG4JJsgAr
QvlEU7FPsiIUW79cC+iYapoBapQkyiVfcOodFC9wtvI7+Jgqo7aaZWKyuwjIXJj7
G4ZhuZkIFiGXj908N3ZQlz0uY1e4CcgNLTLO+URGilMiKFv4yrPsfgX7hkIdqXgO
d2nXxn9HH5o7O/hjb1akpp+24V9g2vhUw8OF22vxCtwNmTPd7bCk5IouEBUrHSXZ
Y+fd34NoNDzN+b57U8o0099ArNUK37gOPF6Ka5prSJD3hjc6iB0qJfCmx2M7zQcZ
HtLXhL1GItefljMTVVgzvQrfcStJWRRoaZ91TlVJcp9l8md0s8+dIE4788p0DpTh
ztUMuFdJzrTr8Hv7QJcQRTjumekxo9ZE8ZTonQdEKQj7SiQI1ekF8h+/fvIjlLXh
fpS2loeTqh0rtL7jleNtwvIhQUnxxIb20ivCw+Ayqe+MIOQiBgjnQPTgGNaPtcy0
NkauEx/W9tb4GJYpB/LaBo8oaIL3CAnvRaQgwBzwO1wmpwpWb3n3u5rT2zSr37HB
Xh8KVRV7IGYIS7hYkWUdh5HgSQOVEXXgiKvLtlhYf3HMtYfRr4hlLEV03BDAOk2O
Q7VNm0onj5s1w1E3i7MfMk0TXD2b1JNcoEvmMavxnSGfeD/NGvnsE9DNHsBnvwi/
mjj5o6Tdk0NDeY0n0fFZesev/4VzX2nlHDcYk5EfVsYd4zksfIAMAdngQyAHdbM1
fSwhoo5xzcQF13l4TH4l0h12YRQnFq7FEJ/O3yAgX7Owkv4I8ddyPB2pSITlhZvb
HLLT879ZTV32OHQXQneuxExqm/zuZ9EonQiO7hbbixA0nzOJkCO5LM43YQMnAL52
yrASPrAnFAUdYFWJTGXsCydE8BTPI2MJlHaF+GrgwXqrJ2inMnbm4aWrVHlkQZEO
M1lbAXMp8HMeIECZJc1jGuyFdUIaFVFQS86yuIriCyz6H1SPddd+w7+Ae4qCdgWl
wmh1gIiO/TZ8LvL2TL88XWLFIH677g5uRXa5e/0A4TZQYxah+S4WolXmv3IAlxd7
K8baaCt4eWr2RX8IzKZH3oWT1J4AKYs8fB//g9kVZ3ucPkrfPlmyEufeDuVOe4ky
HxxDuq7aqlFsgN3Xeqg6DtFAemCiXBarjTl07JR9xZ7caWGuVLaglKn7GdyAKXoH
7fkL8cRb2fO+/hvjHBs1NM66vfajIN/di37xmPFOtAReyaOlg5ojHfJqYNM8rbaT
M2PHPoS3DjagxuQ/ZbdAkEV6Gg1qSz1t1/luEPR+4ByiuA0vf5JP0dwcMV/tNHdJ
STQcTf8PcXHRRhWdaHJCOzjxYeQTQ2GqFOPoDSRoeYwHiCWywkdSOMDyGqxRhfKj
ytg35J4bLqnQFLicQb3XVARLbDb/ukEy2WeAbRWn57+GuCAXjyeSNp/9CSxS33ie
ELt1WOY0AUenc2K0vW51K/OA/7mJBZqik98LkDBGuqFzou8Oh98ghTK39chpoU0V
CarPHt9E98V57dz7MSTqxOqYO8SLC7l6iPJoLDmew6D96RUQaSzherOfctywTEw8
B4JEnCbx2zcVrTIrQETLiD9N97CAG9jrMhoLl5nVT6zDwX7EqODlDI4wz5Ym3jmQ
GtKK76vuM88y5ZuIrPWXoZJqnsbyL/F1f4rbZ0AGcYpNhTFDJoI9vct5mHPTghnB
cfdfooGSFge5z2Vu0RAw0UMtuu28SO8ZtEYQ0DSbZKWS02qXXhT9KFvnhvmGQ4K/
OxOwTaTvYHpdnXLaDhgHvriDG7Q6kscCI3n7sf4vpnwM7hBNcM5nVBy/M7nDPZij
OBUlhvqviorni/gcE2gObUbt5GVCT4ueW8uKyynrXhuEahYTs1x23FMeSajxwGv3
sXSZ6+hcBlrdelT+keE/aIynAtp7k8hsABD4TYBzOcUg+o7VJeQMHToyU48G9z/Q
v1x+0c36Uae5zH8XH8q9ifE9rR55K4vpYKwCBjTQqbdETZ6Auhc1kON68AyrdIqD
62bIZWjvxG5wCUnaAT7eEklLSkpnf1At6AMLNctih4BXrGyP5I4aBaMWzsLUgmkc
jRxViKdnYIbF24tm56N0OkkoqsUWq/g6UivPOK1uPwMyufKCQ28SpK/49rUXxicS
KfoMR3/G7StcBnjtGFY8VQ/LFR58A1Q1bONLupCKNzxGOMwDb2rE4iR15z3F0aJq
5zujcSH71MM5ynijvf2hcL56D33vIsdLkeIXbMRKOns1170jRYPDfCefWjvTrYnY
VkMQ1ZSceLnsh5hnRdpdVVU4rNTWVx+XKrlEYBqsZPtX7ixon/LAqTHRCPkrfzjn
aC5N2Om133jsoSNIhC4x8MIgPhsdRvO1RJ8IrttEk62c0xLw3CdkmRaBONekhd5g
+D0KcXsVr0LyK9jTDKzgymIe/FlOftZQputIMd0EXN+Wa5Xs/cjnZ7oh/PddjCqa
K9xcf/b7gkLTYTCT4x/J7ixjtILGZvyIVi/tLmr+vIeixtvEn3nuZRTcVgbgDAgX
RJIQtm/NlwnjbHaSq0w4s6INPEWre20I0/qWycrIooFtBkd5bpfrk5i5yCUNuEGi
DD3HV2sTJNoyYutTZQt1TMl7U8ShoY/U+Kk0Y5Xt2I6bCTaFeKyNpq9X13bKF0ZQ
zg9vGakuwzKCDZh2UEB+MhNosOaIT3dsHlgiKoUPa1575HfTvfu6gKAEkDHtBtTF
Iq1/z59FyocygQN4fS7io+cWOAI6XoymUTddZyUUb97XaWhh4mGybQJUHqxuBIlT
WNevh4a6SiCwwZJgJ2LLjeb0ytPE/dgSbvkbsO/myLpFXrgli//qYzGsaZcZTYIc
fByAacjLmnCeLA6t+40Houg8Qr6CIL7wkoMEeGmchF1yc3PLq14ToIswPrrCUo5J
D48anAXFMX1phk8s4nPH80hXy2vYvgJRDCuhOd28caL2syDVUeZ2MzX+XePntp8e
kUrMe0McUisNYdLJLsAJy5+n31LevXmW51Yz56ZTbIhVWmD6TTSfpgNLPcWHVhNM
stAyvpehc2cbdMQ6DtxHXkf5rfyqHe2fMLFuB0mMkg6av/Tv52oWokENoVxgKD4a
7VXQg6m22No6RzQnl4eLpWE+9JXsLDp/zQSPjvmC2L7EMDoiHuHDLkWN5CSzDItA
ER/CZUEhtBTSxNAt7xC8oUgRIWUX9IYhU3/QQDLH2Kg5Qui/pmGc4tMi2CN2GsnC
w3sZ5A5SzJK5O56HWHa5gQwLPln4Cg8p0sNFM5zS6Z8gUVb46yTCYjfhZylPsn7F
QW39HyKQqO9ntnMZJVgYfBOnnWFE0d2q22cEtceT6uCK9fe5jyVinZbT8ggdDy3A
8kWsLWlKHksPDxN0vvn5eNnwUXoCcNlOssWD6AblB/bD+loNrr+4JOJSHYeRwqC0
WHNwrRwsHfFsbrQQ73rWhJAEBHS8cJydVXpD7hy5lYtvX6sRsnSYmLhgmYHvCrBs
B0mZaBK138pXOYQXCvh0/AiT1R26NuMDVJ11fV7dqP3huf7UmgOx8ttXCfFsH0vY
AzP2hFalue1woicBGwwAM60xNRvy4TchSln6obDKRh492b48SlwwDLDTulNmj830
10QyyW6kmTdfrRA2EzwgKOz/K/2A31+mwDEO8Qdu62WSoIGtle05Ib8Hu5/sCPJh
IshPdmXdwGQVc6zy1L8YOXiaIhKPigkKIUrBag+B+MaS0SnNU3mXcrls+BdxTJDc
7Cl1l4daLKVKdcRY9mCnhIETuiYWHb5Ip+SpZvFAFUi7gPjYfJVeWmXf3HKo1ejS
ccfmUdvMhwx8Emu774oOefLmL05Z+/7qbCfaVjGybunAkPBJZsrDp6eAzYo1zPEW
v3X1ljRmNvpsrpvDsyYjvOqhcNpfLKqMjbRX5XqiE+7W2j9H/gIxwtGcqcX/uIFj
tANQf9QRFgFsQv0eQP03X92clom5mHCcT2ppEK5748WOd9lCwpHtnZiv+9/Stt5H
66uMWmx4IcPEbcP9cf0zhpnkjI/TouQ4ZpshgbgbMqnVuxbwNntfUImNsq0Iw+4X
s6x7PD6KUvouF2OA7hm84H8n3aCtR2Sc407wkonC7bDAT8SjI1HWrCxv7L9LnHFd
TINX+9rLJnbCTNUX9ExPOd5KH3icT47Gc2yCrgx+00xf0rEkzVU41uxfqd+joNCt
fp/+f+DPgqTIkhDlEZwWEtgFe9G2fMQKKAgCqzGFiWoZ/l18/WVeqld/xY0xXaw7
LzvM4go6DTJoUuUhxdu7d0pZ7ENKvHb41RTk4/741bTIrmT6dxH1oTdM6dYgsXw4
XX9zXikquX1WuWeAAMRQywXZoE5pZ2+l0OpSpPjAlRpayg/LxUxb7iwrVRCis5xP
1VTVmJvamhZKWhbd3p9nwPPSd8LcPCz/Nn3P+F6xvqZhjPOeUdpS9XU2c6aFAoUy
r+HhWpKa3GdzA2PLZqXrk4NQD+tpaRevkDqQrULxB8OBLCzHvI8tSYSD++mXfq8F
M+0DT0gxp9B75KhdP04/80R1OuFJW280qqDdzTxWZ4FRF8pptyTNf5H87hTz0Tne
9kYEIWNWDuci97TGSy7XCl27igDkSx2wMPYqI4lZNWfLpg3mUC0iTHYFPcXK2Fng
qYsdYcGcavsb8sAh3O5AzYIRLVidoWJrU5R9r8YcZbeO1xeIwdX3qm2sdj64fJ2F
89nvIUcMc7QVmPwG5y9eHKwb8H1s0vxwvSyz/h6y2/5MV4oQrzyGRUvq6Ky/eB2+
YLSKwMQZseUPQ5rPiaAEzR7tBoRm9k+P4+cZ2lJ9WbN+OQvC4hQw8y6HrzjrUnKt
vNTKEzNxzT92JGfi42Aq+XZNftt/aFkSJD1/DRnMXENjtWfae1PCjBMjdI2czbMB
ny3vXldfbY5i+iCnj7P3vMmxqRaaFW1HxPAunu4cWKOScekNgTr6ffoG2xNCAv1v
EQHItlGTFmOSMPdDOGoyBC+lTw8maVDb2iYFQxnx04FN6rEH6TtbQArlbrWMuasG
935uM+aBguzXkZShZaMz+0uWH/d/O/FDNYNvSeqgqVONMvZZuDCxO/Ib3gEtemXt
pOrYxFeeWwBi0tl4xplVWuoVxUAuBvlKGYOFPBHWp9xvER/dpQ9GQstc29yELhPb
VCzhVOc+nSkB0Ch6eZlXtqmsGnh8HRHP8kHeynNKIVYPb2mC5t9U/f/lxjBdYTat
wnYc1UaUWpClmWbOBI9pVBJWFA1CyEWKdg3XxiYPrpsdU9HxpPyc/N0YEk4Y2oSk
giaTchK6J6Wd7gcc8XvXtQ7TSTGV5ErSGoolcxpN2cQj6AFTniyT33tOZI4O8LGN
/rT22gvA5mo0uPvIFzMUAdU/8zMak3tBUBrUmIef6IPCwSUTldn000khtPVHVA+R
41Q/5+FtJxryKd3c4+Kj2rdT3DeWo0LBFh9vun/Cy8u0QPNZx+XrSiMC/VZn692Z
7AOODKe1N4zbD0/jR+cXSSPhz/aCuwblYjfKuNXRwOxwmautqVQqBVwqNsKXpyYO
M5JSGlaspXOG7z6gYXPoht6BCVFQ2YZ0mjpyb6w3VbbJecoV9kuPTCb7WMAxYJlz
qwih1AckvjN38t/RDsam0AFIpgdmfKeoGnl4w3yKfCrvp0bm/USTlkK8W4nTSW68
Ps38ZtNbBjx7Ch8pOWz1bn6hT5ktQlf1cnBOCyXHizOQrtdCJR0HYZvE49w1GeGv
KRd2mdZOKrRyP6GV/HYgByDLsq7RkFmq2QVUhgCy38INfRwQuJV5imK7lUwozILp
ITKxQzH06+/x7niSHzmrmX4BpkLzqxzdVLhx2TLh6qTlg/v7GORmfnFuTk0vjrC6
hP6LvjPFXqKBYurQvSR16xzXcDmOQ0Ej7V6Wr+21WlvxKXle3en5E65RdP4uQ9FM
`protect END_PROTECTED
