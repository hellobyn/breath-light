`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iyvm8WP3Fa6RbzQQAI2iA01tRTJKjarVh8tNrjf3DW5IYd5JXCi40y4AWo0jufA
OzXWejfYdBpfNt7W79HgJ2qH9RbbBKhxq8vqYvfuOLGrysr6Q6a2xKZm7CpFEhQ9
Y69JKooG4+O02Iy45tN9xFsCkGuE8fzkn2oyeLTJqs8URTQx1MbfKhukxLhg0wI2
E+fQ4bnnP1lizkd7UWR6eUdugksPQwg2VWijEJ3bA5DkwHkb7mAP9Hkbl4K5j5Gq
jkRGBnmpc/B7VwwMN8Obrdhjix3GwCRHOC2vfSWfgDuOZ1mhpFDZic8Qpl9ozh9x
nTO/IETItA6SiyoAxlGbL+qsOFFSnUQjFSEqxuWTMFye80kJsC7wdDBP/pL0Vn50
30H2Pa7x8+S4rP9BU8JKTAmvu42fGeuhXCUbvAuP/q7lf5JxdOMYqysQxr4wxMyH
Lqa3vlywp2uIWTRuHKePRZ+iSSFTQPJtd91rfj+RVuZgsEg9+MAFqzl0xtxRzjbl
kQ7vbc8ZEOxmlpzeyp0HzmHzeu0fxkZQBxVXDu0wQMOXDVBSVOYWgiUJvcxZ2fNl
d+anPkJEiHcvlGR+Hpv/qx9pn4quMTBPPiXoxf/KgiKLlJ3kfcH63R1VhPix72Zv
l8h1HC4b4+5Ja9XMjnE3mDeFMb1nv2C0lT1gO0CqhoEC5T/1oPJq8vO6sygiXHT9
cueonL85r7g/uwHSWNr1xwWqT8m0gVZbhGTRtg/Ze11flqKIYFJ0kz+832Spq28n
PH4kxBIiveHlxpgEPPpfKeYSciJmrplwGSrV4/jDQ6y2wqnBA6Os75PZeAmafjXs
KXIPkEQwCOwzGFkwK+S9syc4HGioA79+6VUC12JbjKbZoVOnYCMRpZPzSLVK1lCW
TX7D/5JzEok/5Zd1q0OeyghjwAxWNhOwgdje1LZwhR5zSXFHA6iWCobyn16nAhRk
sfChvVIWimeFqQqp9T6TdauclbenB7eNsYys4ZrU32WgDwtcFlL+A7rFiKvRKmqv
IPTMinA5SsaIhE0ED7bZb7xaPXEv98GJ9aHGvoUOBmkys3dsXDQ2SF3EiqGSz0+2
4I3pxe4OmUXyQoYxYnf3pE0V+R8kOpFIoIhaW75hb5CdAvAZb+ALKnZjRLDKD6eX
Rz3ZZVy1FvQwS/w3bpLi+XOoAel73RGMEqVLg/C7OLy2B6O3nXgrtiB6ueLttFXZ
HsmyPf1IsUTiiskuHiIf4vkspZOCyOrUI9i2jgJ3jewH6UeWdeq/slTjXkk5Fqet
n2zeMUHBxS6DEJy2+SclZBVEvSimjWD/qdBgi5BEa1akOF2ZVoFC+/4G1i9yJo9n
Er/kTsrnuI2kacXORvAd+2sdJeVnhUDNW6BFETagsyjO07rPU9z4A0erX1QStBzy
k6sK4s7JCbra+OIG1QlUM3KLdIGUHYUzBW4v2MP+JComol1MYJ6GAQXjdGV5iDa3
wIDOOVr5uPAr3mCigF07iFJYAOp4Nr02tu83z9HF1WgSAA2AgSTvEQyZbB0aivUh
YHW3PU9iCXhdGKkW4aptGtwVhAVT+SFsud6UU7vVeIoRDttE2Zz2T3KxDRB3Jzu1
fAEp3EGxZNVofVqfK3KKyIMkYney3Sbi6gGBs5t8X+gVQu6FjgM1fYUvgJfrskW2
U1MLdGmteXIBKtieklNeHoHh1Na41AFe0GLc4rC5XumvUoUMCzNOAjB/lk+LuPoR
E2HVvTnWIR9GYrdDNGE7vveBL+0JcSIq7UXu1phifdVjXw+UxtuJy1u+l1tkWSnH
HMhCvVH9xEg1pOD1o3D90/7T1eq10uuawAHN8T+qRvUnaqUE5YipBIaWTdRsN3Ij
nw0ejM45bThyeymkYJYtw5KOkL5nFc2UgDQLzrS8JtK58JTL5dUaOnjmtVoj4R3n
/wqih+s3cykyTEUIN2XFLxqx0k0d18q3xwgyvC5nITBC9fSE4/OWdhTddt63SKnB
ThiFIGnA+y6jyKonboAOxeB8amylEoK4PBJmQMtoq64SF/vQJF6YyBfhZ/EF1kaa
M0voA1v8ZOtlDkFMSOLv87HKcjLfEyZxQN7subbPI4sPZ1f0E6xgy6+u3OW1LQlZ
FRAFq3PizEOpSQGezvikV/e+oQG9rbLYj3F1PKl12X+MtLivXkqi4fcJ3wudkf/C
gtABk5ycyiHbgXgdTXiKvLVopVqXUslf0B8p30PR2oeYLvf0AwWQjk0kjWDMCuUq
vDSnY4F/HujRarMTxLG+Pvg+G25fkozHBFMY66cX5PCCSWdrl5PD/dmbb4c3Ej65
RBwb3JVUZWkkSUXJJAyXreAi8q12DubIofNu3lwt/AraZInFmGSDlmF3HopoxPO+
ttZIa0vH4KBVfjSNtFmojZ2ClPyQaRnxTfyGQrNXaj2kC5JoFGKCKJ03vE1oapPY
BDkhMHiEhyEiOd3SE1sZqW8DyPWOmSmn34bpuy0bWjUaduyeDxJSwzwS0m+uGD5U
hd0lwfdeNs1xygC+mgTnUj/hxK9+qMqvbq3e8Oc6nJg=
`protect END_PROTECTED
