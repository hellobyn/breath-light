`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weBsilIskeyp7f3wV49C0E7ZIcr2VY7yTglQuB7fjgdbkj+MpRIm9kQxT8Rkz5fD
ztfbEsRs9fNBgeck4HLpQyCXevLFLKz7OrgIeJp1+m+CbAoUKqK8zVtjgFXGAmdg
dkgNuS46qpclpWbnlSPpoCHpiK0eDXJiMgoLJud92vs2fAdXsEWU2CdX+cV/EmzO
b5tvfa9hfvXwr18sh+3wV9MxTSvPZqd0GxDtCxtl/f2g39yI+bdKaepkw8K0wJa7
kldqhyawaR7HKuqcHDmkbjEr/6YHRCLdAldsDF4IPw8BeI3gSPQKLZWXlybG204P
8HkB4+zdHOPoLQuDLdT6S2cRxCgZtUXHG4GRUVaZc1SywpC5ywYMTkiEFelwZzKo
E8BeEm4fqnEntcR7ELErIx9OLsvEPQWWBB5nKrenbXk/msLvpmtLNXnehUDWNNnW
/9oaLUo55WLtZNUGrtOO3+FydWhl4pxYZ1pB5md+WcVIhCbRI1H6TJqf+rduuDj5
VS6PfrgA8us0fuA/YW/dnvp0wzs0tWIifl6rNX0agFWSJRRQbsOvqqxHcVXMlJ4T
Hg0LmEN1tDHmf08UQ3DfiQ1BXeH8GGWsTT+J7A9/dI8s/R5mmjaczyYgTq7o08Ez
uQWF0aXBa9ikaQqdK0+znukzMF5SAiOTvr1r2QbvsT1T/IH801gYMHbSdMC9ycCx
Xzp74UOoeVpcvGJ9aZrEiLBfZzXURCikskI+MMMKCod9qEkVKMEOOvh0MdRIsD1k
KbhPY9Wz7nDRttvZXjoCkqC2M4gi48vDuj9eY6SHGfV21JXBReGPGbnFke+dSm6X
OoHplwGdQlEEOolbc9piomR/d9mfu6trG3nqoQHUEAlJ6uNFfiWS7jmZFvWI5+7I
eOHWGo1Pz62difu/BvzhftiDJKw+8RMxcgm6au7+irqc3rO1NbQYgjfUi3SDfMNo
R9rMtIM3ijsMHo9lXyZFmrIBxn74he22UjiVl0WyEdKKyrJjjJIgsCEwATXeC32i
GTLS4rphjbQ4AgC0UdWzwtu2w6Opfv7gjGvrVsteK5SfwCwWm/qZSFuHtyipPQVD
wYvAlJI83nb9T8OyFEpf3ShmiSX7o+um+w5RTEHQnuqbLu9NhpPdk6si+obtaY53
NUrjlLzRUq/7xCDEYpOFn7PR4BnU6hMy/gSGZfGMxG9AoKoW8rDgRTWvCcpSUIWV
8NGn4PZYeoR0jNee4OOtr0X2HGJPY5ducBpw3iTQxFi30nyOvC+al04lIFQG6aOK
517h1omEMSTYd37kN1/j3DBs20J9ZQz+36P6IkCEW/6uwzmejSqmvzt3bNlCTKCL
xQD6BlnS38SCb8dG+NZghxpu+mkdCv8bv6Di7knacCRAHQM/ChJfHbka7bZDCAKX
s3/knS4f82gMgCH4Cvau9q3JKhW0nQ6KRfeBoclUjps2eBzELvO/G8lsC2TuMlRf
jt98jvaPIFA6LsiMBx6O1aBwNw/oDcGX5SZLE9lrYBkBVwthYuyS5qaeUgPxrG1I
SJgQ9aPPQDrPw/jk0hPkMUUp109GKP1OY3aWlAX/IINbz20DE24XFsy5kJ9qotTe
c8Sq6zEy1JtswTc2Qj7NUNmrhdI/WqPyKjTqy+Wt5On8lzSVQsl4FUZngluWNLO4
J2xcn9cnPT9IO5mLznYr3EcqzdIzN4QMlSV/Kyu4JiqsDGSOc1xCQWYQEVlVaUeg
1GqE1bHZ1lBpOCqznPK2Bv5jYA2/mqbvbZ4LzQ0ywyY7Mu/9cU+FoJDhsxD5DpJY
phWu+bFRXi8ya9tMq0ar3Kuoyjb3RJNAGaVxu8TaNoTtjYwbwpjheuPKMMXjN/6f
fK7h49IRuKPjWn27RLsJRPwqcrEhwOuZy+THcbrhFiYwDkAq6JCcVjxbJuRidKAa
nPpYByBhDrbIwBEHwPE5FezAf3B3oKSVGuuVyIU+WxDvYjlH4ifeIJAGmVUWG2zY
uqooogMk4MitKE0hCVdElW881KJBYP7uMh+fP1Pdo02COQi+ws8uAYw95R/HWgCm
lVkWKZh802z/GFzmM5exDkyCRf1G0S1J4n8wjd9hJH/3hNPA6Sq4cGHttG347usX
lOQKNkc7NtQbLG/M3AmfT8UjGXtTbJHulvEVhmmOTZ6/Yda9i3kSZ7fQnsI0mokV
Zf7245ivvX1bixwNemOLOwmnoOzdshC5Whjd5+8+cX1pKnVOujeo3HFZMRIJATcU
BxFrRMDbperBTFHmcCZzKwTdWgJfkebtPc+0uHE1MTrgGa+1QuwF5W3NBQILLXyZ
iPUs8wFBgnKV/fD8SO3OZnBXZPgWIgW0I+Zgeq0iyRl5k1Sj1eQq1hONXSVjGgvn
pPe3mXUbYEjpjk3JdE0L8omP7y9ZLMUTLbrT7Xq1j5A6yBCdwM07C5HsoN7XMF2T
M+/WbOZ8tT09bxuBmemvzPw6odUqZ2hlA/+oHzCqEZP1mO3YDP8Q489dPrfk1HU3
M6zIyXSwF8ZIuTAp02lR2MBrhG4BQsWlUnb6bRB16k4RM33Z38qnZmID5EJCnOxU
d18aKbwHxgd/qtYDWujieL9Ozw+vll0G+Biomuyc3KmedR8PziTNko/3uG7zfbUD
P9FO52Qm5g7DsIEtpYR8WVpllZznXdWZ485b67IB2tzfH29ttB1qTFOPxiBXrOAC
u3eIpUrQ5lkvWsyn2mqQbEJaEhnPDnLGsYiVGNDbbL0eyhrnBWIJ9dvLN+k0bqNP
mMt9GeO/tHj1NyjCTQMnsZ17SAj16XgaUMpKpyeKLUfkvMCk4GGz5ICLXPiYfE+k
KKCR4yoTQ5ODArhpT0A5j3W50xW7un/2JFo2OMvu4ng7+LGqMVl+6neA1yJLGEU6
//mXIefOS5PlwVio0uMU//zdiA8lSmaHbIHhRRvGJcXd34bS5gMOdx9uaMFLFM/A
y/XQVAZR6aub1L7FTGlvj70PDVixQEzSsJF5pthqCSuLjcEuzatw7PY7nHhEk/Xc
P8yBBTvb3uEPFtnhnp6zmB8KqDJCo+3QQGzN/J9YDqq2CbqRdqnJsRDVat1rDJzN
EIQS7jITrjr1KNi73PmPbhR3+xOjx5HSWgT86bYFJIUArLvQkTOMn19ntRrQxk/y
JaqETMQcKRDN3q4CK1IGS7oSYOE0bkCTBa2Nw/HEge4qraJ48Rec3UAnjwgxSCTm
syEu8NsZg47UyafG/Bn7ndCACfmTbW1b6vZ7tJATl+EOrF2r8ePys6nAGiL3bnCG
AbVtWWNmgkfSuEAjTrB01mY1jftZwHtF65p4pj/VCFMIRRkTWQopDR2Of7aflgpx
BS2l6+/8lPtKfl3VNlOX42gAQ+phddk9g4za56Xs+uKkBbtIWcgxeglSIBXzFj+L
4XkkOKmEesOtVhAQsjAWX2inArlyruIfUjvP5evTOY49yjrpPIYZ/nZkHAQTQ4VC
puaicMgiKxBQpauqRNoPfKNBQYXrHdeU01gLLpXxRV77o9sxK91MnK21LRkqzcum
kg2/BGe4VbedbRAE1w7VyCcjbL1R1hZ1Ns2X5pfzomiVE+Ml+owBeFR1CBro7WaC
+N5RytonSFJFPe9lmta2fg7kxlRuLdB7oLWEN+wqwReYanCgkxGp9cPUswB+ALTf
Pw3yytaxt04SvsxcGGVHf0a3urKTtm+ognWq5GgC3vdVXZuJ9V+0QOsYjqN/cmZb
RloV24Nme3PXmGQIzOvxKwWKKD6UYEzYMMyXQTc50rEMSoAfcJPqk5ulKoitQXqO
2Jt1U5rC4XG6wZFZqJlvnnoyyJRhpFH7sCMfNnb/NhK2L3XLsIgSmEf50sEJMffa
OjAHJPrB/xnApKGxapFaBHLVyPjxksB7UwfGNqnhF5df3w+gGsPUzT4d/wDhDpni
JvsdWqgWoAoNSIUjFAwx2NGi3RndgV9jJ7UgTqpC554z3dYAOqVm17hVxGQljFh2
jJNV2+pOyUTt9FrQVl1FAuW21rMeftOh68tc6R5/5RDGt1fvsCn6u9oUL9NuRkKY
5NXfzvQnJzFN6upd1TaYqj2V3PosAJpHuk/lN1TTNT0Be2fq7emuJaDHuXlXlw+2
m+rA+6p0DJZMCxkwlhpwgiB+9/8YXAxS02ZqjuGO1+3UZcp/vt5cHvgs/3ASLxim
+6D2iEv0THhPOFCUo4Dp7tGLQU6WevmPINbyoTGn3qtCqVDBWPJlJJdZKGU7pZ7n
BATJP/f+5ojLoe7Ubp+cQV+qCiIyv5ba2ckilWZQajXb/Kkg565wreBL/NiFUBRL
`protect END_PROTECTED
