`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aV4rWsHX548H+CLms8ZeggWIank6xs7zu3QoH3/LSuVbXQF1zrVqLQX9BMbiE1nZ
C/98W2F8aJxVn4AktzdGdJXxKeCh3EfMMfe3FCxtQ1WGEVfgMBRBWjpDBvSaUlnC
2H8fegoAsrfJaq7nbEzpt8O5dYP+IB3z2Gac2sCq0sKUpeEJUR+Dw6i8YCsg124/
f3aoDtjaof4e/ljCfwWzZAHc2oZ/DwhOU/wruRzlW9c3p24Pj56LtQSdZ4qYW6Mv
TPPwiddbr6CTsxURWyLa/cC7SGFlSUrEhgfXZx1qcHaIlpVc5NdaAO4TCXjS8ibO
qNNJ+7yaJeX9LiOVzC7X3eQyEWwyNcVCZuILKdZr9/QTJwDzdGpnOBcI/x0WGWSQ
ojvquS5jtAjZ53VNUTKWrO0Y5tvuRYupH//TLwtaeQbbogiZo4ftKpIhl++pwsOe
d5FYpjEcyHYblZVc0YP9EPHlexIbvWqU+hv7POKNvcF7WDS8IbY7uPcc7KMBfcLL
+e+Wj3Zw71XFfx7SDSaYllYXtFXoeQZJLmWXNJfSlGHb+fMMRgmMTGKay32UdBew
laEEv6tIarAO/JRgVMipbStrzUse/12P2yhTzr8WuEB3JdcX7IhCyE14VoRBgd10
HQ2okXShWiBReUGeXiNj7wqEtjiT1y+Ob2mIevjSj+KFXvSiPS4+QJakZEEVxkph
GC2yMNdIczIO4Ls1jif7102Ec9d3bXn85mt5kCAg5sFOOdxSDcXrA1q7+SAyCDLP
nk73R+/uOAlP2CV+/Gh0dkOGo09KTS9d5cQONuSanfE=
`protect END_PROTECTED
