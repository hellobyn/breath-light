`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7sAOwnygxEcmAQu4mrCj1rsqN9F7+PC8gcvxjprdT9oIjRGjJFm2YUXzm1YE88U
vkY1TRWpETR/GYEpsGL8fkz2sDjH0T2ModjCmfzMKwGrgorvRCZsPXK9GZBaskFa
vK+OZYlJHhjjXW/eTkO1iiSNXHlILVLxgTKamezHcmZk8yJLLfrHOdXSFh/FZNnV
gmT/5YJNYwsn6LGt9AiSm4K253w9uTWml0tNXj95UoeFSZxg4Nh/MsafYrxiwf13
EdNx2ffqikZNaLJqbWNLNuktxsYpWtGefc42ltrhOXZ4arwkxToZ+Ei9E1TQcGy8
DkWQBel3TuyEWQjjARyDN7FG9tmJthD7Nq7roqNo3bbFQXopmuiR2YamUXVvzmGG
7Ml2IcsbOIv/R/XBTJeScrNKYMcBk6vuUKW7C1QHSHVJazIIVb/OZpIW5KZvdRe/
WYsEKA5lkvfjIg9smu2/hFcseq8E/Tqo+RobVxlGXYp+qT/AC7AcoCbtdNxBcSnX
`protect END_PROTECTED
