`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pWHgC/H/M9aqoXVKwDiPY6jGryFZPEjtnfkhBH33/RljJL8shF+8rKk6PpaTbe/
WBpK07VtRcEN0VieO6H92PuGIxhsFfiqXmYk42PgMDFs2QuSbXcdgwTJFvysBkgf
yIciwUzwrE1+vPrJ3a7CPcNXMwWLU7SZbCxCfHkITGtof5esvAz74TG5L1lJ07by
BiJkEyC29V2qUOUcEG+SxXhJqQe2e+LZcU5od4quxdCjCETmqc0zKy3MQS2U32Nd
CsvJMCuOYWvRY70uSZ5zapjPMDzWQk4n5lpJHsc7Jp5FJbKC+qiXRsAr3FVovgOL
JPbdN88NcdxrzylYlNQ/OWc0HDciuJGie4x6CgwF7TnfDPLmP0GQD12WALGO3aAw
vhe3LQvevELFcIkG8ux5fep8fupW5xwOg1UT3193bcLdWwvfcHIJe+VRZIkc3ef6
PPDsQuMcxsqHM6pApTRXthvLVv6/yWdjD886192t97G0/feWO3Cj6RhVXi+8sxn6
WoXoZYuonroh+VRBxxlGjbL2ZwRzZJyx9yTrJAtdqfKeV51/2AlPksrgiUrq6FQT
cmYykf4RFSYx0drNd3m2oyu6E4Bc8cxNw/PJ+bKQgNQW07xkTiNLM6vFUbnb6wfg
RSqPnfX5RJXEyJyONUwbTg==
`protect END_PROTECTED
