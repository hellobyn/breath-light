`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzSs8GiuH/ghbUROrunRSJpHoSaMLFZ+5r5sI6sunYSYs5hguwjT7OmNmPxWABhP
5IBK0I1kMQ1XBIn1JJiUPJGJ+15MR8nU4ouhfWImyk9Bp3Igz4G1BnZ6ORURZXPx
1pJ2h804OuX2IRnjS0MwwuNMEr+vfFyOdn3fQmWPpCx4O8s25CMHDcm3/866JtGY
NFcRzqQnM7G4o89ufmiMxM5u3POFeXd+zW/QKdR1tVtArFR33tWhDkP/5Uwfwt7l
4sVZiPhnpxG/UGUSBuJt8ARWalOE6rqwEaV0zwwz1xaiTqziURoHVPppESB74UOD
rrv+nesc672WKonjOezcCKWzdH7rSoaQznqGSz/FYQvZWfoAACZyMTrwWybEdIQd
3zhUpZcN9Jl+DmKDQPIFJ3VsmYkcHtholtvwRzaR3nf+Pxt8ZpM1p7BFpxSYow5g
Cpz9JSYYZqIcZaf3AIcpZfhZl4TLGodkKLagSSZMsr1kB+WnP7dg4HGPguBMlFo6
XZQVEo1t7v+MAU1vFJCjGulQun6rJvP1DivFqTwPFort7PggdwWoHVRFdHymA0Pn
hqoCzwskBRxevQk4pkz7FA==
`protect END_PROTECTED
