`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PsG2a6+bIbyPNDfGc3MIXaWq99qmHoPskOwlCKymv+7ZXJlcNuELlIAkxFF/zqdK
TScSvcQUYzmM7eIJaFV8KjpuY+LQdqNtMEeMz60COmnD6bkvxDDGSepY6oO4+PqP
ddAR05zI4W63fWAtsuyQxNOqptONq2cxAvGeLrAr1YaTwS2U2Xq+vrFPhsORQHdn
zkHbMuLsxjhm+xzaGpbi5FcrmD+8LGulyvXmypD/FX3vXLKmEZYDXZP4OTpyQW7X
hjwIM+Z4TWO2mfEPXhrxdU3M3joHq1rTUMKeAdekP4R7blF3yfK1KvKTbQFflGES
/MHI1yU8J3d0t8yfCkJqSDh7ED4FSWOJcJMIfhW6q60tqllyRDpsnBs/HPsVGGl1
tLx+jxjyNo3T7tyrl6OVpz72Xru0Dv/XChzTJgl75Buc544o7rLZUZw3tHRKspLz
kIBMLPlRyHMRe15PHvGrLACkXUJ4OnhTEInIqcSAjKPJHIhjp7zcAG5WtTzTPAEC
Am9wbSvaCWWLafMiz/NQ1w==
`protect END_PROTECTED
