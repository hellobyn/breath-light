`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkjA9qY6E6klWX1CC0TermX9WU+lN+MmB9CXwPM51qGMaeJwazK+v84P3oNIAOK5
Ox8+3x9T3g5wLB7OV25KENV13Bqvyz3RGnYdc+utab81kjTndtZ6X9EJappq/Gmk
VvtYxCbbreErgFsytsvLNK6nT0RMR6iCVzr4TejixDI7wo5yKu54hjFqqwfWsmPh
Rew7VB9nlp2UVw/M3093etaieFsJwApY6yeea5tZticaN1O9fDEV/Nqdx/OVKYJB
a9fiLVrYYt//TU+FE58TBNTuq89BlyxKkzG1YNru8nmGNImQDnwuwtpajAnsKXG3
7jKQXCBqE39ZSAkXu7Pq5bKScwAEqjE/inlpN1lx6nGZBf2iaLrShhbKxYmT8kvP
276KrWYe9OllhUenpmFG03B42QcqNV5BIEwDrDQmjGpYhYj4D0ocRew7XHGKok53
nTiYCmtSJFFokjPGoNVl26TcXFDIF10IiQvVLxOGz0LR3UYXGuJ9n4NxP21UrTa8
ZQcyGTt5LVQSiJ9x89iG+v/BY/AhsArBmDkkqevYrnlraEqUAlPs++/RW5WIppT7
++HPqaeDpI4zuRLgziHv5/orTD1EhI92vDvtAB3Kh3aorodyLzKMOmPYyIC5NDuS
8EtmYxeroL6hUF+U6lxnXjkdJplXCSTPWhXKgVxSaDJyFWUHtW11Y3JWCCObE8n7
oD7cOapW83Ctk/0WHI/rFq+2tfAMnHLiMZ2Fx4w61j/iXcTQ17pBg3xtSMNamk9V
ov1IE9xavvrooxBapmzsgtg/KRQTRlX/US6Z6plPC5BoQJp97ddZmjaS/apwPH/Y
zRT5+V347RV+1/UkL7pFVUu8iVXoN8g+xW64syZYB0B0QrvD4TimC+iMWXAANu6E
ZUmV6qyMrz9+v3kRmFQJUXUhBVyLjJEA4J77g3b6RgszgwiQsEN9tkX4Yu7QZVXP
ZgYa4iS1bpWeKiBaQsjQbz9AdshDweVWRT+jrEHLvahlw8f7BEsTbwRnvYAa/gg0
Lde+lbtNCOG+MG4tatOTD4NPo+6/CCB7DPyaXMe657FxWC+zvzHBlQBvZK1gXJcl
98Hnesbjia5K9k9X/eWe2y8byb1shCSqTQk4lbuWPZwlX5f+YGXl5kRVsTLHEmgt
VUiOEIDvdEs075yyKFJi56GEEpv5VJEO7I6UWvr61UUx0CioYOnwUpRK4SvnD2b8
uDohiyPRI9Xi1waIJHcIcIhCCM08/Y5gTkZ4kEbYapWStyhDjZtHDrq0l0JIHdw7
KYZUTlhocsvuxT+tu4kpDhpqXTdLOvvfWaVKRXkO3/VkUwt+H1socDDdXER01Hms
z6iStgYhfGS4AvhCunX3tfSSlq9mYPe1lwdPCFdtgOgeaH4HZFR0FdjmYaoZ9gwd
qfqRw9b6ktTK6bRll/a/K2ButfTlDhbMswDo4MSHvYHCzRkuJgr7lQfXLUW638io
P7cI6WmE8kMJ9DRZxNJMNxnu7nKbbKub4s+EbTcnSAMsOfVg4yYrW/f5xjqpu9xX
Ys3R6Se57I6e3Sf3cD6O7J/8Ol6eYg3lGT9dUm1WSNeZXsGuxu9pp0OcIzLEWm0j
1haj5ia/a1oAYZLn34vFz8O4XlOpevGDiCP2BJRHY7plxseCI5f61e8IvWK4bAcx
/y0NGK2r+qil42hC187DNDJwhOI+DKRp8+PQBx2aQGWZ6YTVe9ajqedthvqKeg7Z
FbytByFlmIQNwRWQBWjjK9V6Ry/WPdFi12/krKaIdYuxDgp+rpsf1dAMdeyIa9x6
Xf8Gvl8YQ90HLKRMrj5/UKyWJOaIOALM7BnJ3FndvBxcMqX9asrXYQuSLnu6I7d8
Qj4mGK6IfY78CLfj6KNgfzKWd73q+5TOdH89G3iY7pgdjHC5QC3QQWE4/ZN0M/k9
Udqv989Iis+gLByrd/FtWRy6Ioj8a6oFDq22Pq3evyovrX+9S7R6VmMDHTiulQ/X
ylQnJZskFAMOgzM1fzsPxtflQg/YLCbOR7Vuzkzb4tsKRasicfBgKe/Z4tD0/kok
pvQojhGOs6lreenSMVVUHRkn6SSRKQ+rWb3QX/ys3C5H/6BhBqtO8NouauPzo1kn
k+faSX2R1xzxMO847EQXmohwfush3UfQqE4brkqqevReWWc0FR0Qyz31Ob4IUaHB
cJkFvHG7+DPc1SWvXGCnbNjwQa4R1BWHVXHTefxgjmvKiYNS81b9GqeCXKvZbcbQ
B+k1TPlWFJ7hkkPH09N2/TRYal1q0yQxFHr4iRWSL2oB+PS39jfSYih+0WTweGtu
yoRus2PxD4Qbc7OeMYnlC80mhyw34UusFQGwX3pzPdAOm2wQc4sVbUK8IYX/KfRT
kyH6W6LNii5NpUD1VjmHa5eU6KXncysUavVkvWSwkz+xLW3FCeO6AlXRQEa4/oot
3pHcb3tvw3o73dr+R2h2iGb8okRZFiGLARe5B4Mt2YU6AJ81lqn8OGnK6XRMpgux
E04E1SMFdKTbrnrclTlJMOfiHfFq1/9JeAqD9llV7kSK9TIvODIrQlh74reOYn1M
Nd/5pGZM0fWWezfnTXVD3c1XpM7s30MrLNRwU0zgZ6utsV9eB+FBexIhmrxCR4VQ
98OF6dWEjTyRrsZ23dc6rC9j+mel94wp7iVTCtyT7Xj4rBFtWqTQp6YhRrnpNlsH
LEi+E/lUMLQJcSe5BWUcc+HmljtkDNSrlKBcuKi7foFRs+/pckPcWAja17irJ3qJ
u2dlOgmciqmbd48KSPysUHU5M44wNRAHc/FzU/GJXkMNWEHYpZjIDg0BSHbTliuA
C1szJnzyCOdJ7V4qgAMsWGov8h13wOmYEoX3B2f56l/mBI+DvBwZwWa9uX6YeEoF
Uk3MK62fT8nxs/WQ2A0n1yPUNM1YH+bDdW4KvTxRjbBbd7G3na9klnmIhrfBdXg2
kUxsD9oPSZjv2DtS7r7s+XJU1tvm5ZLCkughtvovHBELTE4TxRw+2yNtSUp5y4W7
6hbhc7nAULLty8wde+yh8OOZmvxEhU6yXxDri0Y7MhDUjTwvzJ3sxMBs5+KObagi
94RvP5d1lnnePdF+A/ZHJk9HsiKhg5B0G44EnIsZXkYJXtuFG5FeEYJL222h+7BP
J+7tVHKqRgfPU8XrgTcuYGlBlHkVkRejXbIYAwheQYwTHJbOFh1aMFgyjihCCiNn
05z2R7/5y3DS+RaIPwh9Vyi2T3XBFQuhKSvvqva0HmdBTdXslrqRAKaKNuZKtczc
iBGTT38OkELlESlzHpM19kxvPZmZxuHh58lQAjGjsrUPy+ahotiPmbMH1l/QNzP3
AyLpNUY02C1XsnijsIjt78dqQysuPYmlMsaC7V+N/naOVLcTkphoxiqxvJACq1l2
VA5TcT58jPyAjgJJmp1/SUUxDmR0FlOxwhtFO+33tnbOutpnEQenQn1hzC5j44i+
wOixWh51JP58ICqCzMWldV8VX/iyZSq5G9AvJxi+wG8vvXL5QbSSnkPBCHFmCQ1M
VZpYl6cFeeaBt57syrfJ5KyreChx9FIJMfp8bZ/2gnIWiSAraoQVBfycG75BUu0x
/5scUtYY7SUC+P7h+cSRCoOHW7bWLAkGnDqcijg5kN4Mx6eXfRQalBp+G2wfK9ab
4+BeZFMZjKZfRN5wJFLwanlnZhkYg5NLjjaUAQJ4Qp2x7ubRe0eKuFLBR4PovZIv
r7Uprcux/IU6T2PkIGBcDdNNK/VkYQ+YqTRapA/ALFED6QUVXBOB1BleUBsKYd8A
mKPWjwnDRPoWBrZdXMfMe+CE2JTAHh/u6iAtNKWMWSKrCMREpeDnsSOiFVXlU2I0
hOAzHjJp0iS9XrMZ5mXgca0upYxSvmz6vI6SKtT52ZHju6c0GLStx7S9WrtmHg0w
Urf8UM1LQ+y+3QR956ssiDFp3P90/8yzLeKUSIun8UgwukBAKgeZyCkGq4OJVXlU
A9JNBAY9iOfQo2tdD/Yb06VeC3GCqBn+IL5NIC0hk/7FxWpEZVONtagw4Yjpdpwr
0t07jEzEX6dE7Yqj0mpEJ3xpygFVfpAE4J7GNe2uuCUSVNnH5qnU+4zyTeczJ/tP
rGcUorl0Nlley4GfJk+8bIV2NMSfnad2XVnEiV9ATdz7De5cZOZA3iKLanYgj6A5
ErrfLmUA/r08By6bRAN4l4OinMa79iw1vWPxfW41u82xVPhFTkk3UljlB8remuW0
IG9bTbyQGYT+wId5WU21G6RtEXtq913l0avLH/igj6uT0D7VJiCFK6MtK1oZ7YMt
V9U+ytUQO/78MOheyUMkmbstqrCi6U5AJnM/ZOHSFN87KFLqeOp03a7mG1IndZZ/
KxvdUSnf5nHKzhtVgjNZm+xRWMRz1lwg1WVbWKCRcQyxbJjCw54ZNaFiAwg1UgUq
0sa9CuPeJ5z2yTuwqhM6oKJgjQvk/GdFM+1D9ZaAMQq0Hk5df2SNpG9K/092s78J
cV6B1y718v2DbuaJMiw8X+hfgMGnTzZqAB2Q9LTbe4BhHnTOADLNT4WPvw2/kO4c
akSufOX2KJXCUpfkRh/FXbXY0HHHunzmNmIALTjlHEyWfYPXxgrgUSpjdsjQlQeo
5x2Iy7HUP5C/FNEaM0LPUnjZrOEL/22MR0dhdnrB55IpwENXth9LxH46Cu5kaAG1
6r4KA3X4D5nqOaBpwfeUXI7RepXXSXn+1ubi0aaLbaEehyhwzmC512Exd/13j4Nq
eWVOPe/asIB1aOtHrcCEAy1yI300hPhOHKOSD1BCzEPnZn99S7FpK2B+3dLx9Iy9
C1/DtRKqFPnL/I58VTzpUhn9aBTX0vXUOCsnT0aLo/mHrRN7Ea1+GKI4bK0N0ari
RvOvl26ph4p4xruOtZun1UF5rQ2mr6N21n7k7FLDBmb3xR3qymdBi1SzIecoEbRt
`protect END_PROTECTED
