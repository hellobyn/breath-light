`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILeAtbYWn0wpdtqVUxnSmWqAc6l5Vjry1wRusN3zzSVbDrdn1+CL+Bssjj5pDhbf
VsfMI4Pyp/XtlvFPCksec6GI2RPv/QXbOBQLsyEwQeSoI/Ldv2GRIwInYrziO87M
WqlOzEJsyEifQgwoe54OFceW+hrEJnIF3nKH9wNRuX8ZuUcb1R1lzJUg9y4SlVqr
q2xuWZ/hqCdoE0J4axpnnAolTWcJNDV9ZVOtiFCWutOZJ7ww6BqcqNE2w2RHKxFh
X/OJids0/H4cUyCKLJiDYXIJjCGaPRjfN6eSYm52xW/A8Z5k/AMaVtQ5IuC1cujv
In4O+hITnnf1bcfP26BCrDnmvgMtcUa58Gtdt+SCcc0lsrb7QsVm8MbSy9PBeI5G
a8b7gzKcSku3OWzuQp2nnGzwdY9vvYHKTT5AkpLRqZFdTktqbyIXChfPAJo0NLMt
PPYGyJ8h3wZNmnuCXaJTjvKI6ESApIBvmEaWGLjzc/bW70hBvOJ6K8gcyq8o+53e
5WH7fut/6FHmGWewStJ4QZMUiBHupqWFYbd75eHpOi+MsM6FhgBYRvcomqUvnWoH
JLmxwnfhASNk/1rmLcehX0CF3HoT3l9wK5CV5dg0ecMtTtJHN0sAuQRj/TRUKa7W
wHFefMZYAStquWn07rHEPtPwYbWKjZkpmDrUd1b9SCVNSLkMj3wg/LN5zy1VTmDK
7E4gh6aMD538fWeLvv7wtTiC3EbIcbA0VYbsStcZn7TRRt/QisFsUUgU5eiBZuJ2
X2zuwD6z+NYauQplRGEebPiMfsQxH2Ub1z9yZNJI4TGdTBx1TAGYMkbOey7uSBit
eZ5o1AFnyZP/k92pGwAkYwbUOlnEW755G2iIEV3x8nSxn1tzYeC0xFK+Kokig2Py
cCO8BybJQSZzKgA3TaAWg+GKhrXrGq72kSAa7l0ZsJNVdaj6OO5IS/l5oAlSLqm7
aBPYdNKsqXzldATqn/6nqXr4pvoZff6hy1l+ifbfMCnOkuDP99yJwPd14ZweG5T3
s7cWechMsw3khumJ8U90Y30P6Jz6+yV+WB2h53bQNP0VsiFmGJToYrHIy77Qm2eS
ysT9BmgVt7UGWxltC9is9IbhTe5iGB9re/D2h0MKHD97dGEuKmL3O3g+QuSKV+rW
YElgzNcrMlIgxaYBXg8vRdkd47QAyr5QMpyB8r4SsMw4KbH9iQOJDefPzjIHnG+w
u5bAz+AOx+1HLYHgJYjQEULwvfD1Dhoh8i7gwkG0KkER5xKywMRYPiLetaWe07IE
D+bS4G/Jf+MHODQmtxonO85V6BMCHQBuyFyGUewSn8yRYqLqIcg4xweqGWYlYBrs
znyfUeEBzZRa4az92Zm//KE4mtBIcTYxk5UebJ1vRmvg9BItHIMPqjaIM8m1brqN
Qcvp/KsTUX14NJ7eP/OsQFZX4M7gk9OILFAaqhputwveIq7Oz/+ZPicbTZUF/k8H
zQED7jI3grTSAPf1MdHsYojNdGtjgY4k+ZZopzXSUf1XrctuDooMVfNBHoM7/1BG
e6NBpViIBOOvzkc7xxvGCk4a1EMa1cM1KyWmDy3s+mP325dkwAl9jIE7wJK0nnWy
Pgykr0G2iFJI4F+ShH4ss+FFTW0o692vCsKhwqv0lnq0kWUkxu84YFjbhjJsx4Vp
xyEfi/85q65/OxfSm3V4MrnnIxYIHuTqlMZBeM9nkh/RVmzY4DEpDXNya/cU6qnu
WNOW/N0e3VLPujIY3wAjq/MzhsZeKKzL+fw+L+OgfJtohggkfGuHy+Xpq9A4Y94/
PTRQRT6GCjesRRfMDlJB8NxVNni0+uQMwYUwR3rQMm6Ada9yz7YP797AR+dgZ8PT
ktnb6m5kElXB1zVDHE4d5aTl7IEqme+xGZMLQkjg8B3G5QPTdVYF/8f0i6TG+EAa
90/zHgzf+BMnYopX2Ik7Pyo5xw7UT62neRHAH/3D7C45MMsto0nMVL7hhfnfGTM6
igB+ZMC87MD/5DhP+3GXBKcIRP6D3I49/S8nwpI4E+LuoeZcocS2njXgakWzv6Fv
6JmdxQ4lOBUwMfeyeNhs2WFRjAxpl7R9rmGBFaIqsxnA1FmQR6kBBlJcOVh6amXB
4jJ6DOs79hOb9lucpY2blDyS8koO3sEySB3JJBZOCu04/UKGzYgRciTIfXQy/695
HA0EBTxjbAKJzjaJx1Q82iy+0EltgjDq2sTqUoJWe70UVmAx9lWtZsyL0/9nuOPt
zMP1TaIElLSi+f8R2yvnaqyjQzARANf6yuT0vmc5BxtJ9G2einY9i0qpmy5HNOQU
I/zGazF1peu52p7YJBAM5S/WHgZte4GzvgCjB6ZCV1plkPs17LBSK0d6VXgQHj5N
G5uU3hlGLpFx7kFBwOalVlrBhudqBhE1TtKmOQeYFT6S5ziaAHueQ5gTIwufQiZa
E+Lkq+1nAmJtsEw4OyyOoKFPRQClA80Gtmp/toga87jvhKzXSTUEcuHGn3GE7si1
gjnd13MOEow+U0TrDemzwV0sIxYIj0HIgGJCJVEx9dBzFuzIZe1C3zQHpUZrW+px
w1kBwS7gtfw+kTaWdirljKff0TRo6lLdLJ53+ChKj6yVlltvwoGyeIf6qwtXHGGA
KQj6X3b55vPJKzmN6BBWlSKCcyBOQGMTeqbWSsjOeElPweGh6EoYsxAmlXmg1jzL
wNUWN+oWDJFu8TAjaFN+Y2VjeTUVti4jxiIBA46act+gVxF82ApOJ7eKnLrdGPPl
Qjc/CV52318YWEOwQpyxSvUYFJLE8zeI2wQGU7vj06Pe11o5q1BOTYzXRU8xs8mu
rkeWhGPEHJB6fjrPCDY5ibccHlzeHhajAIXKraBsXRrIqvXjW+hoiHNT4G+8Vo36
8xso3sitOy97oU9VAX8RlVdsS3zx60nIOUQ+T56odkOwFHbwruR1eTNvs2hjdbFL
qxbSu0vEp1iqA9/J564UsjKW8r/0ZEr6RcMH1jjzUZ+BBWATkekrNqPRBhcbZCr/
Zs0q+0HlhmhMSI05h193GPGtL3hEITtg50PtPZDZuf00vXcisIFZSmeifmSF/8k0
EpnwwVEjUXbAMTUwVBYJoinFkVIt/NdARqhrPDqHhiYs2Mj89w3g9Mdqr8L0KvKO
Sg3U0HBJ/XSJlOQWcrk6UEN6PvQOXfe5dwy0VY3xQlPChrq/k54ZuE4+SyaTnkgb
/0vIzqNHDafRGdLEJ9A22bW3UBEtXKfnzS30bLhBZfGvrVrBIey7q9GG6osxmAKC
EL4meveG8uDL0Y7FNhPnn0e03hOAQS32qdaJUYzrYIwDn6Q7mDO0iWBU57OHGTCj
VOAWfU7ULPuEzL/uyFz2Wx2wBHeIkFYV7AUKF+u4iSKBQgH48m5929WgeoRKzFaA
IAChrUgc77C77fFy7VQA68y8hLX2RwW43Z/hrdNY71sZZQwRD66WVw2I28di/aIq
MIbuE6wE2nC+ceOXV3UU1fP7OONDijdKTp4lrelsIuGqf1Uy3xrIJamHSI+taU32
tKM7wKM+6r1kobtZefpGWoO+hCjg5eL5FpeCohzxKWRuCcfW2vJ9t7sfJqWzdH1O
ZVUPY0ApdjvZZsqgO85q6MlZaMRvu/qHNBxnyw1ncR+Q9JRWOork3Te7Dghr0FPB
9yBZvrNbt28eiL0D2gD97tIrxWkAsRZSd9aSO6HWDV7kkmXzZsj3SScN/BtWaonW
QgWcX15L8aAgZwkoRagZC5oMfBam2B/G7nD1nyGryhupsNFHWmpF1Y8zDqpDcLha
/Mfr+TDPd6hySKvX342J17NSX9ApK3f/MYIsyY8CB65MTksG/mqYJNYEtpwE3G4u
o3S8hrxurBTLQgYReCA1lc9gv5n3H6dysNNUjD62ROoxvVRknEKJIBs5++mYES2G
X/+TSe6OpVBO82BDcUcyvNrY0cxEfxro7yOkVHZu5a7iW8t/Qmk6knL9MgxyRU6K
Gy5ezXOrjCG2LN2gBahQcfVpgKbPJA1Vb6GYWU5FhrSG1/wyO9Olq3RMnQ054m0D
lME1sgXiKKrdTygAiQnDbHPPS+ly5FBZ4WCesPVgd3MTaHx/6Oxv8twTY1huQXdT
oeRSk8lj4jH+YLbVgyezS0x80GlpTRU1fepufxJGpYaov7qFBn3T7ojtW6dAO7kb
HKCUwhi79qjWr5Ik3yjVtQ/Di1/8nSvAKN75dIlwI6aBdCEcuFqkk0P85slCIgrZ
uahaTHFGVFFX7IcPB+kR+0vnoaIvUE1Ko5YyD2tFFB7OfTrXIq62v/S7J3TnUN0K
HitNZGIwGye9ztbuPQIyCi9ME3vrkvK3SEDj3QB9WYfO4ot83ef4GyRQtznsEzaK
A5XQIqxdf8RUeXwY7dYG6A11fJEtT7oRdNKsYh2+GpfwbKAYMWMhsGaZMfEf1JnN
Spne7LImxGFeQ2VPo+mjHVr11mMY2QKDiwIc+toCns1/Ubh7EwbWgzkkYkRTVKmC
KOyMrlegC2DIpbPNEQxa7BqtN4Njvcztqhsv3SzuAVS9Bu+JLd8voAVqdRMVayx+
yDK9w+zlrx6Liq16JdeA5gWr5EAnLftgZ/UhzByTIe89c6S+agN0R6FKo9CWc6DZ
oSnwh9tG6+8V6qb2iVMOYHfahacrtVyp7YBJiBZ+ZY6w97ZRUmPYWzUArLphEezX
R0AEipYqkdFIFXnB6TQhuEScNCd10RB6EevgQuyB7sfz0zSBDdOpmFoMc1fLm6lH
d4NRGorrVlWn+pUPKMC1aNEaD4y2/raviZ14pSZpRIjfXuHQVfKDezb6Gr6bG+aM
GmqxknzOvrE1ZbjE3vquN8sBfXzsUZVtCC2FYTePxTOMhm/G8LP4mA+p3WVDWtNm
GZcdAUPIbWpmhYs2VC8iyMYP+ddoC7mamZUhKgJ8qZ72H/Buc1ADMzPIFwI3tCNQ
dSJWN41GTmz2i1xhA6LJr8gzVHvGRrocVz3WCwDldLxFKsikaSLGbAbRLyXZL5+O
j2sP+j6SdHyTD4hkyE570fICUTpLoo8GuoW+y/celVu4HBHYtkEJoYQhNQ0r33yx
vjOJ7ovx/lSGBbiZhjPOxCYbjtijCPTxbdz0SonawocW18p0MBdK32Ar4r2lbuyr
IXlj4y+WDGz0qw3fSl9CIVl1Qu//00/nviXrq24ue5QAskF8LF8uuBCNT4AGigWw
WpOH/KTYGROmVBFf7Ie4UND5P8gH8SmCgMVGoTljU5Kj2T8PKxDtgWwsj9ezD1I0
5eGyuOzx7id7fvX/pAJM8hD0aWCJhqu7+z1ZBRJqrVqpwXumDijTKYzl+Ngxp1Nn
IPOJTgaPUaBHeAOnkcdr7Q0lkNw9lBB9ggEFG2kN2JQVGJ0b7FyOc8aFgn07u5ST
ZDIA8ohxzGzdnJB0Mq2aqp6SwKXuDkII7bUCZwI4JqGjq1UMuQEcjKQCRTAXwqbr
4LvFfyt3VjkOWqQysOyE0sbkTiPJAQR/2Ep1Z1O7SmbXQakt8qhiWJ/30PQSKrT3
51mLIbm0dXBVLnddtYzmfbpY/Mx54hdZEXvTX4mGb9GgrRbcneTpmfnQCpeF7b5M
TwLLHNO/5eLMLxqHJMNO31PIGwwJeskGrqG7Jv/Ie40Nb7K/vGcLE9auhJNqJsi7
qcM4X2t6WtOpt/H0VD8z92/yAdH3IQbo/kk9M6b8kISXUYsqrE/6+ufwo53nBBfR
mov91yhAIwTQTaj7pN5GoBr0VART9ADUH/KFWVPshmrBCybRuHpsJwhUG8lqtYmo
twOaXE7CfyZhUdami9n97paUKr6VHvY5BHZSBwDW7j77SyK/jZ8+UUpSjrsbHmVc
3acBxjLDxcRycJiyHbGQVxUSquGrdfHIrPn137tRy927zh75Lj0yqLNxSylcI6DH
hnEvzA9h1UMCkZOstZYlI62RNipY+U30cdvA2hTB/ShQYwaB32X8fSRRf9eXfp7l
eCce6xIco/K/xTNVC1JOQK+JlA5uoO4BzmFwD/8P7BpfcApd3EjYpZgZEOaZY/yc
tvMc1vEYmwYUchsBL21hfMog3CX5TeJdo464ovFQEcBEuJ4Dthf0PHJPW+K83Q/k
WcVSCbZT9RQ3Dp1NqiC00bR1cFDgPgZOlr2hz5ERXs37jfIqlaWe8sWtRq30u8+D
KFUJ2RW4XSJLmQAg81NE90LyfwbM5+9YOKFA9z+4pCVBJZfXuMXLXnd9bx0sV37d
mXuaEAzoZgeJpG7EElHvNXukFG/14wOIfugQ6/O99w521jNVPXAKZ08Ir7FxRE5Z
39TIsBuuSnlfhLPibbw18cHO1eSfUusBW8R5oC2j1PJcCZQqmkYZCvKzMPCyx5kk
HEisfJbeKWcaZrspKIi+Rhhrmihp2cbQ/AKid40tlJ4wudQ605w7VsvalzqcOzOF
NopfLkcWsgDLYtU3bxI0rHyD1U9grNjEYZVmMiA9t037jWM/9m0Kdxy7R65oXVXu
xYX+kAG8lDYufQroODK+OMoew/UM4nZzwu+Zy0sf0S4nrsmSjmTBKgNv6eG1H2Mg
CpBrQJPG3DPwZCafEu5L2Yxr5at7JLm6WukhgjD/qQR5qsHRZrDHJgDwkLFfDoyb
/AHD3SL6DIw2NXkRdfvdwuRNpCLJ5FMHy8Z8p+YEorKI0uOKcOtKdGEqimjSpejY
iqBta7K0KOQWWi2UA2wK6b/qx7mqRSVDUU0fIv2DTmmxf0O4bWJANsQ/jG7R+k2/
ESsEvRZ81emwSmZfvsJCUQPvO2kcEWQoRn/cVMgvDYyyeUcF5iue90FOFnCIzwkr
Noha00DEwvFAo2bUc0D2kRHGEB30w7Op3aVsMk5MIFlu9RMWNMpJeoo2BiO8YrUr
DbH8Mr0RpN0qKBSM7H7UTOGCOOil2ZRtMo6nFLcmldx5U575np3QjBDiz1WH8ImL
NMUToWjxw0XFRNYtCO8wZ+dv8PjOuxjvgM40wjHsvKWQuy2isJe+F6sHc/dby+2w
6jyVVPSQBjhqiwVauGpRAjV2E3scjHlA+TTvQfveN4nyPh2jqmtDKvxeLCtIPeuq
xwJV4r5/UuAf6stobGhKHCfX3H6x9tFG9ARdJ8Cu6x5Lpks5sbkEhiY+lndWmXjs
4sdxPA+nq7ctm+gJA6rNxkiIDrSGUpsDiYYBraIwe+GoamVMCXp4n8DR+fexUqRG
YFJXyogJ0GrxD5v+TrB6Ds8ePqFeK6i/tCP/Yy9Kj6N84QK7Qtt7IdeFzYyBTEJR
yqPT0HSt/jHR3pRGNv2vxo6MGD5HOR8iCfD/EvtMXuPJYp/cxfGAnaufZQaNuBrK
Enz+I1lozKvVcKQVfH59O5T8Ry34SA+3+BNq1GfG4uRxqSs+FPlnYwnHnwGSMyDl
sVOpcjIRt3Yhw65o7Sv7u5LnzWrV0hiexImr2vm+c/T0gvvkcwOYxL84pfrLYmbx
PDWNOpUAoeLk5G9po/7QpKeNKu/p6XSkRZkH38+nZwLz0B09gN/MhFk+wuluOPOg
Emx4C7i2IG7rhZ8hhPnCrCiICgBELP9D+akXb5wBk97PYJDTOgBFIG9bRh9xS+6W
6lE/Q0c/QhvOwl373fRCHSsaFMuuVMNg7/K0Ra7cCqT2qR921dx32KDMFvEsvagr
ezBYIKGBK1iRabjCGktymh4LgGlWno/EHgu7VybjCirG4N+SLWjHk++eoeIvApEJ
ifqE6RItFJeHQpWkbICZ8ndsGsmj1tkT11ZbxGk7NVksHIlrplF4geRGjZUquJab
s5cz2Olr7ZtQHJPIAYa7L4BxelwNWXE7hoibVcjJl3RfHCN6rrRh25lilEn3ZUak
PDodSZ4Kzvi1qhpA98ASierB4JoW6HLyTwnau39MFEIT8LA7xBC7qBVlZuvuxxEP
CJVrdMLA20zecJD06yOyvg5UDufmtNXqJ82/BEXNLw74ciQdq0WIAizeRg6O5P+y
wtDBZC9r8WuiA0vKF8GoWp7z/JUz6FOjpecCdSQtmfEKRqCM2NVuLN/oCzxv8rpr
tk4JA9HIUiQU255DFv8W17WpS4TRTOSqTlIj0io6Yf5n/rn0SHJ86eXWt6XOT2z4
XqB34ExoChneoXYgnmKmMhIshOTyyvyfcJwCvF85deKHEjas2oOve088hbgVX1gI
0nW8SjvapWHSUUvJU8tyj9GRWi15w2A+JHILLZS1Gb9d5lNOMU6kdIdxDeft3Hxl
+yezFKd4+umvpav9FpngkQ0X6E1Bni+PfjxFBWNNZ1NYd0YRXDTQZ2gxi9KyeI2h
/824BMxX5sUrZOtiWabBJgmQYui60j6HlAuHvpIjlWKxXKLQYgjiaw5p2yjkPbzI
WpI9ZEsxGa/laKaoAydN9IikWJpPN7rVHtu01OCPe075PDqrN2Ur7z844kq2YaXy
DvGJU3IAuem+KhToktsWbTK/Hcu/zjssCWG7gEkYs8zAhxMWV0ZV2ChWztrUfKah
PmyxRxpxhVJTyqr1/qzCLcS1MI5T8jjmXNUxP2Hy040R1wocT4zyXkybYIUtAwkg
uEIeNQvNA8voPu1WNuKy95IJIV3KL7l6AQUXHWbMLz6VlXM3iFLawwXWQjJHlZwe
SB1ndLWrlV71bIV7MYnf/YbvimwzglqH5V49hA9NjE4YP7yBPWZZMDBfLFCEcF6n
ykE6EU7iykExNcHb+qItEk7arx3e4iDJnLokUtu5FzBZxAUmDDDqFF8v3dpMGBnH
3rxdjrMXAI1jFiiRDSlh19aDHlmj9dbCA2vBsr/xNkmowjoNfeGBG6FfEYrfpOQI
jmwGUTqUn92AbQKXRhPIc94Qs7/SNwCEAGGCEsz4gujd4gAdP2rAiIEn9oxsKCra
LfDNVgJOiI9Wu7FHg5Yqu0H8LTSTl00w3lfIDPjzMvVboA5MmdiVLO4gpdZTez5O
oSPsPLILZdbKRpP6Qxp+9nxNXQ7I7Ekh+P3fTtkx19RUYgridyg57Kwe3UGPD9Jj
7pRJqijRgJ1aJhWR7xVf0jJ5XK0aLw6DKIZ30v/YCzDSkbATpp/IJq2zySTkxAD8
1oRsd3NLGWt1qFhaP40J2kI1ET5tYec4GTFB6mtOpk0D59JzVb7S5zNZlBZtWw+S
fjfU1kTZdBrJD3nUjZF31sjAK4Zjdo3wss1QKj/GTWuqNPOnCPeBzJ84fCm2VAWr
YDh72JtNWFynGIj/A8ST9giXz48NjGwXdkdlfmOtMakqI5UAdEw7O+J/48wrbIAD
FRanhX7l9utVcLh6/2wq9aTe/OmPn71msc4sfDKR1kkX1eJXDlMSw0A0efBX7oYI
elxHPH4s9gLJ9SzY6NySl6QDcVwGawhcomosnZ4DM2Z53dYJ4ZDSFs63HVXt1MoO
WWFx+p7YEsHG4O54KLIVPSfZQ158iH5HNvgQEiLJ8MwyG8toXVqe35+QLjk7qAuW
fnQgAJbzfuLFo+FxE5sYTQAH9RmERTxnmg9AppfI/+xQM1tAvRMl9WJ+ujDMyzDV
qNbMhvpu9E8ccbcXI5q2CJVrewrpiKtResdOOTOBLwCBKmhOXFQoWrDio0M8AUHR
oEBMfwiRl20ZV3+LK+2sp78Z/7iZYYrIJ9w55Goc9moxfBigXyAuum+zEHaymU4k
sIazuuFEDRLr74DTT9P1XV637MsFxGsXfcwl3jJgrU9vunnPUwLXG6F05xdRC03+
6/EaW9WYchu81zPlStfrCPRg30Bi0Hj0zUEOmBuMq3Cwr5B78urSZYnW3OU8Q2Sa
M/4f4xhJ2Mh7Mjwld1JAPNGGd0b5M0wboFLdgIjavgM23gMGGWesZNeYeVAmqRIU
PBRGOj+1Xtc3XLQwD5xXTt2ooltv1lUC9IXhz+Tyx+nrbyyyX6uny+TD6gO9tVX5
SjdmwmoOj2xONo4WdFN/hbOLg3bZ5dlaAd1AeNSovTpRutIvtjNK7vevCF3W9QYq
wJIYalMvbqObI8bX14n3i3hmBXszjnujVNr84MPIhBlHXIJlIjSW+iop57UQxljB
1aVHboKpq8IwbP8L5gos9w2gDrtWON5kQ+Ls//1VZz7gd7jrxnPG/UInjiyzuWq4
yOTPgdENnajKdaGNbiBc4xrNNv+MSujTjK7TSDXn/p28qUOjMdyroRxQzlUDVXce
q36+eTVXCVtiV/2mEM0VcX4u/1dpgwSDi+afENNeQj/eH2QvnV0xtldFf365AFqJ
jS0/p9hNcsmvRmZyg3KbIzY9axiAxOcem1UneW7NOw96kYRQ8402KBKDyHvHJf51
TEMIoqzjxg6TsfGHvsJA6ISzuTwakx5aC9pxKZfKOPJw/8GXsZycIqxMgl00tQte
6MVgz6jcE3f3WRNh7+oPYScMgzRXv2fFB0csVI6l+uFu+TCJ5/i4ByDMMAbKG5vP
A3PkB+yvTozncqJ2USM6LOGBAFY18yM36g/c7LaR7SLP52sb69DJmRCEI+ryhp1t
WNHBVMRlCfQwJ1UtA0XZZRQxWJ9B3Q6/L6Z6fFggUi103mXOMw3sDUFFoh2YpXec
SrRypLKQLRJFuSdrmk2n4sMImyoiPfMRkayjnZNDdsZGTijt/FbvQkeRW5Ik78gq
thBCv9p8+ssCl62Z/BjH91eC5RkDne00yfU4dAc5b1sIsB0gCu+RatvYBPlVSKgI
KC9qinFYCxMUMVIuYdn+Y1k/QJ89wEiAAMmDLL5MS0S0R+tE0jnb0JUjrzeJMTyg
Y6yumqlPc3ErhwYxsJHNSjC1rnFKQCGdKegJ+AbMdCIoom3y4enNW/4C7oCM3UOL
ssvFhEtTK+zExrDaplgIrQ==
`protect END_PROTECTED
