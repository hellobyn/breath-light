`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFids6f2S7XWZOByawldt6r0C8LDroP/NaR2diZfIaMNdYDIWEIBxLouUFQ42LoV
yj0lHom75qzfsLSrmS4KZfwFYnYBJuXYTunOKRs28LASTIJLTTcJTPQzm/F5QrBk
t27FtUgcIYcNpCqN2d0RXfrEu4S0uWcgWqC3+JzRznCZBPUWkLu2sh3cjabpYpu4
sl0p7sER5ESsSBliWYfi4LnuSvIc92V7cDj7RknJAOP53Qr0ksL3cmei144KwMfO
ZyOWfv4jhzaAlw8HOz0OiSrvkKhl5G7kO0XrvLT8LA+t/I4p/W0AW40Se1LlWs1k
X4iEniA9kqzv+OSSSBwGFOiFoDqmt9WOF92vr07hpoh/tJRKTi8iMdBj3TAm6DvL
hufPt5wx+lCUo60++zzOB/Md3H+80/vHd87pxVGViFys+X6NrbKiB7tf2EMc+t36
3wWKMFWrNzQSJKrJ12tgPWrB6MdNTN6P1IF0155k+/8H4v3E9w4M3GlltDFKlXfB
4r9IKW0VWPmvTDlSp8Nt1v3GW7nV62M6aXVM2SHTUYrp8619NXhfUhQXsKffLegA
D14k26Sfdkj4PngYmrJSZQ==
`protect END_PROTECTED
