`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u192zLabK44Zo8h3AfzGFY/tZkVKak2m0zxemlzSOb35W36w0iGTPHK1T9wRaHGl
5K7TrRiO5PLcseHNZoq/hu0q4l9fzrwkyNreVeETvStN9lxcTL7CONRvYkY3FK9T
4T8fuL3gTssH5gl1uWQUzcuUY0VU9GdT13YkH54KPx0vXJWWeH9iq9rk86j8vyFt
JlcIFOJZgthekiXNI2reM3tOydmev5dYQW35k/8jkqLa0nWj6NMfkgunRYra371L
eYdWPYEVinF0u0aTCqBbkgvYXrUbyb1pbvobvd2Sp1eD6dtRNN2DeFYRkfFRFAMg
TvQZdITx+C3UETulVmMHda41lBvuwx/Y766eIOuvf5J4qhA49YzMCaAdC6s5ir0k
soMqLbdSPheOvKDGLivjTnzT2lkjG3RymPrd+gvYdyQ6qHdFNriA6hct/nGzLDDu
pUl2G+AjuOoW4KJXJafx0IvfUVaTPtpDpIRRKSY66wQHZ1oalT3SPqBWQxVd+jxs
98fAhgp/deQYS7ty+JMyi16ohfPhCxfAcwIaq7XUhqCCKufB1NQQNuWwUaVBbAqY
4kZMEfZ3pmCVJ7TK9SbCey3QCSUVIVs+EiHuRtDbXfKRYWSEPIL+9DOK8b33ySDa
ag2T8Wb5YnOq+vJYkcwb8NLM66hWvjy7/zF6CB98Je1nKjfhofUhyAEcPm+W7H38
AqPekK1q4PUlnGyoSxV1xM/IFMlyAAcsLbpqVywCsoB0rgXzCKaBYm4mX4zYKAuE
EEoVdAUZFH1t2eB9HIWRYVM0/MqPcLDxE8KkeX2GEBLFMiNEkIMnnUMoTWgvnJ5k
hDnoW3PeNzJPAwYK4gV9M9wVFBi/WXQwsG9iUuNoEpyHmjYB0tNxhQe864s6TkO1
SSUiclOWbZ5HzjR50ZhZhLa/9DY507FlfIjWRw9kDibgald3YGarbNIBRln8B9ZE
IBmZsrkrvks1kDaPaPwt01UCVrZ5AEpEzbMo4kXmRm6aHSXkeDzieN3r/4qpVQ38
`protect END_PROTECTED
