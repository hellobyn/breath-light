`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXLPUKRmTMJxxy2vCfg/oeD8mpoiFv0FdsHmcDlcWzPN9ozewpYuIfaa07qyjmfa
H5D+AD8wIWNY0e5B9wvZ72d6XO7naMIIZLLXwjhS7eDw9ab4Z/x36GsKPSNf6KNV
0h7nB8rSaIVxA8V9ztzTW7bkutbOYHdA3eQ1Uli+nf5C171+g/HK4OkvWmPnxkwW
n9VQk95iLUZoLVHuExBKiQkSl99WehDw9zxjS8ejfNOkgUuA8pp34ZXuDkVOfopP
FZESxadOZ4A3nOpNydHCKA==
`protect END_PROTECTED
