`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0j1VvCTCc8H308RQbdBYIVe9WEaYQALPfGDe97ZxvQIz8jMSwErlwnXUuKiblYKk
hfU3SWEz8Fs0mDBCMkC9DoJRMA2MYslYd9BENX+5FMCdqzG5HCKIPPDrNFMG+niC
sdrv1zedqtGj2m1GoTNDJidZkyU/NEyr/Vg+irkJiBzqpv24C0Bw4JAiSH4VTn7u
I8TmvkLR+HpUGV0O+Ilzms2EGTBHitEmQL0gh1RqWgqlyMpQX9khin+ZIhfqPuZ1
yjYha2zfXX4EDHyqaqs3ORkgC3z7Qsyp5ivS6hYkfeMxG/f0ApfvlXkVkigUM7Sz
12Ci1NCMyhcXDkvsmhodNtBlcSA6xjAMaIBC+UEkA1POhD0jVnRynZb7WcNWrOLQ
LfxIpx39gYQitZWhPLD/XGd1Xa6YmlmhjLdD8elsF/CfpxwqZeCOWmEo8kHnlK/k
3GpBSqBANwuuWf9Tc5b3EtWdnRgELXUQfW9Ar6MnyVM=
`protect END_PROTECTED
