`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbAJSThEv553PYzHsWsAPAUrZfPXzFgJ4G3d10DYWy4nULdFw3a5KQWbYlg92QpP
TCLJT7F5hua2YYddsx9ubjDpWZqKCl6I1HnEI88g5ILK0IY8U0oTL3RkxErYjt1K
KDzdKTvDngFCGlYi1MW7cg6dgTcND54/Cgus9GbhutpdNsLHUp7kNH1qGDHnr3eB
HNwG2mJqZNYJE7LFEP5QpkrhilmhChcy1Uix2M8SLF0l0WyXCAtWLZYO0+VDBZiD
rKW60cVHeAdCuewmt8oWY5hvzoXqW4TSWbx4f6oyu/FClQnj1r3yt5UG593VEIsn
w4nRUy5CeyAnp402bYTYk5cazS/QhnyPYDBdkhT/mYQCWhcmh0HKqBZLDPuuNJEg
5oSoxyEQzlP6uxNvWpbSWQUPD0G4HKpBy/l8qkgZT7c1ISbvAWBJfJrutVeKNxFw
Jp9/YuhterWDgdy/ErP7jsYbQoiLUgz50v6mkTEGxBv3M+CY3Ks2L8NGbwmqRU3r
s7uq0T2HiuCeknoLGklb0nB4K/DAQLIE1ETzsXKe0poS6eV1lwO6FUOkUl1Jo+1l
a5qg+L3OB9zO0Uj4hRhAfMFtLLoUOA8fbqj9pphf1MwgbiGDopZA3/rmd5a/Sdn6
hXdF2QWpykhY9rXGmA6H6fEtHFNK/SjWyJrnCVoqbksy4Zos1qKzK6BfdOduOyUa
UfYKTkElhBmHmk7hKN1lqgWWbnvibuurxfu7XgJSeouNq6x+beo81DrSETX4Sd2h
bzl4AN7tPtsMliUuseAPvQlbRvAtmXKliloijx8IcIDUaNjMBXCRz7sl/0Z6YBzy
vEhRBBwz6smpHO4FTjfGFjTGuSAb940hDTYHbZTvulJQ2u86oFKNQJGPYOTqXAzQ
bcBBoUmkyNh0wkQTSRx+jNmOTTkSiJxDhGQhp2TYir1wguz9lutohPXVlSoEq9Rv
4L+q0QGyTs1JucfPvqxfilzVrdCbK3AQ+7CqUa2eBR2HH7+E4vDGLJ00tIKM+mKj
1w2m6ORuB53FF1le68K/9ebzhRiWj7IzTo8i+snLVQu0RWlBXqYr2PFTxGxT+oLz
mhwSFcLs8u6em3Vfl3R+pR7nNp23eZerdrqkB9c+WMD7DvYsXspfWsGG57yExfuR
P2rM/nmo7UZPo+mf/lg27soo7P4gk+Im1jIyeAqItqLbpaOBd5Dj1J3EO+p0cpRt
Br3hTX+pvdsQOw+b35EFE7o0r2/t0seWyeLs2I1bjswJ4z0yJr/eatqbX9jWteQR
/k4ebAfFPRESiTFAR3f+RibW8JMoz6wdcB7ODsnbkwcCLNJIcGciVFTXfapq2WnT
AKysJPGsq6oNC5qjU4eAFN7Ma5Q3t3SGXpgPrQbg1sejcQ/Axl2z12f3F0wD+o+r
KBKHTjS4IBSQNLa994FYx9X9dfI7VjLBmAWGEohcEKllDuJ08SlqvjEJNxOq2GJv
L4Gh1JZ4GArWnjJ2oYTzT01SHJ/X/yJFxGgu8TPBl9pzDlBus2h83I0pNN639XV6
gWJTo/4jAqLFUU+FQTcgOc4tD87SS10Khq3suFJXDk3p9h9hmmdU7NRAPFYBVvN2
WXf+gc5yOeDtHV9adgvyNDTY6ZUsynXzJjJlqlAGd8PUiPHH6nN5sG+3gO3rbN9G
N55nfLLW+QOTrFsQYKIUZnr3t+4taqIcGO6CB5z/9B1Cyrd0nN7nnjUrjEGKIIoZ
kKhflX2qjMGFA922KjhqUPSGtNQKpWnYHEBiK6PdKFxAmfV9etVNa5m1co7f/d82
kS5oxd9UfvqJ6dtt5a31+Y9fftAOfRbJR4a1b8EUgITiNcD5WhmHBNY6KOVfjFZT
`protect END_PROTECTED
