`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RWZJ5INAOqa+6H9EwGEJWYL5xD7iruB02UWM6cTRTIHjhVU/alzhFJYaa98fqveh
Oez8lquAgBwNY0kzSKFrE9qROHbfFZT/Q9QwVhYZBT2xgKOqd3fmMAeMKUrKw0E7
vHa2EPajr9lWWImPdyC+2OW2uuS6OniUXNbVa0WSuIDizru9GQ/qr7hncDPu5wpz
ybymsW9/wYUGztyYZyWIvl/XD3ok7kkLWW6i55ys+7xJuE6d7TR4lZQiMqDqWRfI
3EdzRYwg4nIQPwhCzQZOIFSBfbq2VxXICOT40TGZPMgRdYb0qJXm/0uanyShtdZ1
PbLNd2ABOCzysLxMmSzA4w8q6JyEuWkbUIIxJCJfyLzIg1M4d8gxj+TpBk20QCdz
fnn5EtI3nEkssx4ZyDm+dm6yVjFl0gZnsMkXuqYNfeezDMEy0r4vQhKzmsccGa38
fgnZkefdPEd+OVr0wa+dBEn6MQd79Tj2IOCBdZpt75VNTNZVNCpceOTV6Nsr2cUG
eMw+Lk9xOsjHPW3txCwCLSvEt/dmIQwHkUCyd8/CEaYBKTWpGJPwB5woDaw6nvej
eYi2K5oCSyZh/JaDIB+yrR/PPszhA4ouMGmeWEHIsyOvNdsVaumyUljYX6POD2iw
8Kg1wlvvpDh1VF1oE4kFuo6pbCFIaod57G8i5VsyBfLEollpch2CD11/k52eKlF0
+xcvtJfbg2HE/1PKyeryw2vnBzyJqTI7u+8M7vggbhaOJXpdOCB4Esknr/MFGLz1
LHdDw2pungAdaKi/pa24VqYPYj3U+834peDiWUeWcPGn2PVgwe1kpmi3uEmGvvTL
7VpVVikPIEsLlhLumzY4vX7RTE76d0gr1HktcTXBT3NClQJxVbtnARHACUf7jJrb
L+qwRaLpyMn5GO/O4zZ1r06DwY1Jr4+A0qUO0uDtv2j4J/AQCd4e752QNP6QiBvn
Gg3q2l0Upl0gr7kPbqrteOfRx7uHrG0Q38VFeMGAvbQc3s4GPFrEag+wmJh/N25z
zX5AeH5nEqhff0ccagd7LqOQ0nokCs0ZiZxTU32c+TpfNnz7pJjkmtcyJXla2KMz
VNm8wKzuOIB+Mr6LRSoMV0Cm7T2YlVpeA0idKL5FtRSMoSvDBaDNDaphVb5kWh2o
1IZFs5rRF7qmCpUnjFN8e7OFjj4AR6Hs9zYmU1CWB+FhAMb6S8BJjHOJb29FwohY
UcDl65j5l9jamCQlTt7+dXgfCjCx7QyXhhcM+b5bsPCrtwD5VEk0M3y3+PhsjL+H
CF0DuhAX7TFZUUEVXXMvEFrx7B31JzkZraR9DGZ1du2gZ6ZR5/LVSI2uO0QlDAxR
nXmfIL7PPc00Ykn2mLS2hyFWfObTFiaHeQf17H5LZsuOgAHc9u3vKOsKIV7eyQiz
DXzPC/14g21dd2/MeROXH+8NcJSL96L7waaAaRUp6yMgf5GWiWbX7O1mtmnit6Ak
v34WQISUxseiT6MphBbuaMt5Byzl9CMFDo2P+HWiUB9/ei0Guf+9CXjHXt4ETfg7
oBnU2DIX+2DwkkaNONaHalwPJxeIG6Tiy5llRORZuHPHeWuRjh7OypLG0Mrm0nqz
GiL9qoxdcQfAcgFYQw9r56g/ZNORS0jk5iHSdKnM4GGssdtumWYHU9O2UQerJQQs
w1McPgPrQjmQMxdXdZxpI/95AlPHvAvW0+T+XmoQd3oVKEGcEVfZqQwIAhLcbsEP
oVyapSR9G+fQyk0CEzE3eVa78/EVSbX4lUPRw/g99KkObxbmugHEy5fBcHb12qMh
Yop1cCBFmiT40RKrJLqcxDbEkAY9BDb74BNnEcJGvtN23A7ueEcbwumwaxAVDm5i
AYITcUDHhm4CPRnVkO5Rp8uIuLLi0Fw6GdLRfycrkGguRBslLqFUlrqmsONpwbl/
QqIDpflmDfQ85Q8O3c7+gQmWgnxvfW/r/XMPYhTfyIB00gjSQ9FUUICV5uyV/1cl
FHr1D/Q2fN+1WTIxLrHQ/ThJsSAGbEcVDfvHJz2qUrvoBsJ3D37sVaV6gskupBA6
GY8ZOJCMxMN2d1W+TlS8fiV27tgq4pf4LIhiHSj6snS6wB/HAkJgLbUo+3ML/Drm
8KQJm4ykezDfq4/NJ/brKTIStEnoRB0ZiM5NAImoGb41WWaqHhekzxoq1l1lE0Ze
ubyDThzTP0O7l4TZ74S38zmLF5n3caDvyBAsSHeydL5m5S+6VehZkWPijUtK9VyX
4ATST5jxfNw+FiSkb7gViYw55KN1FnMq908euslQDsGrfKPvcx3qiKLHKlrNFkCN
A0t2t7/l8G7D1LdjIhKz0c41OUXdcbpaHV5Lsvaf7jr7zqICAytMzOF/k1M7ezW5
NuJ5je2fxAfRwENvnMaqlAr1uqArVM+TKCnwXGh85r+uIps3lPEathx2wrO5L9QU
t2JvZqgTVuYC0qlAatzBujyWg4+IxKfNc3cG0lpk7MlmAsQiKazCGVppwY1+di7j
iBcD4WlX7tL7SB+9gabt6IcQ0P14Cf4fvD9XFLhzQAdNZc+8MQI52dY1Q/mSOsk9
FN+dg6llo3RMnwtjAqBeisgMawAOZ1KNhAzmo0jHYaWxsg6Tp7m660uqpVT0lb4k
uzfznVsgtg9XA+6KESYGBDNaK7sZuAN4PF20aHFw0qtqn2C3lBA15dxlGTqzwvwQ
++/MOfxkovG68z+aJrCKct86eguPdyYdx2FE9zuzydkiWVBgud0XB4J8L0eblD0o
kvMLAVq2kPmEyy4GQ+hQw7mt35KRFLlvjGlyFRVwJ7Bf+kblhNCfbzoD2kocctSN
cnDVqtJ/VdgS5lGIXjZPTqgflD59E5CkmnJtrRc0p1r3GuE50F4MtawnzrAhZB+n
gr+1R+u4P3RFxlPJmK54ahAFupQLCt0aAlx7ejjexHiRatH5Yd3qAv9BYUuwc+XX
dhrsMCoMkNwtFWW1nesI2s+p/ooM6wbdsb9sVDOCqP4blcCvq7YCVVHYU/vJJEAN
XN3h5pIL+wCAFP1Dc+6FdtXaglHd3nW6+i3Ih0SMOev3Aprbqzyf7W6dM2Zyf9/m
/cDC0ddMeIz/b1y/fJyO/uPgLqgiIYtRLSHzN0m7bs4BCXed3VNeTYWwVg471j9M
RYn/bUARW5VZh95IIgnvR2gj52eP18P1VhGClNoF+mpNxI2a5arp5OvIAy0nZjbi
R5liQrbINlA5Q4uQ5ZhjmXx/WLjkIu2roztckH6mskfVo89Ryx4aQSrZVJHKUlrN
gyHsQxhdC2iDPSahV6+PWzcSy18hZiAGcI3VtlptIWWWqfy+cYLNNvrCXnD1OAy8
WpMbmsohlSylo/84/jkbD1o3QkbwOjVnb1OO4zjp0MOM1pI2tpXkyYzHE5btjFVd
MstUAyU88wS6Vg7XLluQitgcUcyGkb4givTBilYmiqsck2QIUCU3vTEeubwEUigP
iJJnvOp9hTGFUq/EH/iaXXPezCX9RhywYxCIHsu0eVvW1uJUNCDG7jqKaJdiN/s2
qbsXQbgjM4CIWcagkSKX0eDKdykCYvS/7D0iPeBLaEi6pn1Do8BzBTizKxyRKF2W
m2PSznKnqsvTzG8a/JvAzq+D5i+1svVtxCMAV9DMZihsiFRVJ/1fpGDdyuvgk89C
ncyZnbX1eNDGrv6FWHIdL1hm090PJX74ZrwS+lRN23Bar3MYwzi2Rdgit1lD4SyB
9ea/B24ixN59iohnjoex1eFMt84OqzhzvJG/5/MgpVCln16OrnqVvYUWjgdZNzHe
3QtBbDPtHQg9XcrsvebCFM+nhAlsL2teKVB3ttOeNgC324euRxT2Ft4OPrIIyrV4
hXL9i4CC9FoPWxGKeVx+FGDhQVY1qVuzBf0cSEwatLxpHlA6S8dfQwpN2Ebfm0ii
hAdpAV86rJhpQ5MwOgm5HaBQrgsNxac2zsJDAMS7QcEUTM7NUH6IpWPzisb13dNz
sVIZzsxLF2fa0TqYmEWt05fIH+9zBk7FyMR4vOqLJi5rz6d/A56pPYxprC3oq3Y1
F/INtP48eT2WU7kWAzSou7kOTUH/PU2XHV4xCI0rVx4GYI8NB1RFIkcdq1jnJqxx
Pe4pdsVKfXwsaciw0Sarj93MV8QcacGkFysBqT1V1zy0MxmFLiFfVXATm0uUNGB4
IbAJORKG8eVNVCuxmk6ijHFRrI4VYSl/WmkMeS4GOrhsmhi2LinnW0VNRazQJTGh
qV+u1RaIHqOHlaqPf4E3g2u9GxFcQzcT56D2YE+SHP0=
`protect END_PROTECTED
