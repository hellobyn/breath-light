`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFu62lSql1pmzDVq6Hev0JGXsJrsksyhfjzSDdv9iPuLEcFcjN9s9Ev7AaP2jW2B
XL6ZEkU+79BwfroYtdWCd69lj0IiE5IalmI7g8kWC7W3SyIAbIhegf8AY17ccSpg
KNl5bJ20kasTxZGx2/CZ10WZzx25mYsrKWg4i/88I84rlyykmwFIE6gZQilJ/LeK
p4pqrAfE/4wPoBbKDALrA9goYE/Wrd01c1JcuuBkiF4YKRuUxr3TPDM0XAeo0jDQ
ztih2Jf0RGiCg//TgQm8V92HiXEiL0M/DJySgg13D8TMUlEG8x3dqjsX+pypt67J
bQ0r4g4h9ikxmFtzyqxt0GKZJXTZCuT6bWZUt6lxJtgNK2TbtyYg3Hk9VypSLs+U
84tnATDGABQfEY9zo4nrKwoHd3lE7V6S7q2Ix5IOvw6fZ0W3wuDa2K5qQgSE/913
ftEoOPl5A3hc2hi/tUGNx9pJ66CBOGVDfmGVYNJNpc9CxcAukWOFgG71l6Rf03i0
Uh0NJ969RTiXpDYNTNua+V5IR7+dCQeHYY5l4iSvQ3Sk8gt3xVYNgr+666TiIoCK
gYDSmOCyG9gdpJpkVmqWqwN1ifSYV96+P3Fxt/cbDtWNi0x4RtSQ9Doj69U7LLyq
r2+smhPwJ5ZGm35qxrreH1FCyEUDM7HmUPUURxJNsSyCallAq/zYvAI7UujUcIZF
7L8LPtYUMsZjAKHVFs0Lo7lTUUaWlgkgiJiPaolH/i9W8tI4UvpiAVIXU7qREhh+
F7Xs2QA3XP107tvvupbAG/kFj+MTWMkLMq7xBTZnMC0N0u5MqV19Oepk2NL8riK9
xMzGoz719yPUWLunygw/dh4vv4oyTSYGg885s15Vtbwx83vk8joBGaxPMmhGiMmW
1eIRcfmOxhuiOFHvNkX1nrwbf9ly9XyPl0wzyIocir6XkE8B58hxoldATEKdupz7
EBtBeLyPPHg/ALPC+RVQR+xIbdYFPbUlkyX7N6I7+xSoGRCtwqMyKbVWskVfHoGG
MaOvmy6PtbJ+0Na4WZdn9RMzQwC5tIUyV/Pja3dJF5h63iYB2E+g65p1qpeJuuz4
tXA9rAtYmYUdTatShdl+NVUizZtIeWxnQVImHuTP+7G7CT5NMaPTaenGNSwVpgqE
a9gKP7mIvoiIaofGKgOgdE7BIKHQWAjicadIXdCxfMROtMOf38Ev6TVDRTLyybov
jxh+9HUH5v4LI3JKg4sgNGyZLvb/srlfDz4wgrwCtpYKURTiYHGWTE59Pytvokrf
oaRrYe10OgPsqH3H1f07C7H7j+jzRk7rKMxoA4iJZ+51fAyHYKobmTKBeDJMoPs0
V4f1E9/52hohBwMt6OJN8JGH0pN8Fosq2MCxkvr77LgaruSRtau8VCGJWrA7p1vb
OdLhlsLDAqOo92YmQcqn/AJANW+VMgC/EU2A35dInZwGs+ymod/4bR2sUDaSWmlq
UPUWo/8DSmnYdiomvdx1BPlb/eT7p/0665/tOCzvavxkGSziFXncF6VWKcPKZ3Uk
s2CBq7ebsF540035v1ORP+SOV1IDlZUYOCKXKtiSH5SAon67gcJ3EjzOZ0CDUSBs
nqnVel8VWPQOqPY7EV3MjIfWRT5ZG9VBDMZqaXzu44F5+u/dPYotP7umcJyRCTrt
CICglDwP0RuVbhEvA7aZ34GwRJr0I+4rGSHa8aFznG5NHlHOczzYqfgfMCtK9X3H
U0Ke7rfwEc2OYjudHxUTY3jEx/lbOG0Kr3gUNg9XroAqQqg5e9HzPY8EKmot8z2a
167ufZSdWOhYr7bGwnMCK+wadWI557Ivrsu5CAN0ntIiYsCEGoVXzFJaSnsCd6I0
Kytyxx+RAwc4V9U6RN+Znq+/NpdruXM9pCWzkoCF2TifuSWNWMctmJCuQjlPCd7i
e5IhHc4X9oIZhOCDTiNTOQbSjPT3wyI+GzK91z/DEy3lzePw/X/msTiCInb0a6VQ
GtDTSjKo518LYd4iDDvsmhXej23M54Ua4NjwADQhKaHU3NBIMV6EI3rjlB5woyCV
XAS4Y088jX+waGIpgdrBHStrwH11VbxsXt0EuWaGAdeR41Z5ILWV8fDSBaFrBs8K
ruV2EE+RWoocSKm4NuYSmBqEJbNjGIGtqEpoyT1GA/SgLeemslXYB/77iAut5aHO
uZ50CH90r/j0Dc6cTQUdieOr0L9kFYsCdEV/z7aFaNKC9oedrXnJxdgZMyE7Juxa
B9uq9kuVCTi6VVbZGl19rvveWrywuFQ6+LjCVfFk2v/G14nkPquXc//Dk4Omd8K8
rsKdQ36x3N78MJU2agzDC81BzYy6YmbFkFz+k9P7GQFvP2vvVmu5oYQJYbfJ5mtK
FAcQ9QMLHNgANM4foTM48tI0pkkmSj5ZifVkMn1E05FypnDsI83bVvZKyjj12gnG
KgPOxhNvc43xihyuTQTiA33zpZm4T0NGRHXpDUBQQH4TQzXUcieWQaiWh50k/5KT
V88KwpIcQlXrrjw/iIiZaAlHIbK4yeB8byI0DOU0nQ6rLvBUHuIdWUyOZ7kvlkmc
yjpzA2MIzXzHCaTQQ0reWgWq7Lpa/Z2yqqhycaImMhSbxUQS9rbBfbUrUFiP8rZz
mxAMhVmM7i4UTesU0iYcoQi4YYEUZr7kWg+1YTWDdSDmB5qPLfu+SZ2ObWhP2E9p
b3QrB0fAyNDD5ilHKmgqFXmbFCyhUcDAEeq470n9cVKdO2blqh1u2l7pXG8GU817
k3utgXo9GgU0b3ChhMvfCvQ4XXn60+SrRI0UZ1t4D6fOdKnVVjAGC5OF8D+uUVW4
hL2MNOAYRYDNuXH6sgapA3kS2JAxBfK9yo+XKvOWAZbH7ntkyWue6V0GJseNeL2l
5Wp+fXYim7lOYBoOBakHfvhWwOLUlbiDE6i0/KZnTYgF09E6Z7qVY7ljwV8O5hhi
vdoG56KONHM2agm2/cXjie7vigcK7ZqHMq2b2QEYhAYVfrar4VVmOynpqKPIthOq
cEjy1wjlId8f7eybzXItnEcBpEnuiaza/BRX4n6gCcnobf7cBuS8drpRHjdxZz5l
/+dbnWWu7t6CRb3pRWY+tZurNM+X19V7J5crVbdg0/YezY8u0/+22QrJsJunJn05
qTS5SjcPMsbkccTx68v0u7b6rE5Zl+5Aue8XriyXCzFeklJK4fX8+01dYCp0fqLV
G/cVCPJCJ2RmIoMQIL9gSWdW91ZOeBo5l25F8XL23ecm4pqk6JgmgnzFk2D7s3bm
lQS4PSBgSlNP0DHR35mTjB13kMQ/UNi0GaCGh6cYi3qvLNimEXrrbhJbSj4zkO3E
kSP6P7ZxDCKLyBxWGbVcIhC0pFUDL4XoYs26S/bJclBC+WUOMqoEChQtQakB8hnB
42Z3Rx1ONpawo77ED8I8EO5zo7HbIfc2iTbnWe4Vg63lmoyvvwCDW3ZyRumoe0kA
4ZBj2/0T1zk3LGs8DI9nRnEVQ/5gkG1tmlRRwj4Yeud0gWfUxle/UbS2KSk1xOnr
dDX3b08xkpe0EM1eVawHaB9/8045nDgTpnLJ5abwZF/RjrbDUrOFATugkuh8++BP
7mIA3V/ZJGZ4v/3R4LjczWMhgqhz10+ZbFOUqFDWnf09eBRT3Et9nAULgvyzVCjn
71uAnnB8XVBOZlayNsa+8H5vGozql9lbsLQuIN2ESJMt+3TQnXCBbINQPr5ytejK
HJSnnAQK3A1KuUfrfgOLa7t3Ro1qzVDHnSy9yagHtsinHzOGcf30iIfe8SHWiyQ0
xiTMqOh/vpRBXaiy3uRsXc1ZRAIOTpBXR4Qy424N540Nm1OevhSLRQjaB55jaNlL
GTuiN2VrA8Skr+3s3gRoaqw87dP63W7f4kr5V9MA1ZAaCNUuz7l3kSbVXXFJ/xAx
Ab33138qmHmCARcb8vMlyGM1BdRQrnUmx33ff9dia4jWD2X2Y+ivTd9D6jZPCvk7
UgFeImmDQDDlpz3zg67ZzCj1znHekHOH04I14u28kzrZBuK4zkMe4Bu/gZ1mw4ng
y1kfxOwHLQAt+T2b1NrPf/rOYo5asdsctyMS9vH+hKgrECb3DxZb0vxoulpJFkfE
gmTiDX1Dl4qfaD7QZYP0WJAVu41QHfbbRQ4HqeCWanJzVrw1D3QkWmcQD98t/zgP
NBCOAYq6ZEadpRbUKssOAl2j+l9CsgCFm3MctAiTGqHENrVX5cqhGDyI4gc3W6dX
Nxf/jPVi91ICmbggrhr5EpU7Lp5PCy1uPV+AM9dRr2yRxIVYbKnzce32zR37+4MI
GkVjKYwwU5s8oRvPaVs2a4xbi1Pj4iAt7F2swO93I3LQ6DTWIR+5JO1wFR5V7lnL
2z6cQ2iHEJ8kl2BFLoqSaZvlx9VCCLq0Oc14R8b+82zHBIdXbTOW/iJX3HxXFCkb
cuOPIafdxtENMQKx2SqdmrRL+89STyZs5xWkXe8mUstX6r1XzDvRsJbxqKTdLKTP
gAzkmEHUZbgvIRZNRJujLH0aFXFe2elwu/E593fvH7d7wflXBNSq8Z1NPtw/Um1h
imNuoC5Wqjtui6gv4nZE85INl7Nmzd38ZHstqKbe9nBk/lH3D8+OG/jReT+4Bhgb
jTBzgt8ew/8k1rrEJfxvSQmc9ACw5gMSVoF4uQcN8AkPNAqo1kR/QmuhUXvWKppt
0Tgns3DwyHCFgkfrMRjsnC8gse9gAjVRxRAKWOFTl1AKiqM7RqyR4BVtYm9sQinA
1700UqCabG1lgpGe6f5YBRSeupVcjP/C6/pq+r4ZTbXo6ToEt+PKm/7J1vClE3wB
ruiylCs8/IxooTj/yaANXhaC95583ETOiNb6CjjTHYKSAPgWLnZZCp6vwGRQh9tk
8RLl4x1mXQyKg46uJOATQq0mDXtV5poGnSx4k41P3Khb46UEaPwozeF0siZ+YQfH
B7ScvMPHCDXhr4Y495YjZ+BkBGyM3bcFJscJMtHANz33AR/VTsj+movRqeJzPm0+
0c3+AtX4BlePiU+Wvt3E4wfXpv8yGjRjvjxJxCOqq0ZhzHswXjE3q/gLTHcEJo0w
dShAYPGlQTLtjqoOZdoHCvSxw9RBe50kcvtZP3PV0F/OaSEfVi0LCQRjav/dnZHo
PmYVPHZQKuxfMdy+egI88klGu/s4y/oB7Ozum6BTQxJKUWE9htV5Kw0pFSdzrxB9
jifZ8GFDPagFMjxcoYWLm2M9k0oHWkt04rWB91FaG8BLo/NMHq833mEFydZSpUDu
WaFhC0dZSEf3YDDU8s2I26cbvwZtoWiycUb8jlVsnSVWiIyIfGC8uFkad+zjKW0N
cqA8gJiTwzymvUs4rAvAjsg2ltNV5tAtP7P6lp1Wz8hgHjKcvSDJ4xfsxyUjPAl1
QsfaotJac9pb89MpdqBB8Z/bq5/6nJiUN57pLrl3V1y3cl6zeZAKEMuPWmqq8VUw
Ghocws4PHDXtt1P9gjybICwO5ybbcmpeN28EVLKEaCLPAOZX3tbatcA/6ByWUsl7
xfIhsYh+fe2gayONvuCCHTttVo0+8osABcwiB5kdt7onyV35BkPI2eRaWJXAoDeE
z+yCmfCSsHCHRCZKZ2ywlKmym7aa6NRAaMGb8ehwF9Wvg8lXikvohdRP6R6RqqsW
v6cyHWcQfLzwr8nWPH9Lcgt9Dgxno3u1c5fbcz0tK6SNQN99LuRtUS8fTFYZRzfl
wxMG6tibgjT5U2C8eg8JB0GGn1NFyWjLzxrdIJ/3CnFtVgHpzEKbf5RlCax8IHYA
cA3/W/UuvHptIIW4AEEe5CQtDpxGjN0+UiJmxiKvtHoE3PXkjCTKUwobI15cr81O
WlZpvkEHl80JffFX2mwzKGJoz4vB0fVKgaudJD/u7Nr2hqL2phkGMdzYvmPjfFOC
a6juPxwCn81YSR++unU6os6pK67EWbu33EEttnIIJv+yOyvRnjQzxwTVYMulQAwg
XZEbyOZynnT2BBrsyOo4MmY8W0GVs/XfBmHoRzwZVneUb44DI0/s0qEypIsp7Yim
lOGRwR4bKLmeaNc0or8TTsoXiMmSYfwnLRSksOQXdl6u2qEn7EodzHUXpxnv569d
bP62ydykqTaZb0eQ10NXMRqfkvKyrZsoCSmfs8A0O9uDHi2jiRTak/mXeoTUppFc
u3vqBNwvAPYpYHfzpqkNpZ50qIC2ijCQe4roAuiU/AEqSzyviOGn17oMx3krrB7K
UShHXyu5Zq7PiaaEKdX6jxPjm2LrAMQOA01cK7WAYcYzG5EJWO68XkyWwuD+Jbci
pgjQsxEh365gnIyAohjK2ONvQgvKmIt9Seri4ax9nxKw7Y/yte1flLlfveiwmiKW
irzpgFgxfVRBC04VpkWr8Ua4Fn67Aaa2bFR66XAJ22h15RvgemPVFd/4HqWFJ6p0
lv8JhHWQuML+WnvO8xb1UsoZWmcYvuhs/1mqdEVUE3pMFQ1oE+/GDzQdCl2uUHeu
HBFrSzlPwAAN+KpmL4VlkdtA2rD8imv0+l4H2koJWf15iDWvEMh5lGrn/SRNfEVO
`protect END_PROTECTED
