`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqWp4EgBgayh41p3IdLCB+4eoDXGpj9FuVSSPWkr6dXp5IxBiK01NvtCyNyPnWQM
66YsOJoe9L/AehHQY/0IH+iglSzlpfrgC1MK1nzBYQLBH8RspdqZzZKC3WF0pS/z
ilt3+D0eWJ2nm6sL4oYnkGED3x5nJnovdhazF1dVvee28FM3vGuvIJfpItbrDBhu
xozgeAn3e/P81H4Y8rgutXdDDPvl3APIrI4/GXCZx0QEnIRCAbTwCVHkFpQ5Xh69
GExPOQbmREyOA1NtN1SD46S/6BEPvpeEiI+SsWafaEBEs3YulF0ngzJyxo9WyRsR
RB0nvY/ySv1Ml8w+IPQXV7AGUuBKFPGX3ouef9sMeCFy0f14ve4tu8/qG1BW8IOs
5q4P45cRDySCnpUbHEtBnHoGBE9+gqba8vG2RrHkMtaZafy1Z45jzulfUJRoiMHQ
GdEv26d/5cwx/PPY0+nJBGuUTIU6nhOnVG1/cOvcCBvnfuaV0kTFdcKXuutmjM+u
CM+1LkMrNgjh0eWs8mmj8RKQ1QBAy2mSbygSu9RUC14/FMvgh8ylhgtwmf6xuwt7
xMVyX6cLABHeqL/Ru2tzryqntAEp9gfwyjfxxMfSPGdd8927pTBZ6NngtisP7nFc
BexVblXASj4HDM8LczbbPke9LsBbSbORacKu6nPCverPqkZifGg+At2cL8fZW/7b
9zvaM+nKMSjRSS2/2i4ys5m6lSKATWDO8GUJbfpOiDYNiwgKAvw0hwgG6pWAO9Y0
vi+b2+4DuToDm2NRP47oUUp7cWCDOhPlo09OT1bRMcLmYhDZV8UaFOAvY0+kwH0E
3E8aMKV15MrACjKer32iAVRYxqAAiw5Ff/BAdM0o5bDz5E2JZXAU+AZIuuQrHHOd
d5iT7zqB4p6kI2ibu5f6LUttc2Uppaw7J267sbFw7CZr4QBoYBuPAUeb/jgZgNk2
PyZY85ciWRUgNtI57hRRwEHkSvbf/I36kz37ZcdPJZ4yWTbRc9d1wuEn7pqu1MBz
cqFzidEhL9EgJbAVQo1cl3zc8+hLDqbib0i8dTspms2APZG+SE89Ahw9c4/9++wf
LWjjwUaMWTR7LProDd2ZqKiKKJyHZEWmKvyQ9cxSa4zqeFZR1WFxHzGjyvIYOd1R
4DLC4bGKtCE1CL7kEbJCRk8qYVCJhGed6fQzV1MK/VyWU52/4g96ie6P2fzcDVkx
bEKxYsDuYMrAHHJ1EAtq+r1hfmIuXCJ1MFBVWsBy2DX+vO+qmjp/9k+ElajcSCnD
eOS2SOAzIZo1H0yovToKhhsMcKAcGFqT4qf8VZJjzfHWfKA+2SrudTAaXrkxcqCQ
5TAHQsYrK67vF9VtVczGrTco6XG0Hzu1XPauilIv6tBD0WmNJ2ylOK8MAQx6Vs5A
lb2CoJWzsuutXGPE8E+WVJSf9dBWTZGm2JTF+nSL2AfpCcL76LzeYke4xXvl63Uv
U2OC1dH/FaMrPIdZLqwnfUB9UKrpp+Wxjz52bzgJy6rZdiAC7uMgX4FWOz82JGF5
Z/UAuOioEEbKRCLlOkJ0j/Cr8Yyq7fqVaaiPnpJ3Mj22B/iT253VDynQzTRmggLn
XOJhyw2pcO5KJM9az3rMcI6g1vfkXf/N9MBe/3fswLo7huLKsUu0w2bt1s/ybd6P
Wl+0Y0GOdT+IFklZdMNxX0jGJI2HryiELoBv954HjWt9Eet644E5Kf2sDr9d0DtX
IxcftDsGWYOa/D/Y4jiG72E10lXleLTXPvMTNg9YFxBzThAL5PvmA/s7YcA0favY
BwRbuLDdSVGgLElq2ooIA39kmi638au1KDTK6c56TmzAjNxxwF7azMV8LnYRJU2O
gNS636ifn/zPTMLAuEt38ncZGGeprViwQLvgUWZRRLAs9PppJ9h6wxgkUG5mfOLY
ngOUdkkdel1nVlBuUxh0QQ==
`protect END_PROTECTED
