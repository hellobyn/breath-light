`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkyKqTh0gKIhuSSGo//lLrSUIsQQONuHerSmWwiUjm5WzbnWH3kd68FyfJ9jvn39
7qmq4i8HxJmkjQgPc7OZO/IqExDeEChQpQFOwzk11UDxUc+gTPVAY3D/5dD+sqL6
riT+YIiPxfpqDysrDVhB77jO2G905Ndqt5+O+5kqy/BlL1CCsYCo0e/naHep+t+p
kLpNWOa20PrI2VA4+17BRjLuyq88w1YcSeFFO8VkEmKbBrvIAr7tsvRSOEMuKBvs
YMKvY5s8SstZJmifQMwGvSWhcOJDVw8N1JX3HG7MFq6JAYFYSMZDy94wiGhqea/c
UP+7ta991SVDcyMWUqFDmxLZThmBfILzjBYbFYB6cfNzCMuioWpZapSMEyzwLHuN
28TUAHn4ndn0tqdZ5VNH4mqU7nZaHBmFLderJfmOe7Ksx0Tn6g6QHvBtXp348YK3
ZRxDs8s6bAtjhYUclc8aVUxAY1HRB9mU/MMSb6rPhr8j/ipDm0ZHuGum1/r6CXAa
sI3D7XShKSD3zEDjd59W4QNu08XYZV9StNY2RqWZl0SFDF3J09iPEqhHuLyuzQFN
BxyBZmp4caFU81Awd1UlzM7hfedbHQg4PZuVie8xEwLm69nUal2zzR0e2RFnclhb
gPH9PlbFpm++8QFpi3vB0Bgom4O37MYChzRZQJ7GE5VFkJTxCgz8AF2t8HJ1/I4u
Cb+dbk7iIL2a89rIPmT7+VN3Zx1NYt4WIoQrpunlO1DN8OKyzJxxwT9SsdQwM5ZD
4iYdKL8j/2FhuVx4PE9/pnfScUJ91epJN+6/o3teQdzZ/DG06ncyJuyJb5oECmd/
goegcDnTWryaceqWRpezyA==
`protect END_PROTECTED
