`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3XP2u1V0LZRTWNtuNa8uqLcMGso5wAwM2257R8jol2gh9kv1X3LkroSvfcwRSx3
q5hUZlxh6Rux5h7cHT0Hm9n31g52gIHKjpV/km7fjkzJfEVner27VsswvbWGj3Li
/uM2nYnnqhpD+5wEdxHmmqOHpzAgvINihiGNG0Ay/2Unj2MrvVSOnN46UBDUWAYA
8B0OD2DAWXReDlMxUdwCYT7O6GEglqkHnCb5ne89cA+/IMwNID6G83daXvXUpLSG
owqGg/eOp2XnCbivdSaB2rDW1A3rA6kn1umkJrEdLwkuCcNwB23iiRNE3EnjBdp5
MnyMp1XDvcjCvZS0QfLef/9F6181wWvwHdTqkUCd+KpBxd6IDYtcATlQAwar/qGN
mxDFvC+kHh/qb/Uv9spuFC640WDJXmjMD6CZ4b64cWchG+XRUMOiKK5cUnCjU9g/
Z9cJWkVOWEw0RXZNR3gSYhEFvqBuXW5o5CpdbnBWULvM2EDfcaCDPGMNLchmyltF
RFcijqgeyxGiPwro+NT3Fc8zec7zfdnhMRuPOJEf6VHr1rqvK9uR/zV8SWVDFNlO
O5t6Graqx44AkFsLUr1sMjBM3zQphZtu8HSQsQVQTSk7SPwP93lXv8ofUgoCJSal
Ah+qhpgxbnjADTscGiHfhmLnBmFOZ2zmh6qomN4TXoyanqC4X9kBOGyDW41rM9g+
tTmgaf2C0C8VN6quyjvMk18jpjk1H9IXCIX92lE8R50WQBLtWv7iD/rSnNgGzdiz
IoHZtaV9JowwNMCkiazUbyk0PiVSIGPRd45fqsrGiuvnFQrM49cqECFitG5LVLep
6BABwFrtedVvR8R7vK3uGZF8rHex0vy6qodk9Lsm2RKJxDJGyJfA8QWcmnXyqVVl
m1FTR7ff0hksg8ulvMiQTPvIAapOnN+09WtBabVpkOKYDxJW5KaBro168vKeI/ap
z1rjtvvGKvpONGKYHXp/7fow8AIJZUpIvIMkQbmGgxKbI8At2atiwv+BBpWSj7rP
rJO+aoeUKjJARnPNAuZScKCUmTW7KE13Rq9VbYM5DUT+vg5l80EwUCXONjoU6l9S
Yc/pSVsZ1GonsDuSaq/2m4d/Baz7DVZyZ+4ZJ4UYmiZSvSDvDDsXRBkKmZSy1tvS
PifxeweZAOTdhgcsuk1E62xr3nb0de4kMypff6Kt0K14JL0YrgG2k5cypQzmVPz5
B71nUZmVBJ5ZhM6xlprk0yboY1B6FPogpjnuqS43g/CZh7nj9oNKCSNvkezksQ/x
9+eTrtXn+05i8ZXNDD9zO1FQE7X7vIl/pXTFdzfYOHkxQonSDXFKsu60BIx6XIxj
/RMGVljx5sBdgBcO6iIubKUsry+bCpAePGBaMj+yOROS2RUoMjKf8Z/VRcBTJNlw
S7mj1+jhnWDXxcSaB3XmQcJc/QXr2iIMEId/tEWHYSwkxOtouZP96nRB+gg5DKP8
CeMy2Z1eY6WiG+OoSlUc6lbOU3neT58ejgjxe0boMRbfzRDuCq+ADgXr8dD6B1Eg
udPHlEUEzLskxAD1bZb+qXcP+wnOzeVlIXGOADlKSZcX8Pg6DHn2N8sSYNmnExrW
ML4HJ/8zZWmbDXSqlZLi7TiKxVQPvKe51TnCCW2bmsxDwj7GdcupuaVb/I2onogO
pKNQpamSYKC6UcWnRLNMRPt13JiTNqWo0XSdCiuOkjwEiuJ0kQi3acbYhhWXPjRm
qtFZ1B1XW5eg+dCOh2DQBOimH0FeIYP4fjBYK5x5pR/RjJ8Wm7zZA/mWuLDGFi7Z
HvOdEHz444BwO4yNxvez5Ur7yLeJdn8GebIrjOuQItZLQyf7n3/rtmfx/0T19mc2
gWwC/kCj8+LipSrW0HSu7broK/bZFThX6jEsg/6+aVbOyVSULcRiRCyHPCF4O3OS
I4AhqznlKXSbpe/umLLxlYoMTeDbfHBmyvGC/KZ8MbaPy8jK0EvHyuTI/tsD5v4x
rGWPKGo2KO2pJpruPMHF6N6NkYOsLWDw+XPYLawCZRCY/9A6aBERSulD1wQWYNTK
ZuXfBBBZ00TCoi0K25+Z053BkuJCLwCepZ5uoWYF7D6y013wQC/jAc2zHfdSl72n
3lp0fLKPM/N8shhag+4WX7uxAnYmWGEhjJMHbRr4OTb+hH5X0I1F+wsg1HYMb0Df
nY1fhlbS1StTyn/UFsZDhzlvgMCNFjheFrUE6fP9/d+gyO6qRoc63SjbUerdzXKV
WBVB7zKmywGfZ3Wo/zhG4gXXa3o+2d6HwDogXefMHlsd+E/dPppfd7EsoMgsr1P1
E6z2PjNbFRBIgOofrjP/ycTUXu7GZL7WWoKpvcYvI8Yg6UyUeyu+Q1I45Vj/EVOi
JIKYk+ggWDMFeWc1U5cAxJ6F3odk2S10cWI1Vk8Lrb6aeDVVtCOIO6Bgg3QqfQc5
FRmj3OCEO9VphZhS3uIsZD4olm/qZx8LpbRyt+79PJN0t9+Oqza6ONn1Q0hCUiC+
kX8G0Ryy3DYm0IMS0ZINX89lomloq9JYvYlQKfWWbGkWZK5yORa697vJxgr9/Qc+
rF3xsEVLv2erB9geEfImaUYB6eVP4K55nOf2i1elpR1kWc9hkp4fwxXO+2rmLpdQ
KNKThwc9WNtNnFq254zY7XRjTU6XeEH5ZGlqZ/+dwEjBOG8F7meU/ybPWsg53ZWg
j7Gdgy2ghUuWOtOoa7Y6Apsoneptci2uO8tDzAddcE0utUc0trNRgRbRh5iVBBFR
da9ROgQV7XyiTXNEIG7l1JJ3SCbczySuu+N634Q1jNc9Rtqy6CwL83EsfcDW40fF
1Nlp4WjcDWrCKE0ksUuJaxhwaDOlr/+DK+llrio/PIV3EGwV85ebxocGIJn5i0yV
ax0vkqiwnBHeXisUwiTkWXpsOwiFDd1ORy+OiXfAL/SCM05NS2CsrKHbemo7hMaj
3mcuqI2Aw7K/87O1HZrDbycFyyKnbpcrCKwjdQsb1XJrs8/MrvzL34gnqPGyhgFK
91XeizR8Jvb8pHHcj9UZG6855gSiS6xeLfR1y96zGb89wARHguetLmrxhivJJYKZ
2cPUTFf2Yhsg3VVLDzc4jO27x2pAVGl5HnPP7ehTKi+oS+5Z3qoHYhDwL4BrC5/H
SeQEr5KKgr3IE0vOr44Jg0+Xocm8+QTZ0GbV0aaqMAYdzBd6LVxNIU8dTGjVk9aB
kCT6SiwOj6RfSrNvWkjZdkzB+JBE+9azB7WHX6DacTlZKgqfqLV0qgaJQXllEToj
kF3rHN21208hqNG8WDnrrC6Of0GgSu/ajcVaCqzwDeHnkzXCU0FalVa5lUD5K0cS
j4vMWl+yZBvSovFXi5aug8CQxzo8wq3viWDbKxRJsBR4qdxSPhsBPr1CUzXT41w9
DPYRYjAayh1/MHLhcm7mtkzUTISFcqnj398EMIEDnv744K6aO/lm/IesIdN9ve/a
JtkQu3918wXCVAWr2IS5iku0RbA5exCWRaVYDJ70SLh5KrCIdHlWWwVtOBbZBywX
jf3ZEcnvN5pRqe4zGglo9fEkmVMpEOkiFAKpzuvjvvFpIaUwsPVQE3xXTnvzqeXI
FKpgSASJ6C9bKyHBMcIB1BBEiE7ZaVkKzO5cDTqj48A=
`protect END_PROTECTED
