`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11SVl6uO8jwzVFBK0eQldPqM9V6PMLBtprKM0888W/+Menw0YtE0eDyacYGMg3y5
gU6EwPpDw1ghAU6tFJiscgBuQEa/+mAHQv8CvJ/rsYAzG7jo07HW+TzVzfbtUlcs
aNqNRXje/gpFyTCrglDc8z9ONWeLvrv3KICA3Dbmr5xQdZR8ajw7jt5pJDqo6GC5
WdnNrOf1NYMLuXkxZvoO1txLXm0YqTvFmrrOi/KZc4BJs5AX9C0kNrPlbSpUQEEw
tuvuw3YjdGYgyjBkbhKygsNIH8aAqyoSMUH7bopepbANlIUU0wi4tPa+8iKtZ566
Hg8JbwIAXkSOKzSaasLG1pgqhXLG8mAAu4Bgy1h4gm5eHG2ms95Uug2bej/2sMlA
Zilk7nCwG6+iSf9diSV57ty6yUVxJJbuI6QlUpMb0uEUWAvFEyolqDToe4JfqVDs
RSNHmEGIJ0udR3HLLAYp6h/IQmqlRigKRovVTgC6cDJ498ufTQpjIw3qITSXeQ0a
m4t22FzGT1h5gDNw4AAca8sWXrVvNiNp8Y45s6LjvsPlPfCpHx1QLWqvkd0ZBMga
lIVIedNC/0V4z3vJbPLXfkSBViBVaDfloHGeldWWVQpW78QmCigiQOMQUQWZ/Xyk
CdiYWluPCKdND14Mdnf31KMAPO286gS8WBgnMV1LSR/GAC/OOtFHw/UUenjJfeoh
AdPjWGgo+28qGuonhvKx/b1LR0AmA1owSF8WsM85KlXgjYqSXjgKyqwf41i2rxlk
WeuCIg+otVS06Jq4F+8zeB7op2OSNWzVDIFia0o5n6GsexYChtLaBCuJBptO4ord
AHyLJtJwqYBoknqu5lMoGKv8DphAThCUk+dZ5xwwTbXWNiotW/Re4CAzXb+q3vYp
RsunDiwNCouyjP5pI/eksPuqzxrWxyvGg0VVoy7o4l/rncjzv6iQq0FdhZ6w2Mb3
pBAu4rf7o0rvBnWjCaNQZVXKjoGwtn0v8r4TGatW5dIDysJ2eEVeLhcpa/njOQws
9V9pDh9cVBYuSRnM9Wn/VW2AZq/zaN5w4esB3s6J6kLHUW+nMUfde182wbB49UUC
/Nll1UB2BmX/pDfKT5gOAiAp4onRK6uVEbEtyLPVixoFlbS14iqhyJaEq0Wjemhs
MiChXOJgjacQ6voDm1BmhIayLVuLGCtn+G5ykCqQUW4HmTomydQtx6Vlxw8gJEHf
S3Bcpmmrjj+lxovS103Tac24Atmqkt2MhAa4c8cKUYT8SUwlk0ceYlgZrBsyieQT
BVyS4sH8oi7nfaf5Q8p7UAZNt/iRP5XbRWJYcixFyzUd+BUaCi2/4VmggXbLNjR1
wjqnB6V7YXdkpkCpFQRdglcdKbukRvhDxrbk4pOQ0cDsdGxeRb+6NnLqMZSzx+u2
ahzvla4AQ3JrVRLI9jmtPJQ+Q8NFxH8yCCWajdO3g9dfem3CIbVZD4egvIAikuoG
1PxxBpFKzjSnTWwsqgD5eeeDHtWMf4QCXLJsUmLqhBv6MrVSIOgYex2VP9E271a2
Ys8x+2dpaa404ZSVFbkmTXrsQIgqSEGcCd6pbKX85MYAbtN5KHN2obQLRFwTGYut
f3WIRYC+c25hdE86or1xA8xVJ5XncruO3isQy3la+oXlGR7Jm8S0d2jgZSczXp71
cSXP0WRTObOpjt2wP19xcx60cy1iJC9a5iO80rQPyqzs3IWX8Gy0szgbBjC6kMNv
u9XroceLFs8aIzKK75CsvIi5DfcmGubOFm6+VlhmvVxO13Yge6vBixFCgqHbhc3O
hQ5a7dRVh8HUc0BMe72LFn4OW84si+qw6ZLLiFaTF5qY6sNbACzzNmahi+ozpG73
R46v1g4w0Wjqvr8fZTFBTQ==
`protect END_PROTECTED
