`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHx8XcewxpH2TD0kmOQfb7Pcepi1kpl5h29st7usGxEvb6khNmkfCTN5LmnBc32o
JiObKyOAoENb4xAFiu/H7NEbZprn9q6/+PYO5M4gnu9u/HSsnG5NNbUYTnbOUk3W
yoxIRcsz/osNFIIsSpSAgXnoAM1KQ+UXa9JQN7vBduXa/SQievE1xPC1kGYfVHDR
WW9VGZk6Y1MxUt4/vLT27tbNVFv8fJsbu1j64QLqsiDXLmC8hbyaSZ8PH5bF4AKy
6TztOZv6oS4+w05t5iAUsyLT0MYlO14M32hgHSIQ5g+PyBKu5nFdK1ZBV1rbXtjO
fJOorfBz7nfWXtucalzaFcVunQb3Grw2z8oSbtG16KNhxTTjErC1P6PIvQA4bfC9
UT/KF+1wQ9r8YwpvrchygaStk57brmDSGLMMt3X4YwxPyVi3ze5Tliy4TTWFQG6+
6kRJhbcXLIosfwPM+VQkrDbpa4nJRZEBmrABBx9s83QvsVIAEJ2yQbp6/1kU72K4
ypyOuAMPtICK1eftk5n+jMPBMhINwHWPPM7czatWjwdRuSn2PNCqrSqNs5OaEEVf
ZHHNBOLu3Sh6NY9RzNXdmPc0F1H8pGmtsx7pbmfLYhL4ObQ9uKO3lkWuvEUPJLOZ
66zUW0B4nIeGZovZoC4/r0A8jW3owxGxebshR5lvbuZoPUlWO+rXrZvlqPHfgB19
xrwo/1xwn4lqaw7aXJykjjtLbcG49pGMpOOGgD3cP6DE9rU7eB4gqCCQFznoRg6o
eROZPEVL/S1PTcoFeOKeu3UXOmOdqlHq0aIRz+wvfk6tw0etImGgbnR8wKEqg8ig
BO3Qv4gU9yu376TDGjhD6vgTQrPhOI0Hb6ZTSvnjM71+sjxjNs5Tq7XW/2BN/KjE
iGjxq2gq9G9emyq0g07B9/IJTM4DlQmRLCrTHyF0YcHi9iMeU2miXO7m5PsYUqyG
9SaK3KiZylXNLWgw//2gdS3x/W0SLPqbqpp2QiIVPV+tkEaSi2bAD1HrtVdkNEN3
mONzYiXf3ZtCnopz9nepRRyv6UhSvz6ixCDg0/48N94EXMdqymyrzkeVIm3Pz1Wg
3WFtNsMbIuRL8WgP9G5sqrJkcvBrBORWgrcVcjWz8W1zRNWIIS57iaFJjE/greV1
5/VC6AF/LJQPjdrC6cVl9gbEIi+bVGsxK5LzwL/zXoe/ez3mQR+IMtlj21utwdYy
mHDfwLwdL6NN9UO9h9h+m13Jt7lkVKWyxDTuId7cHVzviij+ZlLLYUQkm2B5qS1+
V0SgxqhX0NrhaRMMZ2TMXKuCHbINT+XLbF2LYelajQpJNetT1ROXfUTjsTrhAubf
XXpIjhESceJV/AcL73wKcEvGVr+XtR8Q2pJ/VHZDiS6h8D7CfGlCD2C68AH6VqQx
XvSdtG6vpvIV5kU3A+2wWXteM5HWQIB+FBhOX+nb2RKSGmpZQbQjadalcZPnSLhr
SRup0YbpprVsQ2YXAF/jaqq/rOlW58kj1HZ7W3YGAU/gVM59mcePJZikewuviHQh
19JkZqUDNfpo2pcoaU6zWuc/07hLjKNf2JqnGtUNVG9E3+97gzUBiCX7YEUmzhxW
1W1B+MlYrq+weTHaXcmRYnLWA27le138UDN9uUoVSVU=
`protect END_PROTECTED
