`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PLe0utk2gWl7eudtD8jclRxoVQ+wkxWZH45CzmzRvqunGCbB02TEtsjG9eXTwv/
X3bW17/Z2VwdHwX1tHV9EuxRmh7d0x3nmLwPu1gCOhFkPlf5IA0MWGGNIcGW2gHW
ScCHh6YxcSoJUaQOyrNmF8VtHtaKRZkQ4jrH1dKyKCihrQ4es4gwXVzqGLhRfDEo
7vtL4GpslHHYyWHOKmUs37Z7VpZy8yUylBRPbFTYNCn9Yl7HaI/Q3T1idBe1riVD
iD/hRvieddHOM0hvrSjejXxzZbTOPn/waY+mWyjubz6JEmtSgCEvNruLOyVkXFAS
H3TMczjKCJrpB3hXidX/F5A8hiSoVm9XzIL2zCmJlLuHS/hWhEsRt/UQWJEOPupd
KeprvfTLPeY8Gkiis/uNHP+tjy9yXL8Led18Ref49f6uIAU1deP1KYwMGUbI65GH
2vTo17vbmz29XJ0kk8snkj9YHHix4eiXZ05SrQAWr417M7hs9c92sq0mH2cF+Kkn
z19qrPnekISojdP1n271WndoWMddVOJFp2020gle4EIvNxNT4lS6DvJK7ZXLYdUP
zUw2qCwDTdGZWkhcTo0lw6v/b1lvulGfcmSNrUkPuk/1Ms16ruXdvBQttRTmyhIC
kyHMz06DQzXuDtAb2d2IqoGSaWwyUtQ8ppkhFVHYbkhyPfRikqY6rr1vBFmyiztt
/xQpUEZ/fMPSZkj82OLN1t+bRGeIr2lJqzpwR2Kbc432dFY06IsL20vwYlFfOiW4
GnPamAG7Er1p7gfsep9O1f/calNRnOcFq/rMf0HVSURYezBELTN+R5aYb9ah4TTD
sxoon2KheYIrZLmPt3+hFWjIyqNOFWrLgjcM/ZIznnyMreU7ydpiE8OFCISL2gwJ
LjnRXr9Pj+7PKbnyKAQx7CZ4npKq0Coc6ONB+i6cIoy0aG9/+alrbsYIMgMT2uXu
h9lqTPCIlc7KLj99K9ccT4L7Xi5LCObITwT9VXePkUO0a4lqapjIf7fZvBHoOcRv
Jcr1BKX86qapNyMdP/gra7TGb/Pj9oB4+dCl9ZY0ZIiJ5RrGg8kOLVX4D/KCD3Nc
y/HB4MmuFjsHVZ5kGhvAZOXCbXVGBVkcs0QSwiW6uDNthYxwW4j62bBFcl1KrnUy
WXSMjMBPmReU7C2O1Lds2do58OGec5bfFcgnWoNk1Ego3ZHJfu8bJaeQxox7QkOQ
2IwYhO0lyFyjPU2gCR4mXjSvqgzIV2D8cuGwHAJ436AcrmdFBtZKEQDLaz5w31k3
aW6nvYxfHQK4WScb09Dtg09VebAwSdm/B2I6oUYeoMBJn082px6QB9IuMaS0ab99
PJj9gZdjJ3BGHDAaF4UebH9/LuWvc9lAGOCbP/KX1jIg6unQWzINrRQBWxud6uTB
/0mfRIMGJs1WwyKvZbcqb3Hrj+tx7kFBc0Oqr+mqtH1Ek6Shp1rLdr/8OXj6zHjX
hKq8DDjnIfqVavBFg5NnlPgXxC1kEh5S/s2mtgLo8hq5WFxi+Gcujwb+ICR4FX0l
Ran/QuUMzAT+0ArcB/Wd3ywVtKGg9GThifU3AKit7lRpU302uaqsA4nkCbwCvJJj
Rm3mB4HbTkaXtNSBj4EwypxBxRG1+jE622LkF0yo3cvCP6fV7AbdkO8aTHowadsI
G7C4++04+Jn1GT9Dy1CrxMrPrKpFk1JPg6seBfAQL5aLUrvGMnmA0/sdBaNCqjaN
EP4hgkJ7qtWcqR2e7lUHjL+zCc7Z+2viB1pYn5r2CS0BltA10e+uSZswDtlc7RP6
tQ3zr8O+4xUKfVJJbCbbkwohc8WalAQ30QGWKj6UyscNwn2bFMJvrryk/loFkzMT
ddfVRVgBcwR7vS28DJ5MnZ/QR68g9dEDDxkUmUzO+GonGPjlpV7Mo7eg1+DvhRjq
CHvXGE29xRLOPuz0lihZt0c76M/6FnkNAhlt48soKWh1uX2mTG1TC3EXIj+VTRB3
xiUAMBdLkrLyzNgEJ7N6TECfA4WW/B9Vj8rlqwns8BR1K4udpyLvzDFyF7TbJcjp
`protect END_PROTECTED
