`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IiAOEsGspPFDBojPl0I6+1tDNVz48GBmjiw6p2aWID4wHn1jo555GllbAqZjjgTB
l+UOcWF5eqL/2BCu0x30jqn6u/6H+8Nn4+AljQFMGBr2LC1c8kEY4KsgUdPw0j+X
BmWd6cVGzRA/WkUPwy4aojfuHWWsVQWlDQtoFzANf3jam9pmZS0Hxz5FVTYVeDHu
qr3rw7b8G9rseBloP6hJALWRjVbO5NVM1H57o24OimU1JSQ44SBSdtYCI/eBmCWa
cvA6t1fcX3Cv/LtwSYBsWsv1MmydsaKxRGi+3DZIuDPQ8O/RegxcMw4v9ex8FENu
RKm09U5Ii+Rd91a1i967z4OR/8hi/rEAnhGzGUp4w4dBsTpfsnMLRJqAx3ozH1yW
PyhzKq3pvU5p/F0mIhd7stP0012b7RqZcVhose/fEP23eEP7daB2qFR56N2ApueP
F6Tr4lQaq/oUuoAimYuloCmwKvvNHeMLL9Oy9Xbcw1IYW3a2tbXDE2IfA1hLnDU7
9RnhQ/FtH8BxjJq5uke+nbhbbZEsQW4cuw0Rg/GQqfx/tAjaUk2dzgeNvp3r5TXC
BfW/CwZwCq2kbOrFkwgWXdk/Z8Jz6DmPH5K7/mnNfJwGD1dRdDFKYgHcBQjnnKB0
jHaZcYYP9Hlh4cEmgdOji5zFmoexu02d58u1czfie/I5xigOzvlNodmOltGyikCX
wwiPMup7t3RIGsjQF/XPkB4CGH0BXaEN1/cHTD67rS4r6A+Xt3qPC7Z//yEbhkia
B9S388pUaw4+JUoY9y0Zj36lFWO1Q0CRC5NiotPPxEgB9upXK1amn4upnqyLFBOE
L55nXsC0MnNZncdUnSZbIywkDguKNgsd5hdI1XzGnsadPhjgcUN8yFE/LB4KrFAh
upd8HYwhx7xBx/6DDZecnm3agl/k0jfBGS4X/Dq15bZqx7ilSRqXNZoHTmTcx7Om
CxZ1ZrtZvjgWYNo0OkEf3KaGByQjrXtF4lL6IO2Uhs8czgxu9fWwQ5qp8vLpDohO
oOKBX0U7B3Sx7rVLl3C3JOQekV5W+S7K0jodKy5hmAJL/94zrIrn9e2amwjmUP33
EMjdoXfq/EN6zq8M65CHtI278h2pUG1S+Tz6B847Pz17mihHCHsfiBlBt6vy4Tg8
gZ8as47+CE/XG7ziLrAd2JTQEg6Umtyaz3RZiTFZatt9ah4LqagjmHyPpQerYUEd
+2NKO5IwpdBCF7UpXzoNmgcAqm7pua64wEvNSTTvc3F3swfbrWa4IdJIGp5+zxBD
9q9hXCZFPnCXGNLcANfuaI6hzzDhucBfOi9NDNVPSEFyqSEtFy9uJAMpdZXU1/RH
0E+KGY0C+S+ih5Wu4RIng5U31Irrmk55266qusjWpb+yB/5/WU7g8phL8edm2EJV
j63T8hBO3MVFNlEzI9f7Q87lBdreZm0MLvx8psjvkkM+zuohj/6RSvlCAOPOLlcw
2XIzJ0Up9yt1P3pmdecbnLh1yZ1q96Y2ippnfRvYIzpY0INpUSR3sgTzgDKm0goK
o7eMKeGaVscLXKC8zwOY8RUBtrLOQRAks59oPBkj3QyCz/ZO8k+iPMA4Yq/xUm78
ITdkvrZY0mvthmlg+68tIlD8LYSeV6VYOZTFMsSuiV62gl3i7eX45Y19Bz9b0Qmo
rM3cU8y+3UrLlRf5g3rBh5AtORLpGP2a7Z4IJNKgzLMIBqWX7Da8R2ShW+0fWuXA
FNOmGUCXTQ0BCHmlWm0d0plo+YC6yXxBbAG4xYeAPlNKdTh/3t8oF9Yr2l6AFlEL
C0QgH//R5jYTaB7bGzc2WCxLVDm8iGNrhuAYPeFYoANMIaZ7x8ZEzPRI86UHTiI+
RCVVjssOquzFSDZImyCSsPWz8MvwL/g7pxSbTO5Z3q/BewgM4pFlI1fxrgT0tyyT
xrAM7Xco3GNE2mAXWnZ3JycXEIdZatm+CwWQZAgy+cMoYW4zncp+Tmp6OoV/oekw
ACS5U/0qG/aWPLTs4BhKiewNDaRdW48aLEp/As6dj0tQD43zwC8J+vyNnOGhHtvf
Zj3BwqgUHmBWGqtHZZ0HGDpJ9yg4ZhEbXGqVNPwdtKNpw+2gVpZsUbfNB2wDK6/Y
Nw1aOjFn4KMxtR59z85herVVs7MRVVT6BKdX8bf56JoSaboZW1E17V+oxG4q/lJP
cugYEttPJb5SMHZWGaKxU6w4mgzVqgKhYKswjJY7l1gKUwF+h1XtrK4xUnw1KvPo
vNEVWTV6b3EPl3zL0F0v1sxIi5+PCyLGKdFOF/gDkIdD29TfdbbqX8EjYlz+Y21o
gokfHls7Tx4601W3B+iWNftJhubFDEp03nk2bXESb+WbHBJnLikAZsHlFWgWep+b
bW80wxwsafwWcu6ayzbgoWYGPPhTo0ocdnqF9yaZ2nfcKeOtdSd6If+3HrOPDbDt
+ug/Oa3lJ8Uvg+Fme870KpnBXH0dJT8xY0h29GTcEiI8RZxfuWuaFW+/alqCxxfQ
ItCxEUaxTqQdQK1Yaam8/laIM5z3mvb1H4fBTUv3W2K6Mqdrun58PQQ4B8V7zvcJ
p2IQR+68Yn9mAIzb440PhnW5iqGmZ8ayC3y5BuqK1qblYuODJNB+15qg7bUFdRfF
tp3PgMbrGIG/VSVYvAeCIP0pHddCETX271G84XbJigmv6s3PhvMFBV7jQi1bnpF4
DHh664UsXmntIoUzqLUtNauC3g4yuLGEnqalWTDVLKkPHwk++wTjzCkouAz8AYDD
a8/uLKEcX1xFOmqQsQxnk9MICXU/dXJlPacgxW06x7UzmIkwIyNisGFhfYmDSZqp
xqCPNc37Zfy9HVxJdggG1PhTE+ups4iE8YR3Y/OR2/kf873Q84JDMiueT0ByKbTP
8dMmtp1iE1pkb2VEKg4PfByiF8wkf0j/5sL3RELlHteNnnd/4mV2EOj2fBcWE9yU
FN+0tzATvwR6uJq+W33Rw3Z4xwcee40LZma/F9kT/6OqxLR64U02x5suEKtYSA4M
csMyotK/TaVsxrR+LTZ5I7AGdKG+th5+Rgci1ewrF4p+cGABsNsq1lXvMYd0JtbL
Xd6kg309M+4LtXnHT0zOSgH75D3Cz5+BFGREvCDw/OzJ+4IlsIf7n+rl27IFCqiO
YYBYQ/AVQcwvYS7vFsd5P4dazMCKYPskg/e7z5Kbe2dtD4R6Wmk9ziqP7s1aG8J/
UQDKvy5k+064ZaouIj/ZkF/QmMSTn4zkGCKKrnTgxz+gzs+wQ+tuI7BfFZ0YF3lI
p8zn04A3+wRMUZfXf9Vt7RkfoHhJNfVwZITFdPRVCP6AzLnCjHYVue7NpAawUHeh
vFqk6FoQGoWg0fRG27fc2Zg8NC7HnYG0nAwHRsi1WgtJbSYlKfR2B5GFew4D//rM
blgEAoAUHHycM75qTwCvDqF9Frkp4eKelT3Fk10TdllbkVPGQwxpvT/++i3oV+4P
MNDwoNCdBnRnORwvpdUh++jufYPubT4wnDi3kbsF5mc04dYeSbVpbM3nLyBZP6pJ
wC31V5gl5hK/e0ynnG2V4P4P3BjpoRUuU40nzb2I0kfcKmLM/C7U649NxvcmDJPi
BQmRxnN6als3IplmuCNz5KBFONo6NvOPwn5YGYxuTJZpQboqDIawH3z8/YMvPFjo
E4AAxJXO7wYkFw/IJLB3WtDBQpNQ3XWWOpeRgwAivKPiUViX903jA2vgVsZNaVjM
vjgPOPLjXKUyfyM7cM3v+rcJeYQcObO75z5ZXdKsJ9xhsW5DDA/EQeJiwxFs7X3n
mGVKBCEDKa/+5yQNqUFIhkIzyNutWCLCxucOZKca9QZqnjF3xf43sk40xq1+iICM
M6o4qWZZjSkGu0ti6X5RX/ajtQMkkbS8RWPXt4U9qB5/SFSOBgC13dpzBskX57B8
9bf5bwHxi1rjwPvQUmkVdukxU/nfwV2+zric5e/BrMd72WebGl/qtMFpCb1lAYCq
ajzMgfThzpMRjSyedp88Ea3fBlqF9cOgytb+MRxjVIRiUdR7Zx1bp/0WKejOtorl
PxhLda9/1V0xzpLpPjR47+xDBE0eaf0TAdWsWb2A+7j8SBowTxNNd+jI6FbVYSEc
jmUmGOyA0aopybu2ktctXnF7Xd9ozqBtBHKIjTn6nTK+tgQ5vo9wXaDYeqXEUjl4
oNKeZMDS/zXQfdQc6FPMdUaGOSGh9aVZHStrwRedvb96dI8O2lJgTjx3dE49AjgS
MD0a7w/zPZRIgYUc3g0fBkkH/vFllvrrJTbyfAdwguK5nrSGixhm4TgvziGH2FfK
1e+OGI4xOi1TPZzeEwAGfKgRUfp7fTZWGaF/UH/9gqSsyucbUqdpbhPDF2s/LUNt
1MU6kNLafNPe5CU/VJDi4MIASrwNi68c/nT0k4pJdWngkRgI6/tPJENafx7TIvq1
6KYs+CJcTlT9ZH6cH4zBKn4hNsued9HAJ5xpyxtUAqL+V5aHTTu/3Kan9ufGo6A0
vSJ2Q2D2Xawa5TEA0rRI48nRTNS1rtw70tz+iEzxEvgDXh/nUfUDA2dZ0TQ6DVcG
P5Sf7whtQ1KrEd7FPkKfhWJccPRwAOMoZykvO+BE7g0H6ZRt9Ddf+HCbN6rd48O0
OClsOU1v9LvWibkLmGzohCRhI+xKtI859c9QMJPp6+kCTn2MbiN7VJDSIP2fRhGp
x5dauJPNZ68bM7RRuV1trZ63KX2Qf7jTW0Oc3g+uFD6g476sebB+/YRtGpSSfaDH
Ukr8tMuqyduRTkQoUjwcgZrdyQtlqGY7qqGlcv3jyAh0Jilm61w5OoEN2I+KKH8C
pJgGG9juEL0GKCwgQsq4VMgYIGXFmMHklHwJQ8LZ8w2Hmc33B//yjON6lEjoWTou
1vRJ3E2iTyZiae30kCCVpf8BxfqG+rqdIkQndwZICPpSDNUA8N78l1z6cTYD+eL8
CX5tct1Nq7+DELsELyXrJ8VBIWSj0/gBiO5ep2CCN8ley/zFBJ4Tky4xdyNa66q+
MMjrVrK6HF0nDBOfc5y9d59/2+Vao/6VwEB6DfJg0SWFMVmzJ36CcHMNFU3UaRF5
5rOBV4o1rWvB4L991m/2IklHIFu+9VrJ4CfmX39Q5XWQzqnL7T5LVgnsPoI9GceK
WHmDG/dRhmw9kw118ffDzrixXip1BRFaeJY/uPb57wDtO99anTNODuhIBUxahdu2
OSJyB8CMVHKH7z+Hmd6FrYJquES0K8IwkVutVDrAnOx+GNh4XqXn5A5jnsDdYTnM
Dx2DGNkBDm1H5Cw6ZnMHLUbWhris2M4GUrsLqNwEuwqwPcrC3aUmGl+GzvkEObL6
rePL4ItRUuRw6yupCKWFzGh3eHiM3KGm1IPGJPZHSefulJoou4qmCi+qyxapvOqq
eYhAMmLB24C6I148Te4YVv3QBZLfBS0tm9NKF61w5xBCa/NwzPbLemVGDfyu0GO+
Hlo7bQQNYp7Ex0XoWebllgwqpUBNVYz7zkYBX6YjYELqztXBPKyexiQKeAVQhdl2
VO5g96zwAJ3KouzW8Z/4Cg2OCDCJg5MC41w62J+x1dsSphkwK1Ods8bSTlBk+E/p
VYLkj4OgEPwOWH1SB2GA6r+cGBQAzJojkCHEZEMmRcIFXKcu1A6nugnYS4HCQK3Y
sxvxBGhGFYZz9U3rwdOOz+lMVm92J9Bd+UxNsURs4wv35ryOev66audluyGoAic9
L2ZIkwmcitUVgARgbA8qGhHsIsg9tCcUfeU8rlOumG47D+uM3gO3HfRtDZ6sgZog
H/ZjVItaK8ErgdzIknT9CkREip2kRdvBIFHSQMH0IaZZ3mzk7f1SwEsxdbMR0st7
1tq8iVTf9IDm+yAbMFR9y/tyfkRwds1A7wu5SV46/+TVIcH3CmAT+zrATj3jjyBA
2F0ARi8nvVFoSxM40uRomk5/MI9I1YP/f/TFwkMa8tv7z9wf9j4loD5nTHYLlUO2
Yg5wnc5LbmYDt9bQEyv232rFyW/gLJBkqN+D2ZHQKlvL4iwuZzJcxZz4o/ndZNgR
iGVwBKX5bb0ftNPz0xIn3tQo9dfB/RRV20uHow2kdtu/hLdDYY59jBW+IugyDUMX
JQFw2Maseds8ZZDEUs2lxvzydiYCGecwXxpUiZ/1kmbD45GJO+gKh2De0Ap1ltHd
DBjcSMcTzJmjxU9WzCn9vXtRQJcZsg4D+JpXIGSBScj0T4Dt8k+6q6X5OkWYYzzS
7Vrwv0Y0GiojnMy7VJt9zQ2sSB0ydRAmJHC+6Qb1pTz3s7RiDO54yQ8sR06haAVS
4VamBdbmLsFi3Z7snQ1u2E9GndDK3Rsz8wyOQPjlAge3D4VacEP5eDwrksl0Uztv
pOWAhQ1AwV3NXWZtCPKr9ulZ5XS7uAtQMS2BQFN0LtNZ1ZMCTdP5xCWKBqIyM0jn
3Vg6BkhwcfWMnUMT2NGJQuVXY15zqWAE3LQ37W3GVPxFE6aQ+xUQaUUSpeBt8zo0
T67FPGVooUoY5sPUd/nGBMPDGDXA7/ea8BtsXVgyDXlnU1sHW0fCSa/CA5aIXkgw
GsTK75fLTb7ZU6g9ttDIMzkfjIbogg8C8BOealTFoY2KWQg9RltDc8ubMx6q8ggr
40EnbzXT/NJbaUJhQ+Q7r1T3Nn3nRCx0Ki7rK5FnhYtJhQZqBXEzVbPrvNFlKkZz
SY3ODmJS0HehLb684D/n01/jIO0mAxPm8PLFYSFr/NVIYx24r2H1XfTq0qc8rJSX
HWtKe3wcMF9+dDIRglkFCgMkKV5UEb/pa1/OsGVnz6yGWowsN7K/aJ87Cr+vR4uh
Xs6iCejRDik+fKy6zZJqqkvorAd9n6wc428EG/S3mL8qzC/Z90/9Vba0td5vLZ2n
Sv6cXleI7NNN/svHyk8C3WBBgTk+sWnO/CkS/I6GLAa0aryv8St5uckdY8WlqSrT
tLyMJ8Lmq4HvSuE4kd/twq/gnFSrGyeKGFqq4o0EWVItZAi6VWvdCPaPR9Rw9vKo
9Ou2Ggh0i8SZSC+rYyPxV+5/tiyr34572SN+3zCc8D9DdN48VVFY4SWD68eoMxzJ
0ZCVD4vbZQwol2n5mXU3ZQjKvO24rpVvzFe3AOMu4WlYdCEcb9BzCdXTBoU9CrRn
pAfvG5JHVrdyHeJ4MxaUm3kWx2X15vnp/PE8WXkf0qOV1SBn1UkqaeX43uuiK98c
tdO3TkeK+wWzuKGYbjpwzIXv2ygyW9CNdE1SbAMIScGoC1YFwXIypFy56P9XHOgS
SjwVXmEfp1LBdsdA5UQI246STG6W388W+np6vTS4f2Ap7p4tu9bDpmquKNwqK5QP
ef9oABMqUjr+M3jpjidfnYe+IjLKeAwCcdyutBxkAr4l1c95z/MI/IMXwTQWsaS9
EXhKfLzQxxvXtZEg56gfnW+tZQ0ONwZ5NBnqo4Wv4euP1k88g8NeP4VJg80UDyKi
drHF2++7DAZZKNm3/HOkpOzZFWCMosT6lsIGofOOMven5u6yJEEm39unBtqLOiJN
IXk3KCXDn3LFq14bqQwDsTx69sVn6CJEJCb/pHZrBVqDemVFkdT6kmj1lyEIeiLm
NXd9Xit1Ep2MoiJoNZeLtAHSUo7WVeA016Eh+cTTQO93ZSdXUFqtaMtsBNDMb9dx
w33TF/RDHxKMJLUd2JumHkEn6jGS08upHZG2OegyHU71d6Okxuiqs4KINBDFUCNE
JGSJFpKd1RieaKajilF+xC+WPIxI0SqEAVepUoS1yrC8U48pPFlFRdRpzATdUPMo
81yOt+OHolKGh9epldK0ce8iWl9LrqDBhfcs74iCYD3gZAs2szyDzyT+EdgR+Zzi
YbKJ87D+twiL3G+GSCPi1XwtjiICWju7MU60pU7gyBPOuTaIS3DLOBjuOyzV++Er
hHspbRSfnBQSnIOaIO9L5pHiAauIWx44YCFfH1wC5vVUzOhRS3cNLzUxumYFnfWc
mPudA/A00B8W31J/GLahT3CLw67t2kiKwednHrTnJOO5PbQt4G258bwbnNNJwfAV
nFH2Thx1HnzDlCu/Z3rvhZk3eIkB1o6JEmwsQvu2lmIDoBvrgLo8oLqlPGdceP72
ZUcegZdm6U/Vjv85zpitHhkBPauN3HM+auCyXs8qMa8j09bOEwRMmk55Je1vhsYQ
XSiqY7Q2zFxHdTKH4YWpU1IMB46arphnHoRxgyUfEsI/3pZp56Z3MxTeB3gwe2QQ
9zaSXPgs+rX8fULy1RyuMN/T6ZPZjbRtESR6cWnGQ41+BkEp3KO90vxnM+KyzzAI
2FlU4wgIAbWOngFyL6irtymVptv0n8SQCsnwZzpAm4l3WjWpNYC9HdgQHRJ+TtKd
dTOEBeXu0C89zHTsb2amxxvIR5Zsk7RZeJTMfFYde1zKrlwVH08WQbX+BkQk4EUY
3PFLQR+Sk40NM54qGG5N1GRWI/qTfJEZ45n01TNJC+aryJnpz1fIILBc7E0+q6uS
c24ftOzRwtDtuf/S2dKs5Uhu15ISfZ5FcTVsMxNFoAU0VBeVfUCgoS44yykyx58P
JqyTUZUHRamLr9ajhRcTvPm4oIFGKCztuOhooTw8pagdip6/R+G0/V9gdBRTLx1d
sxQdu7Msm5MGfuQryFtbJsA9zMzO9wSqKFJPOt96U/Gg12e4aE5DuezdStEGV0G6
RzTag1Yk1YP1McQpI2gDMCLjKE0B19iFXY89YnYR6tHS+REfV2qe4Z2dLGviEWl2
BdF/HHmIXct72uEkw7M//nxQZDwxrGcW/WPlbgQXlAG1ohHhWi0oKdjU5FN1erGI
XnXb64FxD4Zkio+4gKQy1cBHYB/X02K/lnKe+g5udh3achf14luaEyUufEL8inb7
k7Od1PuAzbfj14Su8cLc45+Cjok+57jmSdblBWzKbqHqaIB/VyJdI10GPwdnWJbQ
BIesjK5ijdgppJSU2+DcQaZ1WUxqZqLbNlys0eGlDIrjhmm2vMx0Xw+R1/CZuwa2
mPJ3mpizRjRjlaBLKrfgk9J6CRAMqaUNZbgZyiF+u7Ru4ioPg9QlH3yS12eYx5cK
vRyMSOMdK+qs6rAvznBQfwM4tcpzhjdW/Ghr17MN3ls4mgsuQdHpqu6N9Ue9UZP3
zTTkJPm+AtpHHL3CCXiPSt9s2atq/f1mQOm7qC/MHJ3GPnGeN7HzDs3nvQZkIdVW
KLAF5jG6yOzHhKTr4fUFvE658mQdm67Ay3Cgax0i/2qqOmtKNdJx0cVqeiyP0+WP
ANBTBvzkQ18mt4aOMJyBdF9BV1cnu3Qim+1u0paW/944MWKtiKaImLo1KqIPDiJd
uL4pUBYH96Q2jSdIirYmdYB73Vize58yd9D3yWkaMv1ZJDTdYUObQXa+at/HVQmv
wn4600xE8oPwAzeZwKPyMr69GRjxK98UPgyHLM00UMBz7NGNTPVhvmmePx6xxlS5
DmOFxn/KGEEwSONZrO0wVA4of9EVDEUqb2DmQFeSzf/KiObyBIjSHPw8G1Qll4tJ
tPY5xqy2ZEsES3Na4WDH+rJY4wuwuWgSRo7GrpFYlvkFlr+My2c1ugj4QewPwgQk
Cs8cSochQPdWxXJXzLaPR6Ik0eSEnra3ClNwHrPDxYSi+ETn4aStha+0mcmhjM5Z
SW9SUqNR3ikWoE6D7uWuZqECXnoKqQmyDj3jXG4iFj+O4la2CTp81bpd7ZuRvvuf
d10Ab8ELlJL5QBeu3vJDzqthXU0pCNsZKKVEFv8CWxMFNK81wnsjZ8Rfqwd9XhAX
7a05QOXA5g1Rju409q+9VFb/9ZIjT0hKZS80wD4SXZJi81R4gyu3++x3wI6dxMMS
Dd5JkfuuxIeSmd2RR6cl+noXlVV+kCL3SjUecO0OIICCWPiWjS4G8Rm/HYbZ+TzP
sviqCFMvSZ/qAzo3RX3TP0VCaWrpLailbX7vlpdXn4BbVLV2cONXjHMbIQP3B2yB
1V3uWkRpoQWbftqKeX+hkuXTBR4HMg5ImT/8BDLI6pVVVkZe8KgGLr5G6JDkbsGT
cq6bT1Mjb2fNlkZi8U2OgGN/EUTcs3diihg3xigjXLl2keg5rTwMYlXXlcqVoKCq
oab2qSvzZCsYWLaMDeULq7c1k6IlTiCLo+pebwN+0XNuSf3o18f28RwaTxH7AByT
tumkrfGWtYBeoIWezJFPJ+5yoTNHlHtUq/+/wqDHk3gSax/vPEUECqCsriax7cKi
8YbBm4cGsHfZ3V90Y/dJc3i/4LmLSLMADrvi+p7SE1wasHWJjI8yQ5TRRolnZOME
CvxV3pxZZOHXLppF1PDyxnlZvDyxDtok4SHZJcr1bWDtNpax4b1SCU+HybqLDDeJ
Cht6YhNfJb7S4nGzhuLp15hbZViYLI8IC5JSmspH+ShX7lJbzWvI2Nt1HJfCd8gG
wfExqTNKZDJYpR1vQyQqM8IpAjuQzE0g3Nd3n4cWpFG03EALhFBbI9KEWqNs+Te6
smQhbxAhD212aOjXNT2vwtxxxqg28eUtMMsC4uoZUhYB9jCJQ0Tfl7R3te7AvuaR
+Wc9SnEmd4ug7rGf4CgI/JHJcwWqudm1x32sOUyYCkQ9Vhk2c9Tosb323b1PMc9x
nlcdtd7qcVhy6tH/bQjUwH2iUbwhfAborlrhB6nV5flJFBd6BLL9R4upGPz8RwAt
Q1agTcvDnuZEynRAS80SEAaQeKrfD8N6STsu2tmpBgnzf8/yNw6kjln2lM2HKGzi
xIvLC0PFbOJ+Zsmp4KVmmgqrXMVlyBAH8CVHZI2NmBAH8bpfDS3DSBJzMc/eqIWL
QCR3/bowVnGncSKfMPcbs+qBuxhakHJODsEWv1fJQ6TMml266waxtBHsEa6b0Pfa
qGh+bln4xQpLMgiKAryBNFaZ6w74GAf57ESm/UJv7tmwrvUUXE1RevgEzjjc7Etg
6FmpWyY53EIo/Hhp1x6kdyAP2wjcuL1Mk8rxOEv4aA/BfX8XVS4rwh1+tR5oSL9c
ufUWCUTqRgitAPPqTj3hPAVKSsqjxu2SVN6RhNk3Mx3V4ohEYZ8fm8nTFRfvcYRn
yEwiA49TouxJ+ENidkZlgfrCYBEH8LSCzZlZ7oJrvrRhLg21mKdL+oMuzzmTSOSN
E/9reu6PUOa88164T69Ep9bfKkBYrEMhQcwp69GV63m5GOfJQm4vRBYlJ3cUl3bm
IH8h+pF+NuQXBGeL6KMQU6IwX9HR4i3DST/e/g0Ui0PBNh/LirUXlTpTYdJnA07i
UaJsgnxwVsHorFlNTvlxuqb+VrR+5lwwl90XYXdtfvMey9G39DBifyl+1+8ut1GH
XicvonrUakV+j8TgBqpMf3xKY1ycvP/RDA1bYniyihqcyPnQK+hCqTP6zwnImlbK
39Cay6E7Zv8IhnElpY5OpzFjVGDBwtQbOaK68EL2P9Nn/DRXnRCn0f/VQgiY9IIq
xhPWd3McrVfvfBIOK2FZGItV+WsfMrHKXyI8OqUN9Sv4//w9kEUs0C2P91dL1BcS
jwO5O+dTVK/XDYMXTBE5HN8HIMj5SSGEbQmXtEDGG7F15C3FYbndkYGE0z89qmkD
G+tRkj21RCc+XRse2C+GoEgYBGgNG1QEPxQsy7m3OZrZdlVpsS2vqJUPOUyxKngm
FAmn4b54lm+gGp6dOisv8D+eLOHfpxTtB6ezbDBG+4ip720VOsp8SnFN4Y1SslMo
1WIt5U7WELELZ2tpkuA7MhCMwCeJlGqHOclp7BAiOWKRx1wASzgKnESX94Nqgbwy
07afY7hXgNrP8qHgpsP6eBwEYnwRpfsCeQ2DNqiViXNE+C4a1r/xECyJVGzCTEg5
w7sn/7SuQTABF4UiIy5WQBUPxIxL7UCwTgRWl45q+H27a9nm3rW71uRgsIlx1cvd
e6YbBNkcCD/XvVK3zTjkCXOfM0QgVzC1LWrtbeDODYHJQgBp/enqvLMXYooXu3ib
3CTOmRotXD3U/bg7SgLLQknQRhq6fK3x1J9dAN8U4MyBiYqri/79uW3G8JiYz/Xs
eZ2R+f+Mrq5o5MEGA4mLf7WjyTyV2D1u63RK6t0T0MeSwhzVSQvDSwbAGUwZbnoy
GBj0+Eamd7WPW92AmgJ5gcbm8gPqx+vlU8TBxPWm147p14zJVhjqMpCuSKOBxyqT
s8P0CnphI2dwPNnULqUrpDhPhtuZUAzXhBiSczy/3C2nC9L+QiBUxjoRRi+Gci9c
VnZx1sdQYXlI7vFRYqbJJFDpyS0bLgZuCueXa2HGZQbq8SHUaQL30hlHseNc/uV0
dveWnWJbU/TrCWxa/zPq9v0miscG9WS4LsgoQiRB7+rw1hebWjG3Rw4WTh+toY7r
X0r5erMsNVcH0rbjo2Qm4oRUEzX9w8PUn6t47LHqDER4sdqbBtrP1fghuB3d36ZN
BnKClFeHxeT4RsCxy9s5bNxK0UHeClqRkm1rOaCVM9WMf+19HA9Gcoqcv9v+A1dW
j5Gb+hd7mpyhWtLFDjk/6QnJPNPvzVl3xM6nIOdLDDh1vVjtcsOGXn9BWtvQmKS2
zCmZJlQp7XR/p38ya0gTcOxr5fpjHR1XZCH3Z1e15KRSM+rkFDmooy/s9GB0duIl
WSoGqFkl1jyTCjqSl4Rkk7Fm1tgNI8JTLG5xkYiMvY/7yVlRJ307D+LTK8wwfe/Z
c1dIM7d29g0BeZfghsABSuwVfbMN9SZOrM0GGErQq/cdiRQc0E2TZ6xPL28b6CXA
UtDgYd4OU3GhIhTUanVfAZu0xuWRLyM1rkqvec6eD8J+4t6dNlw+ZBfHW1CVj2Wf
WuAVv3TQF4Qx6etM2bASmiHVFanEIxa9fJegb68rZtFLPH0kiewo6IpH6O/eot0Y
rvJhQtojozdqEh1ez4TH5K73X3LOnKfBKzLVYueCsGdXSUs2pmkwCBfpmsvxX738
+UfEy+q+NgAk9V3EjENBdz3oEf0EbGe/7NCt8Zj1kDSu4X//S1jQu+/B/gE2uuJb
Zp4od5QFQg0L2gdODSOaBf8pu1wXyhIqC1ebpn9lGTKlV9iamo/FQwqTi9pvQ0zx
RoYGOre+4gR43HtpV3JZD4PeOkeYOVw6nKO78j/gg4Q4zJ8jgEFQbuoaOiWzLRI6
+ijT5hJSR+StekLubk0cOdHqn5pBoN5d1+92brIWS6la1Z/uNAAPQSWT7yKJLMZb
6KKIFBLK+GGiPZ8/ZQ4XvKf91OwOIUwdDMexOrWC7XB4V2j9UBQQDl7vcwpmf+YW
ewqe6ewqlgEQB3yw/b+BflWAovMlyuRB8HQz526iu7hsQ/zq21a9OkdIQqH6/20W
BjnwsZP4UYn3GJX7yLgJxT2ojTAi6LrUjPKHbdY36Pts4/NbjkJc8AY5raP2AHZ2
ZjmDX5YSnsw10On6L++SDKgK7yexANtH6pq4rnGMHlhVs4TyMJThDxPTuoyWUYe2
Onv+X+hOWwJybU35HM7fGSX8d5Nf3kcYtgzLSvxIy6/oaO5LSjzSxu/5Lx0fh1E5
QD6zSQGlep/GaJN7YYs3XcFUD9tzYcrS/e8MjcvZV03LuYQ0aTI7yXKAX7Bbp2QM
Uu4f54zYpQCcbg9zkHIKLtBZNkaI5K304AH7aTj5Q4B5D2oP8d6ECT1oiTKEstG8
cMkVG/zGNrX3uYNF0TLtBxy1tMbk/YZkNVnyX3lQr+dtTj6d/j/K0xNKwp/ZO9De
4xNGcGt1hpa2CNJKu/q67w4LiIvLUZoNUr2fff29z4aOWOvBk5w+uE9hfVVi38rP
vYJ/uNkyQ3JF9Rgq9CjGI8wn9KaBTKKWQtTk9ieiWYM1srsIX72UxoFcOYhVwiyx
Tg2fbNoozHQ/4XBxfNDvvVAT0jihGC6JXRWG+cYIcE0=
`protect END_PROTECTED
