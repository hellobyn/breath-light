`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FkaSgAveqPJVrEqsSuvDY21Zj5npjQhZumsMnZy9/+tGpmi/wv9RsRuvloxt3rD
Sg0yaByc8ceFfqgmnUiCBp7idxb3WoROu83SylEgQWDrH7QefL3YI+ajCtn2ezUr
1q66ADckHbKb/vAZXDOI85ig+WiO6XKF8O3AISlVV5Ejva9GnuZ7rRqfvRrcHWMM
4HZ3CgeCbDHZEBmTNrPS51bKpp7aAJ3N1QGITNGB8NiJN6hZLoKmajM83WIkDNtC
CkEMLy9sGva+OjNdwqgiXeDnpjux4Po26n2H6VC6SGayieTVL+5LKiuN6NxKo0i8
0LaZ0OceZ10hXtoKNHQehLUlbND5qnvtENZsxFD+A8GzEN5yJpaHN9BbHYK+FF/K
08vrDvcGCLrEFS7OPOShhDJr8JeUtjs4p9Gn2UyVwwTnfUozIQ0VlittZHbJotMX
fN25+79xayftjGaYcNs/dHEL7j3vhkciplYy1NcpU7Cs+CGk2T+iZSKS/+IMrb+4
GrIz3thnf0G40Rg3TAHHwft6bRHwy+TMeF+kTOJSRvI=
`protect END_PROTECTED
