`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9a1J90J8D1uyttTZucmBvNyB1GvSPcfEurNr30ozzZ0s4udYO+r0h46jo7KVPfV
88CLG6o15HaNG8GqVpQjLQMuN9yP9maiLH205RN42v0i5VIXVg+GuXAAMC86Q59K
h2BNPsu4Fq1e2ooLKFYMcaOQz9u9c48rACDw6GU28vg9zBQ0Dm7j5zBcT7rKANx5
`protect END_PROTECTED
