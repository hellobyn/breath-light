`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVPE66g5Qegu1+xONAYaLocRMySvTY97H9C8ru8hzbmgJyi2RVuTccMxujknDpmK
s0oGsMa51RrB5H7/415woCCgCQAcN1Oweu3f1hmvXbNx8a6mxRkQZ/jEE3QqKP0Y
lEYCj7n562UuhBecnRc4UfsBM1gA8KPiaO3tRa/QUZC1CzQUl7EadUb9TSSpxveV
mKjhLLoc2AfLaKrdf5Iu4PBMNOJ30Q3IeVjskwbwTtaUswwTFJGw4b+2B2Xo8ONX
1IVoZfxMpjlB/0dLqyPO/Wizo2gmrG+piiERcUemtV6Uv21qYJ5G6DXKxsu4Lawj
03Vub6HzttfQrB+dP7nkpN9fdn/PXwlSzwF0Wh9l5NVgtf4ABfvXvtdaSDffMFkH
toCROBPJcD803tslEzdl25DhhZUVtusnRUUSSnp+3Od1l01vrADAcb43Mm7FKzOj
pGs4O+rWmwgIk4QKYuYQVglF+Bni1gKT1EwbaXsOJ1AI3XJ1JpXYONK80y9e32iO
71dgRFM0w4LI99utX2glKDwL0+V/AluHjOENqufSyDcKBenQIhvlDVGzq1/YrDdb
Hvn6F72Sh0+2BgG1TdhiTWrQczzV0yGS+ZrXdsE5isBbTVbecCIfzbQt40RXb+fJ
PXKxhjrx6icpHb7WyzcGjrqtUoKqrlYBLKtuDrXNA8boGdeRd14H7RUpdBp8vFtY
kYhXmLBB1G/R456wvzowMGVSAp34nXCuDhKTWTS930pNxOgvr7uZ1pr5zdcqj4Cm
L00uDkxPKR8V7PvdnxwpejCmbMlKJQhapftabv00Hen0+Z/JeYHBejdSfHAI/bpV
LPi5c/Iew4/T5z7m8YSezsmJs9YHVj6lGuySvnvR7RlnoJ4GHToebx30s2i7g34I
sF60YLkHJ60clykomowXTSQ6D4tVUmYMVFwW20gg5WGcbZ0zPTGlbOuOpmPGEGsi
OI+4dRvv1BdB+KBuEyydcPcLlxbaTEpguZ9nZDZ/mmgNVbPGXjPIDjVfBYzGplW7
Iu+2LN5qVbmLMqjalw9+wHdl28vFODRSIyYGJm9Ni6WS8YYcNwlisPlWEhn34+XD
UOAG8HTYMf1hV5nFUSpsWkglEo2c25uK010zpUFkOLiMiSJJE5tYFQgh3NDlNbxC
0otjXmZ2R6X8kmZBuXdM7yjV6ob6AmB5nOEh1ZzVvr0bxag360jzuveWMWIZE0x8
vj3U2NSUngMp+vHNpAnxlQ==
`protect END_PROTECTED
