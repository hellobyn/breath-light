`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PKSbAaRr1aHmBygW8lEJolJydcsMx85q8IT7iUR8Zx0Bl6bg0ZhmfVDjqP+UvZa
HuOAx/P2Ucu9iuBLeqEcN98mtDIRPlGIVcot1YhoC6QsRNIcfki0CLOT7R5BWZXl
kjtxkQq/jKe8LuVogYDI4dCAtPHlKYo1VSoxMGx4SE1WrHJjrIOSXeg8fJgykZuM
nTYAmet/INHp1rcGNWdTENtMxo4nhp9WS40RRLTJ6rK8laTJ7Hi40Hlyq+bhoWMj
v55QXp1bIa8fIhxuMOTVQ2vr4Kv7LW6awQP9r69nzn+D+0CPfUELkHkTNvBkxNi8
LWLLOvEz15r+bD736WvT0CwZidiO67kd+UvRyMXdcBQUxcxVPqZON70rv5kHGr1p
8b+PzxroboQsdWzYCr5UmUCkIYYaGuSVCxUD9y1Lym23qk8UyCvPPsDrOQbUpUaX
BpL6HCpv7wYdyn4+D/k/ponkUAMBET2CFAB8MSzRTaHTLhenjTU767sOFiTu9X9L
a3lndZHE5b2pLIx95WVXHPo5ch1HCJOWo7YYkAkYzsxOx1EOtLvDn1MoGXBe7XRS
68KU0hLMuxI8VsLnOwh475BtbkZKwPo6/tacyqUj53AM0Jat1AMriCe1rDvYbbIx
f5OPvHzM3sn+xcEk2RxhV8G9ZnOwoa1imVXVP3dNr9d1kio1NpFAmG8UAmWnp/ln
C2iZhEurlHxOtAUrrKc6bG0aLfOnvn60HxlPPmhd+/r1htXELLifNREeWweMeGTz
UPxVM5TO+LinFWCpHj53oSuUNL0vuaVZ5uyCzV9us5CKCZsIUHuyR3zPbujiuQI7
yswEkhl9Z5Gds9xzWiRg4nVyENKAA851h4+O+S09DgVbDX6sgp5y7cxffgDbN58n
Z4+riM093P9cRG15R8bHFP7XzWBkZq03BYMfgnfz01KK+59UU08ZGmNO8uNixw6o
wTWlCLS7ecjtO+A5unMDo7Lv36VDHbFUl3BlwmWCRV49rju6jhw7pgNO/z/Zrx57
xOpUBs23tmgZ2qU2vJJjnMWVUTdIW4yzreLHQSw2ompWVQlNEXh3ntr9nKf+4FPX
XzfF59zdAcJwKzu5iWeUEseE9+Ejw6f8ADl1FRoYrwTHqQyRSpc9/EbgfKDSJQ1c
uqTmLtosmWVfX/0WXInGxdPtlpZJ7ZDFV8WzU1ec5yBZMXUe8THOrTnygNX91eQo
8ww+Sx9bC+uF+qwEgDPuk6D5IiM3PdwXJ3g4oaejKu6zTLT0T8czNY8ZVOBp5D4a
5oLibpI/Yos/PgqcGOVFT4rOkbEGg/NaPl1zwhX6Slrx2KzY8Z5v27uqxl49OJHp
IJUXzqmOWqq0qAjvWajVdBh2IyNxfXrN3BqcHZrkQVz9c0/2o5Y3syTtxsLBv5Hv
wX5EwjTYiIPYCDz7w4na0rB3xQcDg14fpl+Yv0fV6MVqWeYjBZcQHperQR70ZvNl
763h1lUv0zQrfjthMTaLZqTtmJ4ERDkZ6CzZtzEs6iIlDeGrlNTUwzI5xfkexRzm
o5gjCsj/vvIukBaLsYG/Q+47vm5NDN8Z+r+FFiQdqgs26LzJXjKKF8htLh86TDv6
JztYbKHlt4t0EVV6GMd3Yyo4QiZPz2OIzUWxMu7igBBisg0V6qtQhh/ufd6g+4bW
Qf1tm1aBd0Is5J8TkgnbnHXdRnmL88KEywVeSsZ2ibtayzZFZhNq/3vY8Yvg9kIc
xRTGlhS6sNadPDw85Tqgbr7lqKzsfEd/2vuviNU2aBbXr/Knn1/KrI7ndR7hrh1B
Jg9bEBa7vS689AqpYGYsjcw3vWOaiU6Kf4Q042Io0bqUgKxgS/OVrv0k5f5VSc3T
qc1Vohx1GFBxasBUyw46Q7a9/MYLN7mQUGp3bKZF2DbbUzhxMeMM8NT/KR6g+FV9
VRTe/SUHWgut/IgGAZ7vJExLcL0mDr05OH79UOIG/GLh0qQZnd6oZOc2tPqaOkXs
PZO7JoSa8OpgwWHiChXKffOHJvPebJqkYUqnGhh+ikzNvJgvjUgEAMCAoxPgdacj
UxkyQymDN6PgCrWjwSEh1vsobYdmBu0M+q+fUUfZRaEsgwpiqPmgyrESMrk5cD0p
JojnhH2FerL5HfxoEZbejrlDJvNNKNdFb53Y8pOMaxiBz4bwRkx+Wk3FmAXNJ8JK
/1CHd8umHHKjoscOz+fhGelopc9NRVK9LB6MRmrOoqobeEyZWH7tNy/id/UNUy7U
8VG2bopJY9p2TdfdT1piuRpwQ9sm2Eguv/6NitobgsjJmMEmxUuT07AjVDAv74Ml
VW3jrcUz1DrQ/TRaKcR8f8g4Pi/o8//RMaD+BtoRl5h7G382wdg79YgI5qHFNKRe
tdlpnu5wM9ri0cHM++v8KTGIztJyieLm8QVnHbXUU43yJ20URqwWt0ukjhWKvswp
w4BsWtt5gzG87mY0xYB4Zs09eaWRx3MoeF9VqKrYbezBKDsuaKUtVTjMcAkU1MTE
Ptkpw1hgQXkA0e4hevOt62OvVrZBoipqRpNLRdvkLu5s5W3FcKwRZ9PCQp5dao8U
ePn6Sb6I/P005Kx6wgArJ9MJiqDRqZPeQOApmgfPxcBwWtIxl+18zZHyzihNrfvc
Q9Rko+EtSzbuaeE6BEUsyG4KzQeXAZJl1ACwPyVlpEtFL/Mg9lhBY08iIwXyssrj
y0dJNr0c+M2okOOhzx9/+sibhd3PGI5LMtKTl8+iKb4R8u7yCDKgrVmsaK70lB2O
c0VakoJhZsMCpowXgeEdnKeOT0zuGngP39YCzp6oTCZLPfnfMlt6puCLKPHWoGqX
+Tb794tq8b44wt0ShkpFWDNcjVPb/Gq52BzMzERWtXjRZh1CTLKvXWNfx3yJSNUT
pCACHdJ4kn4slIey37/L62ixIfRIdq/vVYEAcC99bykrZUH3FB7sGyZoZxTseEq9
h8RevtzmkxgUJx/jYlM3b2qi4NcjSXHQngqwcABKrMe/KvrrtOSar8t3iyWpoq6O
0tsfnwCt8TVPk47zfucyLfjjJteSCZ0CxYTsbJo81Ph0BwdCnlRbnYdShQyag8LE
MHjrfYsvUZg3KFzMAxAGTOQv38doX36mXMQrhVxIshWjd1GnTk11AvMxWZIjEDrw
Z7vo4SUCcxCIQPkkO4ADE1JyNWD6208OmJEWpUzM4aBuHxkjep+8pXK7feVMcRjy
wu+N+dtVxeDlFmmc4JQor6H0VosCUzjIVIxvnXfEJoJHyLhWvXp6PFGEdQ3e9SI7
8v553p3msdVJ9VUyCNUKqm9Eh0Ad/FfEtlx/1YfMsd+YLvryYkykD+pj9iZoMkpt
wlGG5JPa+rg3cWsX4HTj8hvsoPrWfbqheO6vs1WGr1gFiAsnu5g3CgnsK2c2LTsY
iZ/xOjRiKpwzcGWwcD7I5c47Op4OwpU6tHbKBnF4nLknOf0ENW+k1izP7wE2EBI2
m0NBGTzzJ/Pub4FXz0PP03dOPcDZq8346/85YorT5uLlEzxkMmYhhP9fQY6EfMny
uynO5cgZmyiwaaMp1kEuaiGekuTfH9/5EWKkR5zwVTr0uE2Mzg/i5BkdIbxtAVu6
hxxUzDDw/hrucOoGvfd8qs1I/mbVMycz5PqeowMIEDl9BTfZ/HCMBKP3o10d2PLg
R+ZHaubE35rtV6cznkZbYRC+/t9pwb41awODZkrsbbB8nQAzswiI9V+/T0JDCVJY
p4Ob3Kw5iJM1MMe0N+Ay/CCwHeT8Vg5UYVxoPOAJak2XZJiwukQPsASDDqNShYfJ
m2Qzew5D7uS6m9I1Y0hgSdthzJEEMSGFU59D4knhUabfa6VBR44o2bo1k4KTlPCb
9MYGQEg+0P1Ae4dECSfvQze7z3HULbDVx2ZpgLdIheI5jM0YnZ5eMh7BD2KTpnf4
LSJhyC7CT21xsGel6on8bBh2rOeX5uw24lWvgsh86va0b3fgwNWrwZTLAAZc72l0
IbAyHkwSiJxB2ZPcwPoLNysP2OIVrKi0s6Aj+5FdRmm213By/2xfR4/C58GGJ0Vx
Bvu1+3+MPNSm5tsFEEp6toyGS9K+/Tge5kLGbhrfTsdyzCbYu+kk67JCpx/OD6ON
YEgIIqSvPoiCvng5vHjCr7EMc2ZRQwwDps1+qpKs5xDLUXS28nuVpNVB3MbjGMF7
kt222DXs6JLQ30BpYgF3NqnSbgdYVV6WtTzQ5ZEapXX/3dcuRbiqWkXHGW4YatSP
0jB1Yk0o9EhYQHAPSMur4SQ3rFP6rDCZUtbrd7D3OkHrwFxTgVznS6rBMZB3v8i2
4zLSeTJ0gRkaUyczo8tQalkF18cGO0wSQUMDJ0Pkbn+cJ4etUkiAHzQRFGtj0qfj
9LmCgfBP/x9EZo8dUeV/HcZgzpJXuSyh+QZWpGhq9eRV+hhkSbx4i/Kqb44etBCW
ABCECqhjfZfl3Ms9SedztsmlToDu5kvQNSAMaa8CQiya/R0xARnJ5bnnYcGKXLbb
UNXo79fZwz1hHe1djl/wbknAUr4rOfgs7qhkUEXMSrI0HtFMZZadi7DnvAaHM8zU
+Ze2cvQLUOjYKO7S71Bn8CafTorYGMaSFYBDhhEM9Za93UhFm3l3QOiCp/6uVD4L
SPb/u1YmFTJbcqjBC8+bShktff43es7ctVhT0UE9V+4QjX+QWLbMCzgf9POyoin9
cnK3BUgMOeEgbj+WgHaPKVbtvNKrNk0m6H6YHcVfAWIiX8oQXFdR8r85nuLlJFaI
4E0TOi2zQLjH9+/4PwFF94moH5KTVcnUszuUah3nu/WYrDMusJ4xlZwSApcaYhya
Ll45lKOuCoW5grxcjdRU8++2sHbI7OT6OMT1Gry0X6FL57/qXYktArq+lPUbOxxu
eVFRcg+5oznOObRhlA4VykwsYX8+fJWFiEvMiG8Yexu3DoqzXSjVbaLVU5ZcVTMO
0t/qjrjnAp+1Ld5qNbmkF2duPEbrtOy3FOqk1ApEkv1q0nCJEn8/M/g9RUQZaUej
vsZo5lE5WxQSVLByjrXpu9u6b6sqd1crjiHabXpMPiWsZJ4Y6oGCDSVpK8dyh6T1
VAPnU42r40muminvVwZT9orCrhhLWvJW2gKx1F3DcsDeAjl8wA1ZzPQdPsJrRmzZ
mQAXVlKI/w5QNeFOwNrXgRKziFJd+bifEer1WD8rDkbNYOGwSRAKRLkeWtVM51gC
iw1sqU6dQ9iP/hvUHJ16DDRnqB9qAHpXLt4XCdIGtNUhrWdz5QK4w5Emaj5pkx6a
U9d6UhGiPrEl5DS07a4TmgAxaXDfMoI1D+X/uNVes7mGbh3V67FZYeH1sUS5NSR2
YrNoMpZkTIjkEsfmaxRBxquO2PubzIeFPzYEn1oylzzbL2kl77/Mz/pmWuKuHV3f
mjfpqLpjcqXoT5Qy3TgG5GOs/cVMT67gss1pJHdS1vU7BdJov74/pxPD4TYbjO4/
0N6PA9d2hmiuVzj+XTNEyJGG7ynmIpUn7mYPq13uLEnVRtgv4HSeEsZwfuS2rmAc
exVl5m4HRIBGZ+uEWEMfXiRonuFaprCDMJZMWNBvZoC3hvDX97xSuA+nC3q/Ms5a
MAqeEueobJNtu2W0zzb0a2z+DOnlACcp9uwaHNhIasg9rpyhYSqTIMqBiu46q4AL
htSFM/j8R/uOazV2yNWQPlkEYiHE6DGSknrguNVRyNu7t5lZfqo++XBkj4SaiF6N
zZ7WNu3XiDF6y+iGAII68P4he39IwBVrrnMtNZDoCMUyXgRtUELyLp04XrccN7IS
6a3E1Nje3xj3a/2XeArJrPUMvHTwXJFYp4nfHusI84k4+OGvQvXtVQjjc3lextzs
jh1Yh25UAHKodQL8CRGxr7uQkSGFz7/zvDDPNqLT+/TKXISzgh0TgMi0HYg/aSEj
6qMV4AqsSBoez/WjwdKKOewBLq+Rpn734ISQrM41rf/zfPKEHnG9hb8CkzErkPuS
slssLdT7UmOiZzL1cGkaF3h+LWm4B6KxT23B+KNOGp/guPXiX4eGs2guFTCXOASR
OuaB1NuYQ3JxeckCb3N+FlUdxgJHxodV/0UvZryCkrev4qTdoYuI6fVmH+Z+bQGM
wM6p07F6r6ypICQ4+VHLliGkT/7lTpHRz7nz9IY05nPzC7piu3ZSNJyXuNQhk/bx
sQShtbSR1IoLmcTH/CnRr7QzRVr1382eiYomoN8h+gugGQuRElH2OKLN/ga2FHbJ
4bBiTdhI3driUIDWz32x+RLaXNDKSqdWfpWAK2nS8D5eBvDlylmBPCm+qZTrJSv1
JIX3i1uBEUL+zEupUbxePAo5U/HKQr3lagXenM/GdBVE16VQELa1gA95gkZ1MhuQ
eyPh4QkRPKNhPRyNliUvOY9AN+xwG+TfyiaOVOPOJW+nC/ogjIdZqDj99wOPJgfq
1bum6cOVBlSd9PXWUofJNSNPYctwZ5SIJENfzpyqvsME1iU/Pj8wDKOcgprg3xxL
bsn75Ia70VsZxp2aaxaUsAxy/plQiQzTE3D/ERoJxepm78UqzSHWbMNM8oA9Jk+3
fDU1oCDCWGqX/YVxDX5xic3QHEWHQHnuvzWso445O5MOvglzZeh/Vn8OSHFwk3rD
Qxb2P+Um3k3uRX0qNJ4QcJJlDQ6tkUiNpVItpjo4yFCwBytYLQzgXYiCXNmlf1Rs
OXQhIbpyB7pS2eK1+BGyUZtkvafjMnBd0T8F25J0XfqefvVF2+uqp+cc+YMP6L+s
JMXx48vJhoo+cLD4sgPXxvB9TAamvu1XnNqC/nEAkISomP0h6trK99DV3cPyvXu3
l3ws5apJSy1mygcoBV4H6WO8qUYgjnewCtcuY3V3VtLoDDiITmrxcKEE34LoGfsR
uVLiJWr9KNNx+tzgAan2gq/Nl36pv/ggLO7CqP0TJWXTeVBEUunJT6y7uSvCQZZv
44Kal/t1ig9yfAuNwITtpdnBwZQrG0PXaaoRyBYXiiuw0lM9Anj/SC+oKKE4h7L0
2aVdDIBfM4m5CNByDc7CdAS6dAwxbrTocMZEWlvJ95Kw9a7as6fN9Qx+Sr9OP7X5
mhpGK3mqIIsuyLGgxkZDsiZdxCBWefoI4jwpSxCZJyPQNEoocCeex3SyrScctNTr
NT7KCxdb8HQiZbNXEilgrZ6YS7Z+K5c8wGpRJ/7uHuBdfIApuXytt2YJkEJIj9cB
AYhciH5rZXr0c8wggpe4CrgTKc9GSXO5CrqB8aaS2pYDLHP2Wwu5J/XdhgnlGeVc
jTIw2t1vT2OD+l2aUf700DTRqeaCfKVlsSAff81Ozf6nA+unUsPrtwe1Ppnw61ns
MnNYQiUR872o8Bc7wHvTmnss8xg7GuWbU0Z5g3KMc4e2EG4hGIi5S5yTj51DFReF
qhaGCjqTdcmJSCbedmxBbuAUvjzhIqRUte1TzLjJuXnGSei7Gh8qGyJf8k8t9IE6
20cRYOoTMsD2TE2NTaT1MTA1u6AYrMKAJfzJ2F5fyjjMkFlkuOIgR1uRUrY8tUii
6GlszwdpR2XPU1nEvKpnJ2kATSMXf4tTL/H5OiNuyUTze+70+PzV0SfcKI2Ofo7A
wrhtdpxQ66G8sR240IDCeoBGgZQEqkQwalVK6qENxhaKAqQvZfh4D+Vgv/jXjtS6
aIXXB/FbAbjY9koKGYGORlS8RQ3LvNppIcheD2FUuaovw4RL0uJqOMBknWsepdqb
CI8CurB3FT18daBvYRNG9Ly9FeW7kPcza+2zrsfK1saoBIukqiDkoWFhYvZoNtsD
CuDiGf/9ifqUZBxCdE94O+M953plWJ1iDlMiDuaFTEdcAX1qJ0f8BvEudTsbbSGm
c2HfnMuZTHSaaw0QEb4jnWFiyzNnSIsOag0XtOrdvzi/AHb12GeQ6RmK07qYUWVN
rYvwW2C3JQ4XO5cwY4cCQApsbPyCpSwLvxDHS+8mxZ2dpMZ4WDLLqrY11OmjtXLA
TBug3hkYF7roRLH7HwDf8mgVBfSm+GNulR/Kxv0S4hq2RPz5Ulbay/dF071fL/KP
YaDsPzjshvoEahESjbz0C58GfPdOA7WlDgQ9atdROytNavDqu9E+K4SYEOsOuXiU
7jwkTxdl/De1Be/vtUpl3zOjNzlSSyoT4+9GbRbP6xIXbtLaL7nIa+HWtd3UtqnY
ig/hbqbxkgEN61bjCa1FJ9V5MnIU2NHVxL0q2eqd7TvpEq2H7xHGDMv+n+b1xRrl
wbwm4yT5B4eYWHXq2yqen+KtRIQ9qii/XP6640U47Sjv5UxhNKnqtXrA0nkTQW5R
swTsKcjvwDf8wW2l/hKdrWfbXGy5CtoCfBl5bZm9W/1nafzEsadp4uGwbK3MXD2Q
nB5c8S95F7+Fpp6kkktCwpzjm2uxpFPgV7llMOz7bq6i0FcY+z0/PUSX7OR9G9si
4Hf6RifD1BVA+YUvTVKUYD3LjaRRw+h5kCln5r8+Dk+thao8mmmVq667a7GMd1yF
/wXjICKrURcS26QulbUXCGTWpKO4pEZtugZyUMLsiNdyImkbe96gs9tA2AwMK2T0
TgPQFwd8M2ohINNQSruImHuYb53FdQ+26HEAAnUC+CEI2l88MNqV7xfo1P8X+QT1
Qy5VE2Q1PQn73/y5Hx3KmUG34KUAzc8PvueRIwxqOSDFf+xv9VloEqVe3Sd8ICRe
qowh5y/uoDkd0+kAlpGrvgmU0vF2mKihmaoReeDQRfId4mQmJPkgf+jYYpfn9GOP
qY6EcOwLzynk3Pp3ZPdJvoKz5jkXoB4hZOlPiEvNIB8yPTr3+4ew8nD/KwHA8iGa
0BOjQnIO3gXMumd5NQfixSfIaeKcV05PKXvCfVrSxIqU+3qhh7Lgv2ZtYG+UtUQy
Kn1Kie/5pEqGh2M5Kw5h5t16Qa0jCFFj5FSJq2HZuLunlzym/CpsTd2cu8C68oTo
QTzRy2Q6M79Ngay4v3eQaUJ0xttOXlxi7dnxCEkCbiZT9Bag03Rpr6e6WS3qUqba
njVpECyW05pCIcoKu+tzFCXqnbs9dLVFzJZSMeMj2XCIPraYQNManPwVn+vq1I19
Xx/r6HUioK7YAUmFRpsrwZ6WUS6mR+M9qdiMFqbmjCLO3X3Jb7e1FuV7hhkrF6dg
z2XnoXzFAm+rmKOmuBiT5s8HMxKqKJCx1wMZW6x93oOkAUVtQD/MWGObOTlzVPyg
TcA95qp8msCf8mbRLJ07TGFreMYk5bExkzn6oFKGMvng0mfNU95YSfAmoJNCmwPc
l9UN2/nRNIg8sGoUbE4/TBtH/pSDqedTpBjUY9S8pWpqWwdqvLSRosgiWHTXwUt/
uKYUKB0zsB5vAYT40HKkkTK9m7x1pQT4s/JMfKPu8Jds8jNSToq2PnE3Knd2s9oL
hkLnNAVoIMOVjMvMVR0eJ3HCE733niXHJjrGOGWh5kQ5wDrX761mOxBL5WyhzQIJ
+gKQ8g3z15nUgpGWjyDJrJC1udslOtDgWkW0wS/4mwo5i3BJPSznE22HgfuCHEw/
19Cl84nZesHzVYMoySKaLz1hn72zi40lWo+Z0UFcbIVGA9/j8jH5S3Abm64vpvLQ
A1Agi0BIM3vraSLjAV+K4uEe2C5uzcWTrg61aSwOpuyVPdXYMPW3oSJMMFofZxAt
XMbrrfB0YUNVxCXoUDd2mp7wVM7YWzugCEtRB/DZkVkX8nRNnAHHrV5UBPG/5UP7
aCauxGE/XBl4BhGOvhqVBezYQiqw55dq+P4pqjxakvkGcDWnn/7Ee1RTj741f75k
WvhIwI8+e+brMOv/sZGhDPisB2tUo0XwyURRqeRF1pag8mgO+Oi0Z8tbf/XdwbP5
qeZxIvA4ynmUpTvccM9WsQFJ1WLLaDqXp7CyJczLvi5+NkPns0Ut8NtAZp3EXejA
nXc23B3vhn0NLjKH8slBfE53+r5v5CVD70emsRNQntrU14W3LXeqDyI883bKwXFK
/Z/OBGzBLtF+ljdAmAgLAPFvitUT5E4+m1tbHGq98chuTpe6ieOKH9hjNhhIFGUG
IpgF4Y06bhKUC29SlZx1uPwHcakgYWgx60iJnXve5MidOiYtCI6kJBxHU8Gn8dzW
wMcbasndMwgwCYNCbCVw5S1LtY8ny+qtnjbm+BhtvU5h6l+VEv5sx1H3ASKwd9Yc
DW1Hv9Gpm4kOLFR8YyotBwJn13kXRW2qxqgJZBRA0rXD0vz92Vv/WOmlQ3HiHUoR
i8VJbztBOJgKh12RQ1Sn2Um6g7WB65vFxXl7SWUhQUoO3eKQ18DGdl68DBi8bd1N
IVYBSWK6EOVieUlz2+oie+2MRhHgT7VzFHVsGN6botE9MbSSgJHwh4TqZw88yNEg
Oy5z0idK9po7x3CIqVZNBuW/HkHuG3W1vNe/isoP1yXuFWRTLF6ZcQU1SDLVAtNJ
N1LpzYRljxuR38xR9t3iRGEjvppv6+QapatyNSxNWERukkrXw4WvOAJHkBVm5mif
OnmSFdqEur9N6+Yq+lvtoIQwTRivJbuRxT7EqcFkAc6GUpDg9eJs0KRqAjwsyFw6
QoLCJ2aMlxpxC8tqzfj/h+fC7S34/oDg8E+oX8I29lK4+v9sh4LxU7w4nK9mEpye
d4gQTDFQck8pImIygQYFwpfQTLaw3KrFI3NMa7E/rw1B7Xo0fyeleJ83Aue5tU0a
HnLY/ilwaFPCnXh6r7XFULVsSBprKsHZljbk9uoAXcXhMS4WLqzCkFl5e7RXAO1I
JccIm8tsTPfatczBjpgTXvfTV+VaU+liV06JEMaO3puNywIvfWKGZZUbRpqoR5Pj
uFs5mFNg4a2AbyVfHWP3MRMkab4KKJz9t0SvQNXKnFUoOcm+j168Cw2G+JRxXdxQ
LGieCkY97uVzu64rQes73oYAmYN8mhQrRjam0tfi0KM14EaCioAAkAOXPMsilwx7
ogFMbY9KYl8XJYTJLgqF9vk0MYAgbV6ztYMCmmXbh2wtVoIi0jrtCKsyKIECxuhk
wq/oo3radieo52blWmvXLJFd2cbneyW5UtZr2K5KYANOg/9miXTvKII3oLJj1DJx
B4TrC4nwx1jBDJ2KMp8CqyojQI+LipKqNwwnNP+cOeS7iEKhm/4oqIWJbSS5xsbH
u8JDU1T+5RQ/cepd+Gn/pBxe/CediXBadRL5IaXeoZwigOw7x24UF+l55wBvG2G0
HWfmHA62FR7rcCzF4yGC2EdrtvCYpebSJEdVD19lUM4TP/9f9DLTHMmcsohLrMy8
44RDtDRmlg6RmkC49DPieD3Q7rudhLT3AqtuU/Ad9VDT6edgoPtnl7jlXZ8d2UpS
EdfrWDmw7UmRtX8gcWgXiDnf1b9ZZbR/DaLumpX00odPrN5bBBV3VVHKwnnrD9/e
J20mRu03sfPBIUDxJzqhLDfycgMml8AXKq6FKKHkNzLD8uNXU4865/Z0qlrRSdya
sXDzP2+GxVww5y/znHP0gW/V+1Q0jQvTmxQThNzMUgkWfuL8cMVB0sIAZWIWOlYd
/4MKKHZqecczK5ThTfhbCtcVxXoupqyjwym6QNzIm5xX9LDDoKcCHscPaj4P7W28
Qc4ZoralDKMiYCN+K1SGtUmA7tjrxP1z5z7HHrp5nWvQqWXIgpiQD+Amid4qDWqq
NuPmOsrxfGse73Etfux7Re8Mjcoen7ojE6xZMs/RYEYuN/kdKLUAu3S6FEPdXeEp
dmQExOzaIi5UR9Ahq64cvzDY1roFu5Lc5uoWHJtuvwOKikV2cPySG+ozpH4aVjrh
uFBvH6fMe2QLFt9rsaw/VzAg9A6y0IfaJmsZ3r3McSC90uxngX9pEsIEUwiQ3/PJ
JUw8KPgFTp3z8r7Df8dulr0z3cGyht3mvo5cyjnP30OPJPTigSWq72PBffkAsuv3
Rm7tpvcYciUGPGreKwQH+cmwl7gaYIw+QPZjm2dMrbku3Y/Nij8Nqy8p0a7iG8au
esCSDiUs//W6FZ229QhXeGbUReM0CnVCKtP1MBkd3BK7fG/rajgpaZgxgzkretWb
NFl850hnfy6yeAodRAl6P9ZBiLdrD387vAUEx5sKdLyqz7YYswKEwBNk32+Qyj2E
0aXIaZm0o/OOJyIlaSguoIPfEGCJD8F1TptAHpoZoKYaMQRmgaz4stBy/4bx1Ex9
xDnscYD1dhO/LfemlzoCNycsUi4juLyKMRqa49BTP70eqhmDFD5x+ERe91pHYEGe
RUZzMrLl3R8xlThN1kH3yiEPk+qTkEcMBBKaeaongPTuMsg+9oP9iF7GK3h4Ch3r
EvnzKGEFGLm9eZRkRb4gKLXtuydfdxb8jJHvExNlF+mVtUEJ0Yb22YWpeLqFdA+a
2RH5AwVYE9ZArL4yQuoYZxtdxBELQyAUGImGkvwsBeCMM7ujRcElPr67Bb/Ieesz
tYHRRytZtmc4MI8J49t8uOirMgibVIY7jsrx1kmLDdytR0fZEk6CDK0q5MTHJM0r
QNRHKhLYdKZSpCCD7x/FcxNm/uRBJ+t7cymiJ1lAUEXhR2ACq+vYA0A9Za7lcblV
5MqyCsu3jS9147Sb9x1b7Qa/hoHmEDTbMdDNu/vZMEpg5/mVTwhA+kpFw2cDRN4M
tZWbpa37eR5UJy9/NP9fO8K0In1dwEwWnXV9auGS6OpEMooA0U1EKKviaIa23TDi
WqYaLRjK/KvAongsfUJjZgUbJtk+GT0w6O1H7KNsRsCcPAxp4Z/TPO9Rd1KuSIC0
Q4bXTbKM+jWeDWBNChfQSPyt//3EUyEL1Gj0qBl2lDRLppLRZDd14FBAyrh/cQ43
2f6OiInE/a7aX8FTTWjSfX5u1S8+70i1HDZNAFtSnT6ctjh89B7XoPkTworjDLvZ
uPGQ7UhfVQrtMVUmQnWccmpPjQjIEiiAPKaU5WfWRvWDtC7SQyFTQ6KYxc7td4SM
2ZqKpuxF2Qh42+x1K3I/+1gG647kY9CpYGoV8BCx71zBjnvZvDuOWy+Gs/1dwETR
DtHBO7nQTjvA/TxSNQV1tiCfIUJov20DSnyECx22l1nIQaTutknTwbZ0P0bVOyA3
2id55NLtuH65tB6qNSbiAJf1SWhl8dXd4YgvTmgKyxXjbuOcqnJY0drPwX4vcGxZ
Yi+9Y4ZZ3nnz0feBMWoVQiaOcmG57TilxRM8mw5khKNgrlV++5OGNZGv5dgFH0gi
eBtxjxS7EmYmTTdMaEEvdUOVPM68dQFcpa2w7/vPoT++Ab0T6W4bfa0dSUB6N6WW
OzrWi6+fow+GTqcDx1fLt6anGVHwDhbxbMv2es6ghKRS1XIb2ZNUaF8hMdlaZL8o
qTXwERvuiXf35Wm+et64WICJ0FgPKlsAEQWg6tVQor+fC/uT+ZTSV+aUZLR6wzYy
NjSEvMf5ctUALtqPxsg9/xT0pgQGmZE4QNYdOupjwIiiUstjnPKSvrBs6dQb7lvE
a+5MifXRLbJ+zby+4aVv4EI6MdyTik3PnCKLAY8XMYfz2rRsnzqJ2gxMnt8kUFjB
o8p+BIXpXbDFjq8UjG64+MeHit9F54GkoxuyRwBhKdYh2z65tRgSb0Pt8260Uis2
Pg0qETHnMIUmRnPtjdgLq4QzzZcDMEIPPz3uWaCYtnolEXFcd5Yf9/JWGJ7shcm3
mKwZJeT55YHgJw+DPbPSPoi0CKws8sbILILR63lLRq9rjUojDodRiydgT2t8PApC
Vl2N+3Hwh8JxZRZiLNPKaAeKZG7x6dtPSiF2wP96X2+9KNza2gcYxleG4Z5Hyrrm
AWYOlvJFi3QhO4361nylVQAfK1ysFDWUwQrqqGMWczImMeYYMwFMQ0cLnLaTw43q
P+DbbEvjacaHLDaOaiouOdJFBNntdK3+8icKCsb8ZcBQ894fbcu4/WGGRgKrsWSH
+dJ1En6PJ1jzQCpWTuwM0w+67TVTNhf02+zTn2iY7p1MbvQMX9+3oXge9VzyddpI
MSvtPRbYJ38cpd1zmm/3W7BhB/cfT3fVOL4YdgzH2MZw6qel7/yAMZCqtQji9UOS
UHn7zXGNIW/NaOv2mqb+qV+h4uUIhneg5AFkfE2U/Q7we/0hHKMbv1sDr2dr/98K
3WQ9w84D9x7l3DCaf/Sn3+Kqpxe/MFw3sN9M1WnMAuK4n5r9AOAgfw+qHCSKtxLR
lrrgy9Wv7G6dVMkXaq1elBNgJ3nk1DyLSOC8liBiNrhM8s1Y6g6SVsP9gp3vFZ99
wfUNPKg/7jBOQ+fWfPUJO3OgZBWlO7ff6hl8MoU9gbwM0mdkPpAP/49gvsWML+4g
ZC8g4SWtT1TguVieEMX8CIMCS5i4AIVB1wEWwg4VErIers1X+g9civqQy89OzWCz
tsBk6KmgsFdBA4YUA6KSnWr+iQ6D/ZAEK4/CfWjRFGQ4+5o7YaJVj1RpWE9EfD5p
JYFmUMhRTlSKoLlji1xjubjeFDe4fEBdn77yZ2ldF1DVoS98m1uI/TF95ZK9FjC5
o63UWIUYm/nooU+himWh/bp3UxXS7R2PYtq9ZZV8+ygik8I19MSSeJyIGdOTcf1L
VhdMZAU+GFKnR7ZFrXbqP7tEtMdTVm6hR4Bro9lMRIN6pmD/Emq3d7wYEI5hDxfD
l9yGuJuNKw/zbUzDG9dUw7kRo6olKKwKDdVQLsWFPz7uCpNYM6z7Ke9Jumqp1F1/
lLG9X8iiRVQosR5NW2BHYIa03KT7sjQMNdJSSmsRRJVZ7a6aQ6sGUqe4OGz6iFW0
XoHuavfoL7XUg1JIsFDPpIdIQeGo/fI5Guhix6+10BEKZ/LMIRDAn8XJs+eQcDix
ZuifvWbG57JpOheyXU0ay2biZLNzKEMTAhsj2ix/3PSxkXcGdmDpulKNjkT5GU7n
UxI9U33PS+xVwda32T4Wa6QIjKmOXb3neUyyKc/iNlRJhtzLtudkyNpk/xABZa8C
ox6jBUpj5PNOmhyvlCnr4jRloaEeBK6f1lDiSZ1/DT7c8p2TeHWttA9uwQ4dhP42
s5OAOm9ipB7ZORYDqkRt/jSfmqmQHNYNKGivmabi/IaBUNxhf0Fca89Zo0mLhFXK
8MP0hsCC2JC1RvXzc7fR9Qfo8VjZD6vq/+zrh3F+q9Buwu6cCh1+RxKrPaY3UEM2
/Q1W5hBqZAxA30anpBBNhxKuzPK4YLXHtBsfzNXDVHk6e2ccMjk8JnsjXcwdIdr8
J0+5uH92Ns/tL7/iTvrMgYgt6ws5sB16Y4DWAgFgTOVifxOwrt/NbnclYnwk2dep
mCISKx/HaeCLoI8Wm/1fvujeMsXpl7hgC8eft5VulwHlfLApfRcb90Owc5d1i+cg
vGk60PXZwoeBVZiHxd99LqQVQmHHHXLKsdMl50qErrMse6+jpupuaZxHXH87GLjj
ldyKSaHP+9WXbBI8iI3px5J3GamZLX6GTFI+vCHaCsa4Ya15ZauGB1Jk6DMJSIjA
AFs4pnQDoA/7JgHsO2zSwwGzMXGgYpJ0AxyWr+s5KOeuTwJ3R3eSdQAccQMktvqW
UEbmAN6nadLtqffU/auzzYa9CJKPRwMbmYHlmqJCP58i7vqwEFHpYAJfI0SIIQnU
+aRBmdzL57F+p9a/rFxe/WfVpSrDnbHWxTwwRwEBDrJzpOEYywJf29Vpm+wz5v/G
MqvwN/9Ldbl1qQ9Zmi9Gytg3AcWl2iQhc6dvROpbd7J7+2FO++LDvJFyoLbDBSgU
kZsMWeKEb4zj72EvZc3QqZ96VZsu5iPylN2RzETQAr6bdYGpUE/756Ow6xs8+7jv
KCFU/E2omDnAQMZRAQBFg5gJAhB9wVnnajEAneHFg/c3VEaM7vleqUH5vzyXiRsp
8zdJygPF2l9nnY9jeouxf1lUr4r+0c7DwcONCysWxJs+HmNOBaJEGGqkblF0KiRl
MsbMxDGo+S3NuvdcixhiO7P06bCu2srnO9AoNHY8XsvJMdyAjnF2R7lN00sGKshV
DjxTt1FWecfaQeU3H+V6AXvLqpx8YPUKNeS6xaz0ahn0ApULQqdEr72hrq+1Ippc
L0Kadrv4ucjzXpXZ30ZkZTzq2wi59Gs2/qkjJzUNhi2L3IYeoP++iIhkfTB+0rRe
MKMsKtee9TrxXb4nnFaxqSfv6cvyxJeHTtde3O7qrSB/lRb6QT2Kz2Ik4cbpzP4b
Ww778934goA4c9exARtVAztQEfImTsyvLN5w9Tpm6v2RrbCOPrVZEfIjf4dKLpLK
0QmWoxqY4qgd00j9D2zLTJi8sQOA0ndU6L7pKvzyOIgVitidhMbegxLQcx6nAp8m
hkv+q3qG+TyM5T4a4bOYMbxt9hmDrNKyCa7x2WDQOrMr6+wrAqV6JLbEoIqLTcAu
wnofdRPrFzNdtdF3phiEh42uFgqM5/pSN6is/myGfecInyaVaxDOxrAL5Y+KQjXe
jVG/c6B5xzjwJS+1OY36x5zchPP0edLh5SjAl1gowIBFiEfHcI1HNaFYOr4XfxMw
wQACOke0p3rd4ItckqVWwohaYrGSmXvDwH6XX1+JojUPY8S2oUeTgFdA5BC6eWjT
z/9jemviJbEyBxBTF4WGWcqVJmCa62kIV2JKDdCX+EJeN3TBPV6mHoGTK61BuoxF
tJzLnX8ROQNHxF/30OKx27U0NOaevilkDJks6Ovu4zDsN+YuY9QXhqzjzX53UtMT
xCXOAl5za5kc+8SIltJsYGf/RQ+IMSuoyari0IlbVpFHzoJcn++8MqdsbkTIe7hf
5jmC4IW39l9tRyhx3oVfgxaf44EXOWdmysIZHVd3NQTMxnPpRdfqJhNcLx70kTez
ot6hvXDlDslpeMjZibKBuzz6ItVKxIRr7smf4tZCkdp8yPEtzEN3UQ8SgDLCxbWu
+Ezu/2f480VVb4JOlwX/pEMV7bZtqP87N4TCuLG+4LiY+7zhdxvtRHSHktTyBHJD
fCZjYzTkmue037dkB8OjqwhnaREU5K2QwwhGQDtlfVodQesRmOOORUcriblopMBQ
EcN6LRgdni1Z1AUNnzzDanI4kGtvuMgscldBY3D3xuAZF9Q01WBw5W66h0kT2GVO
IBdzGVV5tsFdIhz0QlfFfqesjtrZr4t1I3OR0VONxDgJ0+D7padhAAljXEMy7CxF
V9+o/fXmUPVsM5rS6hYbnEt7cfkLW7NOq4KiPcHpfkxFNaZAv5BoTCSoBLCteBZb
zSD+qU/TvjhjzujsL9EkL49q/Mr+SzCtb5LRiS1UzdlkcKePka+3iC+4FabBFtV8
kDLnQX1Kmm16wL0Ruzoy8E1bvB9+hGYgVvwxYUW4m8LUC+GRiA8x8yYqbW2x6Tb6
D1sLYlnLIKOKSXhYRf3olZlHCSKDACv/VtIbnsE5PuA36lqzxqr0KzqjkhQrB4+E
2p50Iu9w9qcr3Nn0CQbsSzVYGWDcxuhqBnWz4/AKvlkE5mdPLEn/LfCXlTWzia/6
CkiuDIf0jUt3LlRvX2rr86sXFrG1/7U4GWO2PxjDJ5ePBJLT0+Ojuid0+jx1HnSF
BiCwqZ+ZaL7GxCuRvsyc0Ha9V+83NH/qWgsCviIq/0OIKnCAViK3EgdosreiqjQZ
t8acFNQeqA3uksSmQAY6D6LlBFsbc5ZqUGWlS16VMcEq9qb4pKsDZeXn4G0caTHE
ThHVKAkDjZ33tkRlaKCUqFQ6u0PoNiMbWRPhH24yNVoAeA1+w4DvU4r6QIsP/dT1
pHiYi7Zg9eNmZAQDNrEGZl2eVoQVHyIF/elGictiIrZHPRmv7Vo1uAqRFYnAJHFc
bIgjjR41yTHKSUpdoJXuL+m8zgoaA+t5JwU/wm5OMJDJWYaGx5Ib/R63kVfgTSM0
wRwgiyPjJ+KasBytPXlZmRJu6sOtPAxTF0oxd+6HkjgID5SUi174Ucn9kRP6/93f
q6eBZn6AQnh1uCrzlDY6Z5u+dnQ11Ktrp/s6kyuOeMbXVCRt+DXyQA5pTcOcDanO
5aLf0QehO50p5aFFfm1pFkSTnJ+G1HhQWB95l5rTZ/0YTi4Le91jYfXCnXOQtbkj
ni+kcJELmk1IkikI74S9x3/5ota2b8Q2Lr1pMj3dxTvWsHIydouqbIENR+1KmT2Y
D6OvDu4d4HWmiX4upt8oRrUX3wI5901z0RH9PO1UaH6/F8yRqsnuxm2vLk3ahqZY
O9gjuXHjhfJEcvGtBlScm4CMelTnOGlBvjmiy5bIAtb+bNrWrQ49se72WOFKKZBl
3JF1SouVLnZT6/LZFcLglf9vuhp7Y3k5wi0sL4pqQfPqaFD2mj5orlkkbBNaciXh
SXcvG1u8UzvIz1Qr+VUDnv5afQ1LTQYBL+OWqnZwXK5v5qF9azqMGHNFw1Eor7sI
Gxtn72hQHraqUTYangJVNmSqjhrMnFaE6NHhwT5eV0HifXhVBL8pyyz9FF9ZzWiW
N986G/aZNMw9IVV0gK1dt0LjSkHrzsuJkCy14WgmQl95s2EDmUak5smV/Kgqyhaf
nJkPY5dSYr2gA23CrzKzEA6GdWvf2aY9aAL0rvcOQ9nYU1g/hT9OMlp4QYWhKMav
dqRua7BNrBKmb67tHpbG/sxdfOI3CoCmw5409Ni/U5qGj1y7IPBp1uGbKxizCMFR
90Gk/rLiCw1hpP+pfmpIQ1nLuS3pVkZY/JJ7xLkn/5i8WhoG/9KvBzWjl53hEi+k
AT2D+O7agwfLI2SuC3xP06Ci3SNSoVFkddSaSBKTrtdkuxDRKRqwuNs/v7STCqkX
+bbx5RN+8dV6IBZZrBLlB8IWe350i8pWakiFxF52Soe5sMEY0m8dPkupvyMgFpCu
lIoviBDJAG0bB58qqba4ewtM4utOqPv1vKnhny+sTbiOJ+OoPvsYzabypqlB07P6
JtauH+qK6VRa20/DVO6gVeI1BRLGySvw5zhKYDpRyTeIZAAcd5ex8MudGwxh/gMK
2ZOVADYfpuHWRKl2/15g0cLnn9GJkEuZDgsbcRSQEFHR0pVbS1PQfxSho4nDUnGr
N5i3qhQzxvSLSyrpP8f5Y5YDaBwjiwyvD/E3Xx9aiNnj4MUiXEzza4MduSdevgmt
ZcdEj55qQMx6OZZO9pGyPMYPhvgRFnlZq8RxRvBPmB+9umoqL8S7XYnA8ZpAMp33
jLKbXYkRfuCFaXFVy2w5qFlXYoFTCZR+POpRPhmCCA7zfNrWw2Ebl0qk/EpU/B9v
C5voziVP7dVXZJe39y8Yren444mapm8SaWL4yaocVAW6QfvdWuqDbsOEJICkZx4L
O9eRPyqIGKa1kWAyitnFXTz1Bf80ZKp/R1aQ3BKVkLNJ6DrWBDIa1/2S1JZ0xoXb
6DR4B3IORdowmalXLl4lfkoWDxLtsn/l45ms7j2n+exthFCQNanv6dP+YalLyph4
thgOgkLTkuj9zZ7MJm8qxlL9ByqMUABsOGFPFto5Cb3+PttkOi/nMCAinWnLryC/
PmdN9WRkCOBlyRUXuR74IJYiTX/0G3dypr87MD7ujuFN2/webn6+DXiipCKYN8qp
T+iQjtQ86QlKI9oGy5eygzmOGud5jM4vTwXT36nNyniO2fjqfsAV/RKwY363pvUZ
XAr4pqo7wYHRlH2KHPv/FiLBWWohVSYesVejo+3hA6w5yAuLKn7ie2Y5hcNfxQ5L
+Jb6hHH2guOTOibHeQtpf8RMIyC69zvqw2hyTk4qyDI9EV69C4Cbmf3ZcS8Zeecj
kiwKHPvkvcJCA+tJAsYjrrqs2WkZOqt1cwJ7NN56O9uEif5XZwgHwOXIhWSHZY9I
m5CVyRZUR4RZy89/rsUh0UeskHVsBi6WiNEjCYcko13Mf/AxNSKg5djoNczTmnaf
KqE7xnHqbe1qkQ89Rs4hAbNIRxiuai8jbbYVOh0Zv/uh8ORFINmhWXRtZ60H4KDI
H3yEyczSy3CNZP1+mW8za7Hv3gqNHiBKoSXpEzlrsllt5eOhXRIkzhkUwIXGKj3r
fya/cGQ8pC/oGqGyC40yLqzbzFV8qv4nFYsPkDXTfcXHbkVkgsOeFYNh92Yy4syT
CZFs7w1pCexNMT7rN9+g4rB5ly0MdT04yi40lwfB+P7LKrrcPBmUhlv+XOd2hHKF
3MK+uy1XTUN8SbSAX/jtE8oo45jJqUYr28azfeobLGvyzKBaMzyT5Z6n/dztuARR
8UtoZ081DN7Yx+LTiaUHjubkSfu5UZNcOYeVN69rJ8uxi/Xyg5Sb06Enxc6VJeYa
zk83hdXI8k9ybSYhxVWqixW9Yk7lL39DMQvyqRskAJ37z2Oh4GkXmo6SiXVefzh6
1Prrx4QbRyjL2NNsxcSwwBsd4NL65f2nlHILIt45F3TmTGFjVEC05j2G/2a2pZ4e
VFlmA4EUmpYyV2hxp1FlNC7F1Jc8vo393/XrQksMNq2rry9T0bUAvaoRm+46+8GB
R597zey3a2wlU2z9D3kfcTEoIldqNGd3htx4Ec+8hEKkGMsNWzNxLxOcnX75vlAv
dUtLFa66OxrEqWWjOp88iTqBtThlnvUNw20QT7qyAzYkgOOenDnRb+2DADsjFkU6
a52TW8guLu8UGS93TmzAQMucs15xOEwstGH7OaYeo2zLEd8p1wLV+E9tlltpnyyo
qOQRL5arUs76zMmjISS0nZYcbDh+TFfZYR8j31BkAqkfhAziaEMVoMZw4LOat1Fd
9v/3lYVs7AcZKVH1r4f2azpoKVHALGzwyAj1qayg/AuoRYYqFnWjD1efPs8V8/KG
tVn+lDt1Xuk57UFbb/SB6jyXgK6F4TAQXGtazvUtDSxJj6R3MSzTURGKzCBI9gvf
0Nkaib/ve9W1De6HBHsHUjLtx/8Lk53LPU386kPJYWltJSQYzBWThMP6G5+zDqzG
ovAtb1NKuBd82IRO/5te7QX1BrNS53G6prZUR4shp5rDhz9XXokOKz1EbNMi03dy
bOsd9/aH3xuyo+nYsVnEBsF62ieeMbUaBvXZWxn38jttVsYcNaM4QHBfDniIVFIb
vDICdGGJxY9uwICfvPpd6L+4bJ6Fmdd0dZ4Co36k5wt7iGd/BUc/u6f1z5rF4K6/
CVT6p/3f/8VvKuig7atZsPq8te3uoE14nHt+Sr6o0LZqk4+2Hs379Qaa9o8aW/47
5uiodm9YTuyuVEkM2tqsi9IYvlvHLnvqqNeR/zZ4GlqlDuWBqIEIodpWLZQZIO3e
Aq3EDppNzV68QW8gJzkvPkBfQS/zPBn66WF6XZ0yxlmE5ZhcvMUC3ujt1VV47R4t
iIjAOFDXFgkVquCyVXQIGO6Cvf/Y8xs4ROUkyNAwHp6RlIMV+VSfTPKtCItIyRpm
WhpH1pcrFQ1qSUta5lgDp8TahaWf6BShArt9L98L4+j0CyjA4Cc775TBJHObarCN
nrehqW496F90lPoYvWTh2q3B9TULLfSVOpRgauR2aWej+tLkd6uvss1XMdU78MjA
6/DO02xZfD3zPtLztUjDKANLM06uk+dymDJyObgqUQEi/idoHxCL0fKEFsMpfdD/
YFtg9/zkxQzoU8EYXV1CEVsJyL124tgA1WnosXY8HU/QRafCFMG2CtCr2tBTNKav
acOiW7fbtckrwRQBTXjppHnw2NbcG9+KqyT5t45xvXmYicBTglm3sc9j3/NJ45H3
VUdUtdghRU85+5RVu/CxXxRYGnIdTAPK4KL07bL9NYJCEqpMGAq+1TSUAMiwBJXX
vJ3ez8jiA2URgZA5XW+QhHD6i3S8gI3iO68Pp3shoIb4qiPaTogSxbX/hzVCCqYR
X6yEbBCuQJXap44X0sBaU6waRKdtVLwPPr8VCmHyHZ4bRETQJtdL9Cq3PyjFhLnr
qItAjBA1Ykckx/Uyw6JxXfHYo8uPe4sbCoMZTqZXSxxI2bWnkNjWr43YFBZvihI2
huw2ihFY8bani2jpRV8y0PPczTO9SfVbVICc2HtDyMAtPWgjcQGsvL+qx/dJ4uNz
WkAekUw1oSUHccYRpUZN1uydjQ716tYpI+zRuxbzhG0Z52SekrIVneyoGe9VY9VW
tmJ2vma+Bl8aWYbBjnAkvBniP0nzyBt7d3iILOh1F7A8C3vNceo94ZXTjwcrtmmh
0lAdQ5af+4Kl59yMjhdE/VbeRYGL4jHXOrw1o8G0pzyewuOOy5Nk4QCU8KdlqfA8
dEo2pwE68n+C40sqkbAWImj2zWWk/+ZMzDguU1foPfpBsGiA0oZWYbvdlBUTP6EX
3Bp++iQTBzk6zf9JcMXUBQUFS70K/dhZqEQQqojjsiLaTzxHJE8AGdlI0smGEnxb
57J8U6Z5OxPQhhmQnd8ghFIfWRFuDWZ5v7Z3u6/EY0qs1Msu96TXL8vNdUshrgIj
wiGmUwvagkUYzHZ4OcWgBhX2eD+9BFtPDN/gn9GVClRy5yjaf46UXMHVtiYjpWsm
L1TiNXUuTUr+WDYewS2Slp44QtJ77qQwLpUTUfIuslEwn/eentSCH0OAQ6Ql4pG6
TSH8vujM/vFUOehWaIpGKLDHI04716fId1/Kv9vEIyed2xtKJ4r+6R/asy2RWVqD
wDfPIJV6lnZ34w890Hil+Sb587i6KoqkARHFk9CnWRFSEXWUWfXb8o3PQP14k+xs
ddPq33CtmdscyeX8uoeE8qEgcIH9vwa+iN8ZSs0DlOFgQ6Z7Hgewjey0kIYLl1r2
tIVK1ADnMxR9oTCjpN0xHJe0yDLH7zBhYYpK1F5FJQrwoThU28rqwKmijAKjFrYD
WHjzbblsuje8PyhtWKn5cOctHqLECrBqPW87gQLtb08HflNojP/YR0SjsIBb1ZsL
r/yoUnscIh0x5boCg5fZr+RuA+qHHi/zvLT+CZAQC9rMrZW5/U5u6i26Hm8qRI7o
rJhB5NvmZtww9l24JS/lfs6BjOHoLR7rnBgJe54K66Ig0hE9ewd5cnGqqYRKmk1H
zjkYMVTTXDfyEURR1xiqyzYoRzbTLZCUwS1uAH9AYrKudWyI8ZSNXr2uYY0tBI2R
WddHm3ydvnCh+4uUfcuFwX8fxF+JTOtr/9tTAE2k+qYyubS2pzf10ZMir0q/FiPs
ckVT+wtuIZ9mebcBcL0xqJpPszPXS/33/QxX5Nj8Zl7SNkxPqeF7y7JGaTWk8JMl
3FkrGVWnJnjWPBHgg0goBnoEaWTrufLJLbSRF6cywPl8zBIs2C1eTJeECrhNE7O0
flYW4LvV8NiwZTyJQ9o3JXvG0Jt/M5Xhy5pwMt/MKjPyKmELMRE3LCBGEDq2wJXG
oTVwhhlfNTQmIz0IfW5rugp0aTyNg28KgPqE22407KQEQZ7Ea7KJbRx13OWsbXuR
oyQuHBVqP7/vssVztty04Iv2RB0+VNWp3fP9cmBcpcKI9J9KRISiwOoN/H3tsqvV
ciL2mArCc542VbHludsgqbGtiTFZ6vlPSXLelx5xUHFcVgKxS99tYXQG1ZzmyHLV
UJ3EvjVQHtMs0+s3VS/DeYqN/TDI3WImaYN51fhj9X/8svDWic8NZFwuhzVasDRF
9PLEQHji0bcSiQXE/Fe1/mRCM0MOQ+S3zQONV56nWR9wzBF0MVEDyO8gxwJ6OFVX
QV19FQVhwtDVR8yo6qR0YSse/SNKaWOfdRSEqM09W5E31fAxuukdB+eSoN6CuW+a
KEo1UeKXgC+5LeQyhNPyfORNOxfrIgIajOV+YiM6lyCTFwj1PnzO3gJfUMRYC6rz
K3lYAWdS6o8+qry9WraKtj6JpHdue8LJ2rfSh4jr3DNS/PPJGpkRSGX9x6PkC7Hl
IdFO3rkFFQbx23coK7gqf7QKD+IORwPztFOLaekWbXWpt6/E/djLn02ZLCSkjFTb
9UeQqgLcSv7aoDeQ0UG6ORpN1QTipCNGmrTjj2hYRIylGlQxAHuyv/tP/rdZsWZ8
6lsUPY2HPOZ1pbhWaKhX48egsn5a2/WpkgxfdR6ttOpywPyAoMCsEggtapXBmYzn
pTOJ0qOR47PC7llQOCJR2vj+ucIpRC4QpBd39E1q99Vv9ORwhoZJHTzWoIoUazC8
E5lobLTeJ2UBjUfNc0FJheWt2Wl+D52XIfLxlfsvfJ01pzjwM6T0UDg2GRxzV9jg
mA6wsvxZhdR3yZr2Mu+6fh8HSdW8KfOLF0cKPLrF2nPuuLEnmO+bSz5gKfi6vPYy
c3x+ZjV2vVRaCUoeThG+1eL2I0w7sIDGkZAs097gCWJGfZdMuTqxgVHqPD72qvNp
SUAEqGyGrs8qlfHu12fQudAraOv/EuaXFMIygLJxxF0N57NnJsUO+CVVfHs3FnX/
kZV0cWVeyKLeinAkx/3+M6t0KNhK/6wxGvdv8EAYIMQSUBpV3Q6jXwaynmOa563M
kb/NV6/9NAo3Tq5y3YqLe1Eu1iv4CoeErkK7wSWICoF6gVKqjWEglK52UjGzSlvp
ajdOfmr/ZQ7xmGw2TzEcyBA+EC3B87fwcvNXdeouwXZekgxzkEGo1cAMgClTz6F7
LUpXnuMUWHtLDPVQJ06Ni2FymrTvuTcWEYytNMLTABo2mBnj1W9pChOyjOO+7Nxt
W39zwUqhF+Do46L/fDlUYlq25tY9UvsOQQQYbG7zgCSgVSkA5/UPre+azUJigg11
S/LLdgxIwXejyG8TriAi9WGZwQmTGWEon1WFDNuzvN4yosqJgffVOWKvp7NOeW4P
d26kDraf4ppF/CVqAgX2Vljwnwh6xLTT1418Sm3p9gJ3LUs/4ZO73n7k0Osgt9ky
HR0iAElTGAIBAkyNnykft7wnym6hFFf/YFaz4u1/dqx0uaMUz4MzJcqQ95bAQCLw
230qoHQZxAABJL5GGWcOIkmA6aM9wNUcyjp063WY7WFryd4F8mes2O6/XiHoxRJa
8cUJgilpeBXv8RgTR/vBStmgz+jnh8g0SHRO0DoNxExD9QUMK5gIp+nxNd/LFOjq
/cjgYZ4de3ogCGN9Cses3oiN1y7LwtCPor6+qUKg7ZL6XtDObwo4BMXMVDtM9ifx
SKPEbD1OhPuqCl7T26lwbEoEr2nNL9kLweHCbuEctvhmrCC9/uJpiJrIhQBnL8Mi
lAGA+JRYgwltzKOiWUuP1l8xHiN7xNTNhF1EwmRex51OaJgRwf2HVWjDarSklHc3
aSbEXw1Dzgit6dEup1ZlEX7A+Q4LIWV6wFiMrZ1RFrCtPSeJADQUozM3Un8qZBqV
6ujat//qze0OCocPXw79WbYLiEXpVTHHQhDDoMMC+NwIujfXOgAmlAXeukZ1Rn2u
9U2E9XnG4LR3t7v00AIDFNTNvrnW62yysKS6xlgDgEy2M78z7E58h/xEXGUWbb7Z
Bqm4RIYcWpO/WhXYs9EP2f8Aw8z572S7CX4Y7KDWoz2NjXf6iQYa8nTt2VWpiO/p
7Sl9KOFjMTC/42iGOmBmCvEUYcw8CFGOcyGTn1lzYkW8u+LoESw4xtfxsOwztgEv
6Gwk8D3PCHjLOJ4SwSc+WIPPamG+aXPD4OnGa5q2GoiELSwSPPfQS/AZW4jIMECZ
JA0lfhaFYlCJHKT2IJMdPJ833FPWiE3i94ag8xzWsFqhQhhx11K3SqJU5a4zPcrw
GuIYKQotgKDhqdtU7vSCFkTJzg1jjGmZzSZtl1aem5a3ILvhJtN6nZkhbNv6CICH
dVLWEnTbgZzhduN0v5yvu+TZuwUYbzjwS2wF0gL6td9MX6neUo4dGob2DT7Ra3zc
uzM+OCyfxC8qZyWMn+DVCkxD6uCW9ibPuY/ho2tNJ+BNRp/R5ENXbrIsLvuCHgol
JOzopJHvqQfj0m3SAvmFIrPAn2oUS15+mJZygVCl8seW6tcf9XKwUi8ix3t81kNv
OBJ3l3DpcSRo6P58lrnMhymcF8xswBq8jGnrqlzLJP/zbCXbsYs/1zQYJhr5VleP
hNWe9CCvgjmjsxvY0ppIcubbYpuCDgK0nR0oKekk5stVylXW1XL9jwDfHj0F4PsQ
SpsUI2oNtBZ+XDpVRfScEOQs8PRHMiFujB5UnEGsJvJ1/lpURY4Vbxohuchqn/P6
2PkjjNUGp7P9CUMxtRxNMfPiPhvANn6E0qse9K/mrC6ozL6BpQbQy5VDAZEYiN0g
J5segX6yMGRXQpYDqqt5jWuVqj9ew73ivOXeEGihOyZ0mDOrP8A6S5lfIVgNq8Pm
JV9bzYkILBhsM1/TCjXuszDfNoi52kSEGyBvkVZduIcU2dOInoxZsMfIhDIT+HGL
tvTxKyHyAsLCuUb4vZlbyTrGJfb+2CVnZKm/3CI2XkkXi5ehyaYoKhkgux+FwCwD
a9U8eFfftOSKbggnBupm3vlYiKmqGky9eqOnCzJRitvdObKG2Lf/g0NoaLFSykd8
UAUPnEvvHZWe5nhxNSlPa+CLmxVyeweWHV1ApTIh//gaIxfUNx2pilS+KFVF+dJK
+gJSJtP0B5hEH+dGyJg9TOYWz6guiDXx5SStrCOJbY7+zfrLA1sI6EIx84TCg5P8
B1nijVahGY45BSYpC0HGCM7nsV7FTLEb3nFMCsp9eOod6eq3VnSxJs2CD8VWIXrh
myHNm/yDlRqleGIOqpVCRwFNLPUlbcvx07n1M4elArdogc0eTbEP98nDYUXCOXZW
nF85nbzyp3Q4e4D29qYzepPaoZfZGI6gNOFnRc/Vw/hjqyq4z1p3rfRuwuQCjkif
9fAnHxHUrV6zgn+u/DKBW1l6nZVT4hgtaXmdCxeFamjTaOkG/HHQOYE7HFihsgrN
qGHJ6cw4BzIwRlglBwU1UIAXjJaEmEywTFTPVEbx7rM0waScgfr69Sd0YVkX4p7y
ynBS3Phe3hmv3hNtLoaZPQ==
`protect END_PROTECTED
