`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8H57jkC6bwinHA/3QfwG0nA6tppjkQ5tUtfiprW0nRLZ0ZhfgKudV6yPTaF/AcSI
Un+8Oa1mliHB0jfuOsquIw8kCTrpvnUpUYrFJFswmT1FH+hOVbZvBkqqCURxlL9M
sg28ikcuFDnWv7/Hm5LMkATkG91De0KrXkklaTmlOXYfi+VdKUq8kXV+DkC4HWVa
JLmEOxXma8ZLmRgXBdunzAUYOLfHvU0W03v6SsRa9TTEpMkNpQDDYsLXqay7TcNZ
KDD2ho2d1Z+tPfVpmbEB17/EsuZ9L3vulpzpyJrsWqgmLwDN9X8WAR84C4CWX97f
Zps7ls/jVYC/aTG662Ier1QIzYc+wJyD1zZIaBd0y0IGyx+8jDc4FVdIzWKprlh1
MzlkUG5aXc16mKjyjdQ206k+WEDZBEfeI1cNIORB63pdrET/Yawt/sJqCQCQm2M3
b++xcbMnIAxDD3GrLa+e63iQZ3EJtSR1Z2tgGDpfCBQt4TODYckKGT7576OscOYN
rIZSM2ohPG7ldYmFncO2BGLfbpTc6ecalTw/WI4exqtAykOV8zQi4oh2qePB7Wfp
HnmKOnWl2i973W99Y0FthdAc4dsRGuVKqmwL5/zjHM7C+P2+yIbip6pkoiueLhHR
yfv4KvQDYNz3A7w3ELxmF1Nyg6hZAgOg46QnA/XOHVXJxECsZVp0EwcVDBOIcp5T
RtABYJxaHBvFADYtMxDihw==
`protect END_PROTECTED
