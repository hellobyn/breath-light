`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SX5aSclFb+GlWaOJ5pj93nm5rFnwVdRdjMJdonXqB6yR5Fy9Lks7LsjmybJjmd5N
JLxYzSc42KswVaISodyXb4l4BtsgJd7Lgeu6kPGn0tTPe9xYt0e00DSYe5Cp8931
jY+T0qMGhcai5IxbZ2sU29heWJVLFsu3GuCsxtS4RyKFrE3jIFHMGLPxNu1b4OEV
qktkvgec/DqR3R1ntRA/5wI1g89WfriLsQi4h+3B8tAEGrG5WrXPtvkcsq8eeCcl
Yjy/GdL7yEKMg9DaDUDbxsU7UQvDeCQRhrBHjXtdZr3GYvER/AInUBdJW+6KWKD8
6+fmQdVSXGE4QJ5C5hm32vDDYDLs6MaqORFyk3V/xqAFN9yFePMvpsNklrUWb/7i
YIr81lYx/jIT6zZMHhJQ2SAZZvM+xXGWZxL9RpIOclMDXfFItYMw4NXBg+Zv7NLG
6frOQ4uuTT9uZ3yCy6Qu6cR90jY7LsMP0cl3ue7KEfNQIOQw+TTf5C98MbGedb8O
kcM9VMmqAxlfsSd1TJ2xmSvuyHQpAGnD4DeVjub6MmZPBz4mTRWDMufYDWc8glnL
FlLhG6+VH2GoZdEIeu1CQHy9b9giqeia0cb3Qou5uiEGEzPvZ7l6nQ7crjvX3Nfq
K/FwimE20GI02aph+z7DPf/YoMhSUVQCP3+7VQRGM4MbVVAtpwWdLUgKDaBwkok5
zQe+2t8osRZ1GCOw0EV5J/Wmaah+VpnQJx9elQ4ds+kCO1OgTxZZjXy/H8SrAjf5
vE7n5SsJEDef114E91Iu92c1xLbh+TWFdIQdAG+D6HIxAcYG5xWtm6FHPOjqitCc
NXwYqIHfDeLN1YXpVSdmqvn/MyH15/ieiLvnD60r7am7wKLHOT486/cjCmgdxPTS
inwrP9sT3kgvtRSt+U7E8ePget1eOCHgMqaSq9IOhxYKEk20JeBpIXPpHexxtFUw
YMMoC6whzTNI3z+6wY91QOt/FV1VXIoEFsoxz9KFf47k2bQXb+Niq1iIKm7oIVRg
huqrLZsBz/Q6fuFUTF+wfj1MJ5JjfHjtXdixydT7P+JEKa7J4Ubd7ShIHkBdbTDd
4Xp9yjgGNHK9+D/qOz/gALF6a6tIjXQWvdhrJN/Q3+HEZwb4alvD8Efmn/AywQkI
vcPalwwSpwJkME/KvcUfr/Aoahlt/sh6PpodL6O6+X0aVB2LN2fpmUKjE/b+hys/
9l9BkQuSSpbTWbNPI1Bv6i7Qnnc+4pElH+J4i2cbktw7ZkqC2uN09w9JYH9/aBv5
CUe4tXePNnFOi+4Kr0kBPOWodoq/qPK2eYOAYtFL15bbk1uTjfVPM4/ZqvDb0i0H
fKKMyF4dg7m2WF+LULPBgNyYLK5BT0D2lS2sHbpkYfyjJvc4OD/FPMHxVen+MHOC
24qPhAx7mskfib2twIeqK3GS5n1VPaPeqSqQGwtH/6mFKnibStyQIPU58e72Emee
jOVU0DpGuBCRA5qaenFQW5RxhW65cilbzjLIKadINmhOlgknLJ4vjsr0slUHAXmm
7jcXoyiRBSiCNe3AhqH2Z2xO8xrf09mVdOt8Dl7MskQjQVaf4sxUMjuxQLyE8ddv
6M+jA/Hm65FbM79XB9UpOrQAtEdRLOiFCSiwlMKlIyeOKxO59mnWhRq1PVso+I7B
uZhVaecAvBWgW/h2BGMtZxV5EuHRGGbtWyB3nlxiuGpJ7qLiRQREoxt/ArYCrrkQ
g2wHGhqZh+pmsVTAvp2I4dg/asNdqjwyXR2CuQ9YJ0UiHdEAcAzQ2j2eZ20WL7zt
bvJc/LOFavu2qlfLQZtZro46DKLoktI8M8WZ7i5b2fJbMppKbYNMUMbs+OMCNnjx
7r3WHKmzuJxTXFI1XaYGfif3PeXoPo82jQ8W7PIJe9bMbdeiDy6e5SWQn6/MfnA3
/jHKk49PpXk1DdsxrPqmfM7EEh6sIGxxJi9wT+Rxbk9bmP4EVuz0PQjXCfYZZDO1
56IQZHUPnOxyXmLgWYBrFIZ+Le2ff6fpUsCHk6m29zCFdHFo0/w4zkhenT/qKw5P
nJ/7S4hE2pcmzaQOtGBtmvi6bLuqAS9mEe6P0e4n2fb5pJkDohmW0u39PNpRTWyT
0vDfPNItSDhldqDPZzyZLA==
`protect END_PROTECTED
