`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzmkbRE+kvRPFCbNUeyN9xZSAst617uYPKh+EJre7baJTNKFtH0YgailU6UQ+eWR
gGBqb7aptyCP8Bg+ktiBBZ2gJOfD/KEmL6X41Iv6VYN7wRUHE2of+gXzT3KuK0O/
DG4lrPiayUvSJTphTbnjBvfG/YczyvCJyUQQBzVlD+eOU8BOrishf/98jJdUXt32
CnNCEu1ljk+SfGB+deOD0jqosBfJ1rSWH4RcwAjcW/+AI28wSfiAU3kyMOOfRW3D
i+kT8fpJUY4hwSGSziAEtkQx+lC2TJiyr9+/fqwb7c3z8qU49W73iautzUiqsaVT
bkla0jfDsY45O+UFkCGaUpFsBI494CXLqedTMVm6ck258u1lSLxQsxwbyQNVF6nt
jfhJUlU2IcIAI79pE5iREX8kpJEySbuSlbCMfN35XFIjcozFLfzI7bpSyFUPkOON
nzkMKRIcvO9PPp0Jg/dx8LEcA9bAXxfBUID9fZaBNTqohQjCHG93NJ3fxMQnE0+6
TH7rdf4qwI02giTOz1OMyi0C/mAEUCgBdDWADVYjxbgimr68mJjc9/HB/rhzywwb
3Zpg0vnjsjNG//KnkT0qvuyeIEDJvENZ0ToC1Em4qwHYFFO8TyXUjvGYYHFecoFx
/MMm1EY5XRqWb2g2XQjDlL5cbaPmIE+IWgTZz8+FAdja/098eWAPn7IBJORNzLg1
+maLKJKJGLAl/cFw7KdQ7BQ7/vztK7x7XFEr/h4ipWG1fjsf/uWmkViuG7Gcelxd
e5Jd/chXsNwRNRecdeTr0kQDgtZa17tQDa4saI6E1nASJ24/f73gEDyZ+z+XcgTc
rOhVPOpK8b0pYRnlzZYml9ucZ+oQMR/C7QMJFZHBHjzoT7ziVYU+ZVKQxy76BpEA
fZO+4ARs3bQYQbhxLqKAss+oMny6LoBzVF+v5a4JrWFoNrBRvrLG1iPPCnSsGwUd
m5IdcXfPjyJdsG9AOYqruo4kAGGFOKNOqY59OPHwR+WnfLPPHQknrMLJLLj131DC
PJwrck6hkN/LG9oejGlVto7pqG8vBdDp1blSlEy2WP4nJhwBRKaIxBZHrUFjm/eb
6wnTK2lRLMp4VsVSgE5mVLYw1xC2Xls3TUN9SyykIKKTgjpGOKcW9b2CTjOz/uXL
DZQWs5PHv2ZRAzTuxQWRyOKm/kCGO6xaar3k1l6BAdvfC+wjkw6XOaLWEdZYANMM
hHQhUXOGHSaoXIwOpuAs7kdeJVSCd3IceBx5b9AmP6PZhILe9T9LrlhrECKrMupG
tSSq3mRw6pM41ApODHTZvWlY+fYzsX8tyR99zIOLWKNRTpIhJZlVNCEIM5IpAODQ
cEd9784L+h+5Wwn/CTichEVdVxDWxXufLdYzP6gfuN0N+wRH2xbGXoRNbuxvDJAB
nKqsO6uEh6colKi5uZb5dJCFVC1RGQK3JU4GC03q/kx4rFZ36K94Hpb4cbpveYl4
CJCah2oJEHyqo8M2ZaZBWWhVIBQkMyI0HizWemx+nFvitldTwX9x+jqppDbqlX+W
xrdrfaYW3K53tNpbcHaF6ZtxMN+iKVSkYAdel6xMcSKekQXap8nVApH6arecunF8
cu2k4CmzOOmox/H+DuCsr/Qh6H7NhnwnBI2rNmOkfyJEdmThxokayP4wzn8iPHls
Qe++eRDigX0L6iNnE4P7kLfnhlfkR0MzqQroy1kLvAHhG6fwF6lRO02XrjWt8P/+
A5XUP858px/3PnQXk01gExzIvlYLLDUyLTCmgxcJkraNJasDWd0hHu9+H0uA+Fcn
lwVQ/MamOICvpUU5or6kgb+u5lVgJPFpHfjShGJ0noyXNoecVneKh7CEtlKmDYup
JbR88MBThMCzM+irmGvPxirnXz9GaKBM4z+x/ITcIsDlZ6FBJvRDOgASU2YuFPnS
ny/bcoA5J0GRRvLzXa3Tjt/Sy8MmU9iMviMdi1KYPpEut8bLpBEhdRyybyxwY5j0
s+nZr5Jqir0mYPL337KCyOAQ0JA6lOvj7maICgeNqvoqaJDOu6d0YlLMTiB4o29J
ENLkugcXCnYxJhLWdN5B5uO+tKBV33lLrB3rpxcwv69VX8bvrLwFQ0WmUGDZpZmh
PIBdFMOqZpAcTEw7jS83W13qMPV++1sJoh4ZSf7y+C+Mlku8XO27NmZA83/Hrc62
2vMEuwMCUNjRrVFEN3H0dXCb+1dct2shuQVQqlxxjucPmmp5okQapumnxGqLXtos
YHsDEURbouSeIYN1arfNJsyEb301Qhlj0+jMKW4LlIDmCxp8GVSPsBuM1x4lDdoK
fBeA5YQ5vUffrEUSdN1Eqzwvfho9eJyPgwMiQogPVYOSnrS3fVk9A8UlRyVNqM9V
5DIW7esiUUeT9sZ64d2Xkhva06jX82JQMvdsTNJ0q16snFli5oNkJVorTVwPzMB/
xawhqNtD8CxC3C6q9GK+wbLXmC2jEpKqbidyETfilzl2bQQNeFXu2R+/DADB+9Dz
5Yh/Nab9WtYpmo8+KDLPomIQTPv9mqDdmnLxdsegJbIBiGjXYHQ4t97mw6YcSRA9
xjoujWx3kN0EA1uQnEuInA9H4qwhBwD5bPy/EYNxUEA4bKXPJ7DmwTjfJ/Z5hLCJ
t7IvaNT/uquNSE3vHt8NENltc9zQv6TucxzgUKnK5UDi+0xh/fObE1go/Avl9faL
7CZ4q8Dr7n6YNgHPzkR6pddONtu4YFf+IlYE34y7ug7oLxiLtzY665nXGv/WROOv
VEebmN/mg0e7TRU8nA/sd457UVQhXDsl5M4y2IBBfR5ex4cXlQ7Oiaf8fZGFtQVH
b+tV2W6mdtewaA3ToSbFqeuff1LLIRzGn33NKfLJtuu8TpR4OzSXI3MH8O3Y576T
pOwkC9Jnin6ItjQVqPLl8Hfx8eUDVNl+8oDwVeWwgCL2P9dSolPoPo5mEYKbZErZ
eLGERgKwF4K0PZyW+5gK6MMmsIQKOCn1x5/qrbL4hPbUMciSYPzswFoZF5tGFHB+
dYGOBZAK3tGXc9zNCnFFVRqQSpEMf8O2R58WpIP0ZoHZ3gGDWqivUy5zUNqez10D
xV35oKIHwpzx9mu0rK1PZLO3sldEPd4FpGDoUALjpis57EOv7Z9zoXRDIvWOgeLF
AI2aZVL2uQb/YL0sFX5aqZ2Bx1DgKPUnEY4VaXih7o/6w608GhVVXSnPhtl/6Jxm
As4VvvWpq0FTctLuP97D9H6EoHlwmjBQY8YpZUM+3cAZYc20FuwVXuyS3N0RXUv/
SAU+u98YKKjt6DUdh/72MRBVof5byWjZKXCoqsg4sGh/8/1D32ZFw3h+VkE8eIfO
32G7fn9+XJjquGVYVwL4e+9u0TrJpBBdPUB0t27YNyb2/r1jJFi/Qe724b2PaNPm
A61Q46czml0saGkGfi0CZCTOU4E7MKtnIdVAzMZm9mdqPT/s0wCuLtCGrtVjlVtW
eRjGJGVbZh3ljvNo2jwKWTeAF1+Lxz92b//uRfZp+2JRTqDO0j9Ny0mSSPQNbb6z
N6EO4wyyr3Yygg4rVbRgP80Nk0jOxcALRVgcsmYfG2nyd8URZzjvL2W4A5oCVbQb
/PmHTCnP0mWxuUP3DXzL8T+yoa2bppNKE8zRLsSLM1OwhW32rnEZTcgMiBfOC07X
UNtoxxZosNb3oaazoXETi3dwqDSUV0I0NeywKksvddpW/oWBBTLkntlObHX/oB6U
O1OATjc7sX9kkq12cbTZ5GOAFFj7N5rrwEJIDP3aMLXrh/pNiQL+qfN6fsDa4VcM
UZ6kHIig33hu0v9xGs0TIGJ95aknCbmXiWH67Kg5GnUXj0ZiHAnb6uQRmLmNT6Ig
YLT2/DiKVFtQlHYGNr+0/xEq31Ag8IK670ayyrRytE8nq6c5aFzg4daqvYKyt7fP
3X5AVa3GIho5cVM/Uxp1j8c8cC90Eh9UD+0p7eTxWqo9d7SJF2R9iSFOGn8Z4Z9q
ME6YPiYvo7vcmaaM/XaE7Oc0zo7fOfgg27TT3F4BTki4P35BbPsTbyFag+e7pCIN
BKeDmmuUcCO9BWjqkEiRrdFHzyr03XThkSUyjut2NpccaFH1Z8d70OX1CXqAwXd7
4hfKjXwtMEgy7WjqU9qFI2XFTi5212GQYovIaYWx8SW4yJV+A/sVm/d2LyfTFE4K
4e1yQObqAcn5Vi43nXkIzhPGJujdlU+lNMKHTG0CWtSRpMOOZNmCjgrjTiQ/8+y7
O2ty4JKq//DpSSO/WKm/b94QFql2BPw0tHrsAaOM8/BF6PJq0J6V1LU8SDJBsucf
0oxafx04RboKnUZmUCzfKsbpYRvxrOTMp1g6EImhqf0tTH4PQuRx3xhbuoL3lZiU
mndultD9fE767Moa0LmkLHnJjK1bvOZYHZA3SpDv5TorSm/LndVUwP0L5V2eC3yF
Iqiuqsv31B1CfBkOKl/pJnNzfaET/w1MqMe1X+Z/d4yR1YX2d0MJibbSCfx1eIVM
GBaflkguVXRGfXvqewfOR4J48zKvb12VRDUlHIAtGg/nuL/9x4YUyLGW8c9SOQAr
r2XPbHTz4JpubK3aH9L96iO9I78gDOLvSkHgNS7pDhHJCZJULM2wOz96H4itcm3y
NR8gokqWp1cV+wE9wyCPyewHs5VQSzhN1rB8DIMieV6noo9Z95cwX/oZ9uhghArJ
Y3hOwtyDDEzm37aTnmMXszkvqcHoLw7jG9TrZdtmtOG7Jht0ey24Q6sLLcdySjQG
yNetFbW24h7DkKjvz2P9TQBvvU6Yk+9T78Beb/pkNAtuF95VdX6zyTqn0c5oFUoH
rNfMgCA0x4W1b9Y01BKX4G8C1V7KBKexLG+KHqoRC8mCfVeDxda0sKXbV59gaFMT
XaoDFgZ8ar2RQOaP3/TWZzKfweP2+cs+lPumk5lhtPQBYrTitMhPj3o0Q0aBNWGu
rVM6pz024RWzIwayVd/TqKpV4L9QSWR4cgIwt00VmZyH8OeKZ7I1mfWFQrtDQeea
adXCH7CzUGPWD8+SytrGlD6TQnXeX8v2AUJGVJR/zGJzwzfU91zXmjJwkI9zwCop
nLHwIvbrwo+Bs6kuGIUTyg8kBbeeSqvGe1hUnBr149tJ3ywTeXxOtPhoOiu56ImJ
zp2TP4AJUItgCDgiPbk/q/3RRSDFNJbm0m7YqnF02oP8kAuzSOlG1Mmkxdhycjjo
BqaZNDDhGgczM0ygjxOtwiqyrA4UTIJ61CLpqgjiQrCkEv2h30l5ngF4CMYDxepQ
5vLGNbMjEkPnQrIS0F7/75Y0wIMLjzKe1pAfDzpDNS1p9ez415hyLERLOlwhuCdU
mVsykXiFDPZ1rRWTf+6PA7hVyqCTeX+/o0dtbsf8IMlmEdcT2SSZZjDCxWo7exVf
H5KIQkSSEr/1lb5Ad+aWoveCw/l9mMENHh+ruqYuILFt/G3Y/t+sJMo3+0B8YC8m
WBpT98lmsKbCJSd16wi41Bff9lNk/mnQ5navv2DxxsATVU1jCBA7uOvSBnXOu9CS
4drr4yL25wMiqL8d3i4+9NcH/40IYG22lYKAijmZ3VGgMHsz11IWEOCOhd8d95FU
YjKAfWkjIRIe5HuHEKGhpzEraAGwnB8VWSAaff03MNuQ0tjwQe83Dw2jE4kY24zm
X/c1sn+eEnhBUQdKQJ7/N8Kg57hpYz1MeFjLNper6puWhl9DSfiVtRIl63RXmVMR
0F3UdyicD9JlCcVpC7Htc4Aw7eL6bgTfg3iF9zEz5hS0xT5oMEMhkqNBXToaADqg
p2SNelffRVlDF7CloP4hScqanEQ7+8pBY0l7HipgAFmx4cqj1r735i24HVXlb/Tn
dS3P6NL3R00eIe9KnLay6hQQJhK8zcLTB9PPscQsY+1fw7h4vzaWCQpeHWNMuS9m
dqD8sAEHZApkNuq/7MeBDwCCVIxgtInB75zAC84YP2YIuiLZzLVvC7I6e7xQuDNC
kbKJnsCAC0L5+3eWj3/1gXSViclAO8OdHEbxAzOYON2T2j7rKW0lefPt7XZcphj9
0tmJU4EptoMhFWAEIF777wVRN+4QUlmELpPGiEncx5yTVgGWq1cY9jK86YT7nHAp
HaaorTDHm9jx8a5M7TkTfZER9T6RPH6i5hIqJSNkGxaZ4i9ApW+p7qYLez22zRkY
MFK7WgncUv1E1qialCMpHydWlbSa+J4+Lig5Tcs8VmeaPbWFxyOnJzwgI2ZJgome
u1/1T82OOEDkqtheSrFgch91m8GANliNQGDgGqFCjDkOXVyCQkiJ8H6/ymy0C4Or
RRvJOft2bIVttoHHhQXZiTvecFPUD1mfGbDKC5jinqyB0wf0B6PtdhzFEnDGlZhl
JFA2s0IqrgMy1IFEDGoeMU8NgIXARhcrieOvpk6Z2bN+m5AzUxXeoY70spfrM1R5
nUlff0TeuWfHuco+mb0gA9y1LlAfGwWJ8up3rQDxM79RLVzP7kqONeBlmBUcyJVe
nRPS12kJ1AumphWK/hsVJX+8sTW2CqdJj2gENjshhrUhz8tvL1JhEThpixawI8vh
b3EqR6jTa9wxU8DSdL0pidH2KkRfSmQQj/RJjxYiwdkbLJuXoHvYGcSB/AoD+abc
YEC7f/PJoarzGXm/jiNOJTtdtPOL5ODSnxYOzm25BtMFd8/JSnD/nR6M+oxFLXYy
VYcgtEbML8Feb2ruH+lWDo2BBaplNKLytsEd3mwQx5VUI3GjWfyjxI/A1HBw27YW
MRAP6aDnqkIa6cUXys/6+hRqewzLJq/xwsr0l4HmSwc+I2GCSXDqXX9/IBL+yHBD
6v2MP68iKEO1LG5c6ctk+pnDuWtanvA7IS2M4q3v6/UdKACq72DAcQsWw8U5BIva
n8rZ9ODw2ZVV5aMCDjpK4jZV1B0uMRNZ1gLx8Kc3OYsJGeD9LnkPyEJLnhZ54Ncv
/VSAO9JtqrsAavJhAm4dWCPEOxlHzDr/WSLbVWjwvHsdBg7Ed9tHuB2nxXawn8HY
GtAu0yRxW/GcSvwwRhkiqfkH9kTQwOF+iz9nZeMq9fq29JroZ5uobwS5Jze84Z6r
GJ0ttP9jKpC0xIf7BlGl6NBgkY3lJA2viDEsEgoQwhMS2zIV8bpi+iVaLGQXip5S
oYW8WqdNNI7GKsE0kUlg8pkF/jWTTN9KHjq0RjS2mcK/S+oabprsQny3WsOjWVDA
oTaPkJTZ6wlcfAVqBHSF59ZfQD/dGdjsigOmnnkwKOwerU83UBfEw23pHuxIzNyM
bB9jCEdnzkOtgzEf+uST2gS7apWYrMUFemEXgEUZiTBMxT9iiMyIp79IGt51l8bc
ESlHmK4EsNEFI2syEcKlRXYrpi3wdCRejeNXn3OmAJwOsbxwKdD3iHlzfopdjW8e
jFkX9AEez//yI4U4i0kDDhIkc/y6QwG+SuFYep50gvTCofF5GSdc+EizEZtk/HgC
tFcVhG47ac14z0Vc8Xw2bQvF4l8e7ruUbAQe+Xe5xPYXeE26zYl/4WPQC90ynKXV
nsZvYitM4WVdMcY7SRjVBj0ggHBRFpFRG/xr7Hdp0U/GVCIGKaTfkFFzZaJuKU7/
MrkAxZ9VT0gGLJ2D+xwa2r8LZgIsJKjdCybB2e8rRz20cNMPp1Up5vzLrdNW75KN
O0rpMZK132yqKJiQYWLXfokp1AzeWSVNgph1Gq0zgs2cLnxhfWQK9/r3EvKzKAze
rHpRfSh1pik1j7acDbf0xTDNmNvMyFR1HM7HfMNkkGC9kvn6ctZZZqxUfO2pEUlI
ETlwMtUqUya1qIA7a3zrAI2uDgy316jg0Ny8l7BLst7V7w0GngX4omW/9aHUvKi+
SVBv7zCYXcw16L5WpKkGbQu0Lk1lsQg0u7pxk9gFPOiKhfAv594RImK5vLtQTMLY
QfpaOuOoBsWn5o6tt67IqlM94PafqmKgK3eqEzvJw7unSLdaCnsknQTPxPTaCdrF
hxlFqgSIZ79lgirWZhw/x+jRJvwxs6IyWXhDzp76P1y8uBVppafW/jt1kj2dHWlP
0T/EAzajVKj67PqLaF4seXrzZQonvaHuwld+hiVCaTXcrfrnYdVv67XhhBRDLtD0
G/HAo4oHuao2WlNWEJOcVfR/CwAL/xBkSRgyLI5KqaszQj8TvfUaRTf2jwEYUG1x
bdzA6C+LtKP53cWrpYmjOal+DMIU6W55oDYNmOBOHMyEs6a2PIiBOhJRjhJm5WDp
wy0tZ1zax2cPmLTBSWzefOUAW06YVM3pB0VpsTIWKd6yDCpS9XrlkS4cN42EK7YI
COE9uPoUdebHUALzvpYvl18of3UvOaDQg4Vh1bN3zLx085BVep3e/RnGep6hEeyk
vAErpVh7Qas9Udcdt4dtWGo2MhN6WZdVbAJVBskEks9R1Mxk5pDkoUveowgVHfbZ
g+ous6Cjhw/uLVEM0+uHUySanCh4E0ajRbJiSbvAyctvjmJgfCU8xRAQMPp28XzR
Ak9fdAIKcEmbTs8ugsdIAtLsVHWdDij1XdfcL9+hhbWFI10Fx/hd/+1T3b/mG+T0
tSKxTE21kajR1M0YSD9XinKJ7sSqCKSwRso31+IW+m0C/7Oa5+rSKIOLzvPkheBs
YdhdZwUj3JrTO95CZ/dYd8HeLBA1S9SRar6iBZEodWv+ERfCe0ZH2B3vJn0qyUWK
re3Gjy/055Qej0nfyl7BEVsCu5YVluTtTeDgA09QwkcypQbkaL1Rtr1t+6cC4F+/
qkdYCdtM9T4VD9fN6er4AqNWbcUx68JvTH26MHLMwEOXpr4YxZpSLCItgXYdPm5Y
pY+pjlkcoIP8Oqzj8yvYfNjIAJ7MHiPzdizdq/seFtPd191IOZ0lkw6JiQh9pxh7
7TLhBtf55+PplYWCEb7ZwD7YWFaEzt2Lc0wo3u8TYsu/sEM2NtUluSqu54rH1eoa
X6No38p3DJaLeHh8jUo8wfLKjdVnGITu7kX71dTqMjTdMou7w2PiQgiNIBwEvT6p
5bfM/jQIQBp1P3tIFccq8qd3/1Z/G0DCqxYeJ+ZR5qKiNOKqVt8tKO/L1s52rzsB
5MkiOvG5AWT2RIL98H2vimX2RPxAuMRYp0d+/FJIcuQZm7+0zpBfyuCyMby7Sxn2
V6gZ2jjqnsZMRiJdXc5xtJuZQHrkuyfRCrTK1xurrUBGJSh2t3zO1E1Wa3WYz5UW
fCbNFLctcY9eS7DDN+1aANm7+1qf/BikWREaiW12WpqNYnbdAarEFNZIRm95n+E4
D6z7PgIP8WD+XRakiYrRmXGi/+FNst0cgkJqeQbETnk7byimBoFRbujhcplNejeI
bJDI8RD+00brqWV54ZT8i9OUEnPWuyFsMyyxYCMGd6MFAr6xJ+1nCnAuIvTM1oLR
Ddih7mh2bucYZ5Xhpu/zOEpW7df1HnWzQrK5tI+oFhvyNxaS7jnioEXeZnfepSn4
j6as57noArTkf9X2vkjaoot/v/5wqUqOHuZJHq27RjkPEso3pD0GjvVTc39NLKqJ
XHmUzD+tYhqYEgCsqNIoRpRb5mL+T+44e494+4L6M66HZIoebD7VnWmXM6gn0AfT
8AcTN8Ppo6xT6WEIb3kAeAfccqUv6y9uUM8gmYjFa6mvHNde9RQGsNkzqDNZPyvL
aHLosUkfyFdnw/Dx+06Bk0PUHs2R7XPTb1dGlu7SaidfNA5mPaIb2+V5VqRq3hkX
fZSsRCSi2iIM2C9c8iEar9CjRdwPOGBkLHK6vLNgCy7WNWJyydEpesFgFXNuBtOZ
ofGWSQaPThCG9r3Dp7Eq59R5d1O5K6uNO7yF5Uebh4IFddd6PWaVNQcKRBD6S2++
yqwdCh4W39Y4bLBwlMt0pq/FNMNZZRqFRKeeTN9y+q8P9nWt+jeNJq4qKGqwxTma
jU1Ud1UD9SD5kCgnYg8SYOc0/a+oHx/p24abishdITeWdOA2mNsMYRctVBEZ3JcX
mkTnk4dbkhpCgXJM7RKYKo0oijZjXSuBwSriGHJoVWhfdGkm7dJyLAarTZNh5kQT
HCSbvKmPgEYxJ1RgUv6eMlOu0syLYDrCL+w1xjwG3bD1bg1knMrd7crY5ia2SLhn
DsUFx/J3uzHeb1S376m59CXJsZlTevM9JQQnmETvJsY/mOdjYo4cgCYr7NAiDt35
bhk7hNAqGdLuEcCVzz4bJbHDhFuzquCLhbf/aFl7+pTLtIiu1J39HikW4SAs0esx
6SGKelUPKwecJU8/cEu6GNlqPKzwzjETAB6rQMADh2zTsHGFbhkz/5bzLHwsAXLg
VBIEbOuFACRvZK7mgA35u6qHCKjEFmD54eYydiK6Yr7chNYGrhoSTLpbbwOHmpBJ
CVmMKOCDulUYwAB2L4Cakd0wBUv+VMVB+9Uqvfda/THW2jofXzNaQoLXpl0D3nRh
U5ZRuHsps8XC15tbMj0BpJIzJJUCSNl6RV2InY91NrLzwaD4kAwndP4Cf8+u7rX5
hYXAZGOYr5u/BFXIKHs/bNvIVOqUJlo2XqAB1yba33JBCTrenFNUkrgG+iRCxbv8
as7km/l4GI11bZz33PjxEWXfXkWkmS+AdcmqLQUsKiRqXuHCCyBhkVe7gjUhYpL0
BK7PoO9ZFifN4y+IgZ+nR3RKlRctdI5OsejC4FG/zOEbAqdwKBeMjSs6r1B7Vso6
Q9ZRVLSrq8bRxIyzrB6ehCYagKl5+yS5luWM7cr5bUSAe8bdZ0nlftWyTIXORtlt
VC9QL0a5WgeQUpGo0iXrvyrpJpW2rfTZEddN5s7TYJB95TSwb0x036RVl0WG5PHt
cfGJCV4KkHioKcgbi5FwoIJ8iV+ro+slMx3apsMLehBAPUij/fK6Aplz6pgax4D3
m/73epUBociDjeeQDJLz3ya39cwnCsCQAmpLxbbmQeVJncFcoz7lk97rN9neKYO0
LwKe2mmkBkOsZcP4L9/yPO4qhMFfL8zoMJxmOtByO+CjuXr78dorzmfO7UDcHan1
E6O3fPH2Y+qX4EDKQPhaugufmDY18sEltwpjuySfJ/xu2ld565Y2nA+zKG34oD2H
hkK+c64h7PBzJ2cfROn28KWT3sz69vPcbkgy01M1nYNA7pp2d/A+lH6uMdxbqZkI
eeA/twDFRaA00NOv6zmnpaOL0b/MhjAohRKZIYSXyCdyxxJU/axgvgfSHoo2yiYt
DiJ88ANENy/T22mGiuDxVeR6m8gi2mSiHTbY2z1qd/4kFvpxely6Qa8ftMnhsKJ6
JVnHsVeB/JEJdPtiSBIR+iRv3MXtKyt41C003tJuomhkCKivc6Fnaan6d+q/b2R2
BhM/o3lGSR0S8v9D4H/gK2lzM49XpnPW/dvxlgvLfeG0SQEOHS3rTSH4adBHzB1d
aKjNpVUpkLqNlww0W8LVGNZMP2rG3SRZoI2HFtc1HS9STQazavIveVGwJraH5z32
g5vta7Dtc/l22IPP0pdmQApfiuUky7OcWIIyItNI0+XT47BAI2uvVl6HQ+gUO0Ww
PvP0IIH/YAAWuA9qdwI1nOq6n7jCK3rCGmHAhmbIKqno4F6P4qGjj/CkwUhj7SBW
iDXojiQU5ygT32xE65PgEbA1QTK5PDjZZ7npFhxnKm5td2iegPFSFoP77dTOEXr2
OM/6WSgFWdRCW3ShDRRKyKrr/dnWFEaHBRc27Uk+lkOTF8t7b5GXHOKnrQjqELjR
bwBXpQlvqp5sFNZwbZ7rRJKaTlGO3ad2gndv2JBu4vNJG7rMhCTG64Lm3cPuzcfy
i7i2HTc6p3LkC2eAghfmh/t2QmG7gw0oHc8zk6YgljzCY2rBQTWPXZJ1aSbP1LGo
zX3FA6IdWqpJuoMnnjINBxmzleMnFeEliD2FWRhYPW/0/R5HvRR3fJ1MltMXIfDr
hFynleAPm8WHrhce7NfeTTRE7d/pILsUV/xxFKXAvURefdd+zxd4Jlw4eh3yKRRK
d9/Jmm4Lor3EA04bV+bQqG54al4bl5FZMmE0FNOIAvvkMqc8g2c1LMcPMIz6iXiB
2IZq0LbwQjLaEGuIsxF+AmzVtNx5stClhoC70oFoSC2cyognlJuZXZjhvcsPleVj
HsHTKjIu4W1zz4fuCax97vY+U6u1qj7GF50mlXcV0I6VC+tVtclY3EiMwqn1YK+X
QUJVoWQNkNW2TWsxf0D52l77PWOJrI5X8DZ2MipwClewX4vvkOPeGTPrCqFB84v0
dBBvqnlgx0zuQnICwBlv+xTLa0ElFeoSZt09axzLzWwD3wOa9OiztLsm7BkugaOz
u7w85Z31Xofk5vB90uOj347VxP+JxBSD+GuBPB/2+MzC0h4OAIs0J2fQGRVj1gMC
74lnXZjy2pGjMi/Q7WzOEdqOsmT9SCaygSjqDBOrV03111S8ve7xaEDTaa6W7LR5
ALFc/gaIk/2IAhXHaUD9oaP6vsO+tEGIi4LXgUWgZ0zKS48VjqILUer9kps+IMrZ
eE+ebXM9sVdGyJHzr9k4SCv5vQ5KfecsdUaHc2oKbGn70G6cgkcM2Yz8bZY1Huol
oykqo5/PSigdVt2UYY3fbZYgdaNQtSgZxYs1/d4/bg2vdddGaDMF8BxZ/WGy/kJc
jG+/1ZTSUJPOHLZc+Vadiafezkq+sXdtRztAPWhBb8Wh1eYhdFTA5sa7Ym6gLvFU
3Ha7U2kEjgmFnuwz3G6R+cckvNSFEmDuVNez2K+TBeqHNW3bZu50ryLP6t0osiks
CVMd0ZkZn1rNw0yx0Wp4Z51Ob2AHcb8PNI1eIm50nz8JTPgjtyBxvB+owWKpZq6Q
R220e57axUrm8+tTskiFqkHqGB6ru4OqbdnCzNiofV2W/HTi0Giyvp3jsdG0qUrg
Csa2vbKDiqOmLTruHLsWscCzfqzlLPMZPraBhibLNf7rzwkGKmx8y6d8eG1QHGGQ
M5vCi7EW3isr5DJ96iBkpNZON+i1yTOe2UJi1ESha87HVxMPkGWLgonJBqs8qaJB
zU737loMNm8p1Xs3t0E1uorapEiAiU8lNWAbJ2UL/OLcIHSytSuDd0oQGSZ4WDzT
5teInwg9otzrTErnELn47pmcJ/ImQnDP5XT/ms4Or1qMumgchf77uGfjA4zglNZJ
pyuWB1l4l2dB0QDO96ftdsrDcXnAD9CcZsgRVFUTnkJ4RQ9D9qbb9CicbEMi4xBB
hiim0TqjhoHnTG0SkI8DxlmLcPbQGlEWm+khNugU/8uiKKqVegM0IM0DO+A/5dtf
Vh+6bM5gkDOLycstHxtpoC+85zMThMjW+y7j2zBNYYU9+Jwv9PFPVkU5SGXiRDSx
Z6oPvoPcuY1W3vffsxnH4kWkUoO2TgCoehT6hDITsO7VOH3n0/3S5o9Lt9YN22MC
ArCvHegeNd2DR5WLbUBAvxgk7TqYYy2XnAkBnfRudu+LmL7mH6n40xCIB0yuuBTk
klZQCvWUi7EUdHie2beILVReHrLk8kdaZTflE6EingrR5LsBV7dka1warzMmYf16
TSDdthvFy0Li27NUk/PjTmzjuu1KtOs7j7FHc/i/UAMg2UA7s2x14SEM7b3UeCH8
kMnPNayGJx/jUhFxxfHHMCyPZhNdSIbKFtRkK9kqSSYZ1vzvtefe0PRbDiKz+MwU
pAx0VqJs6XtoRakINuDqm2ugrBPFSPdyA7pYnSAyl6pdb8UDkABzcai/ni4u1y2J
kQ2tBId2qT+3wGoe+dJ13eLKTRp691k4yOafJg/H7siLsXm+BW4jDHo91hz/ayUN
tz23y4rraKpa2b3DlK9bxvWbS/Lhpgi2xQcb0SwmYdHDgWj0EPHvJqXAgRs8lu6e
oXlD4D+o/DuZK2NeRQxysV9ST/qPzk+PEo23OOc3UOtW4O8SRKDnXjdorm0uS5kT
htYslYc0lRbcQgKk09QKDUP7AhHtc8YBC4O+ClHf7JehnHB/UoZDHZs42+OR7+lC
pqWiRGbWhww4Hxp+LxSsR+NNEnZ2mZJ8+xOahc/Gg+Yq/U0v/ujZa3NDnaldwYzQ
nHlK/qEloy+FlzbdSofS51L+Dpmn51WUskBKwgFC1QzUolc+LorG8nS4JG53+cqL
ArKLnQEyXsCvj87d38yRi/HmU3SZzVnajdLqERamqaS5b4Z6U/uS4vqZkGpITiqR
avSpT33FnV+P3GZEEHZKbAqbOfCIOt+xqxpmZKm1bQO4K+gsZpezmJ7tRo6djUtm
j+UT7H97QKh2/Qad7DEVLdi8SO1Z243RE51IqfD3BMOwnrLgb5BRx1x22pjmCjyr
7I/smRV9KLukUW3BPHMPYy5GPSyN5zjaDUOjrxC7jGJmx5H1s4203BhUmiZoA7s0
A9VPWObwq/rmgiF1DIUjRnPinsJrXm7Canp+VeIsXRCvov+sgj7U+//URu039UKa
z42m9VJYjUOxEm4u2v+qqllTFkDatzAPpVMrHSjWA80885gYg912+7dCyvU7uNfX
3Aqw1EVg1hiJUMbjZTMNWSDvbDdZzp3gcaVpVpeMXXPxff1HIH+A+9jLDt/C7aoL
Gny86al+oTij8jsZl/+g4zAvDNfiIZZhBzIDTcATbgl6wbVsWRYo6GCEGanKGiyl
OMFokNe/9GCol0ZxFdS5AHU6EMfefmlHMwxek3S8oaat0MYPLEcHbDo40rplZ0Jp
eCULyz/MrCdVE5pVgUaSCV7UjThWERP/BShgguB8avAvdHyVqhHfLdj7fHOrn1q/
dRJPgRsy3kox4DEn17tto83MwnPloEoItkAD3m6oJDZ07F3hsMUk10AhI1iJf58O
pUlxIKqpk/JdchHymmpiS8NwbrFR/B7gUvkNCyRi0PT93bf1K2v74M1Pf58Edc5T
FicFGqbtDeC8qJoIX1L8HIHqy6fEPwya2qRJrPdr92U5+msK9GcQdiQUwgGB+HmD
4NdHUDUN9MMJ0A3CbY98xSN7qsLA+phBKGwOG6l/PrIZj+s45jqXOzFE+9uiHd7C
hx0Iwpa11cF9Z3KxT8kDlccEAZVVnMoitvLXGTpH63j90NHU+jE8jf20bxgcSvGc
PATQiABpC5BWJ3KJxV5YyRoktkrMtIClpa8LIZB67mb3BSB/WYcVCp51lF9Zl+lN
yBW7p26Y6ZED2Bf45ltOzBRzbkOOPT6ZGg5mFTV0FPGdJ4hKjZKOFxbip+29OaBl
YUQqh+23IQuMkfUaZ463DzVEyKjCeebeGcwc9PZBK+BRCnJxjLQQ402qTUihWgqg
RghOHX6/eM6XR1XJE/spIzPHaaVz7mLIvYMWsdQY7wWf5b+MtMGAAoMXL4/gHkN5
LlTjzHep7JbV4V79v9w2uPcqUzKiS/CuQmEdZPW22V45oG8u0enwFNd/sTC9N5M8
fcoBX3Rwc9qtZCkGHYoUzC1Z4NGPouHE9Scx6GbhrtU38MQYC5QWQ+qFbB5wDYkR
GQm7JZEkctN13Uzp5HsFJK0UgQROoTtbU/l26EjRpXjQkIC+1RMuMf2Q0VFmV0mO
SdXzJ+JcEmhTSCuEGMMNs5jBtYQVtgsI8Cx3RbfErUVYX4T/aP5qgIso3sczbEqe
SGdWoDHUwMXIyjsopvSrW55LtA8Lr0jMsMzJ7VALsTAn4S7A046OhE4mYSLtSJwm
9CCP5eGY370mjrojPE5W64J2wUAImCkMkCBA5In9GiKM5gClRadlaVdsVdQ2MCMF
rTeL2fuPFDdgYL94I/ifb9GNnDe2vs9IwgHpJaniHK00ECxLqbxUJc0b994ikTSQ
elyL4iSSvTOu+M2CrafeQ9tiJ/2Jq3phytR9soN2B8GwqoYOoXsjPLCqtkvlvYeI
JNS6jcNqmdSWgrcIMErT2uZ8CHBIO6redYUpjCx2saKquNBYOHj+8ZFJG4jqoJCs
+NKAjSzmtWwK9fn3pqipgafz+I2zGEOYrovB8hB4klhWkLUFqK6u+NsjGdui/AHc
wrbB1jo7/Ym1Nvyh2BUyUYBDTMsd+KDmEZunUWOGxjtmtV49Mq8fA2sHNH/+7yNb
B2PW1k2RlEv5MtLHPfL1j+0oVpObX/iAEy1eZIIAETBNyAcceKG+5oon/H2mu6eS
U5V6rRJRzdXlA4UODwHqxyLIYa0npuMqfPkGxTZpes6qV4CPfAYtDHPMrkKd+Xd9
B5uqepmBmaER83OeodAH5xc++nhewDBLhTkE7iVq8DyJNcS2RgsSTiiWINt9jQhw
r2w/rFn8BcgWukEfS4EkvD5XfjdQRpVVTKkorxWHzgE6X/z0ki58f2DazNxAVOq5
5HHtK4wnMRqYs0uMlr2s/Th5Qfv06cP5+tcULB79E4q/NGEva1z0z2HbfPHiNDYc
4CHhcnQQfqdF86HGST9yDGEdcIFNRm6D89MjtT3JWq/lZMNkHthO7Jk4vWA7INOm
SXyRdiXotCBINgAjb8z1scypLEpRFioTx/tK8nVKnZR637RlyIv2LjTMFMsF+kJy
BDzY+3guIOjEuW08i+hqWgEeSZwHHLXO6kRjxiHDiYGbzLLHX5/Hp7EbNfJ7kNWd
oZQF+IQgrCRFri1F89Fp3ti857oIsCj4OGncQashXL4Cx1zp3+zawkC2fH+RESmx
wZityJUif1TZs07no4bLR1qssorUSVkDF4QuIvF2PTr9PQ0V4vx4JZYq4hpXIoRi
16JjM2PQRSWuX5ttJVWOckcLHpaGxHjYsI1AOV5bWIa+S2vy9PDszSyAv0Do0kKn
3HBkaU37kSucRf3zXdlt6hZW3l2W4IIQF6/FMwm4u54DVIyBbJWlsjuz2b/NHYPH
v/knRqAgC7XWkGYdnHXQFNcOd7Mbes5B3dS9DJKhCfrtr5OEc51YsGFlSzhtXai8
SF1Qpci1VxTE9wgGeTrKNPIvgaXhzsS2F9fBE1+UT/Xin8Cg8H+VxTweAbp/z35L
WpGbKyuTeHDiMfxr7CrfY5wjS43E3+j8Qtcu9lAjTxS+jnhROb7qLt/Eq0qqX4jR
7Cd3ZCekDQnJnXU4x08sSk+WxO1OdIklcG8mErIxKekbjmsH+/S/AdpCih2lhYVu
bZt0x/i4l/LazTrjKQuFoCKSN0W9Iif4J/m7iXJeYfz/3Dbgu6C055jS0M5A0Ckc
V3cJ+MvxevJtt01XWoBvbNNnCkpMie7vUHtrj0Y6Sw3WlkUsCCNbg/ky36hKUyjA
d716wr7Kq8x1hOnp+8StIBYsRfSbVVQw8D3iR7U2HfOlWfj8VaEUX0Mk2J6qyls3
h/kAxffvSAf0wn2KeGZaCqU03BGuOJ+pm94AaFRvigkZ7YzUaT41pG29GpFg7UYH
UV7O0bmpOI+mg9qoo5RGJqo4q1Ia2pv27cI4hs3COvqFeQzx5+uY2JEKNrHCeMbd
Qqlf9SZzxoKkQ5dYlKIqb51LRo9hpiKLF5EteDYTjQEzTuzupbbeKhxvwt2pAajF
sltUEbTcGOHzUtCgNKwp5QTKCkwR1NaD+ca6m13FvZgCx6YtuZCDExgE/1sHNWaS
11W8Akh22GsYavqhtY5mAPY9pROmOr74XjF/ltEykb2hf9rb/Zyr3fH+9YczYwFX
b6a0StSgnJdHHM6KPhBEWjehfwsjMvrR3YQNSisrnw6lpFlJCyLr/C8ruDnEmXAR
54mCV2S7uXzKG3ZP5z1SFp2wij/7dSC7Hf2q9TRZY1rnM1sxhdDuaLKmA0soP66X
VDp5o8JQ+yHL4VsWqbYo+Q36QihRCz9u6DG0N7YAv1N4KaiZT/NXgIJvd3NN0fhr
eBAOtMFBPb78H+OmjIx1BiyJSQgE/ZuFmf2BnfipouJ2C1sCdxZw1Nh4nVjXcnlT
PA0VLp0XT6v1156+Zyz4KJwqlikehRrXqi+k+TRba15PJnWzGl4ix5qcARTtHK6H
FkxLL6RFu7mWjPZChcRSrj8XVHiK6w+S2KgdHNJtuOnJw6wtYN9pmjemXfQiwNl6
ENy4TisiSMj2wz8IIx+f/rbQ3rrsviO6nQ4iaE7yWtZpLcnbdXXClVYaR+pySSBo
NasGfh4Edaqto3oFPnyx2MA4bWYIR7gx4zqD6uN+wGHz9Lrop8n6wAsDkWmdgD64
S9cpw5A4z6xWBMbqfsFxMRluZL33QQdGnRLQ+yAniZaa/PW5jFN70oopgi4MVe6P
/aCgdU4nnSJvAznBfCW1x05Hj/o09ErhDb5sECA/WxWGHhzKU9RsshXXlymREuym
F/Nu9envPurDuQp3O4x05U6bOaiSgrHPLLxTpPUXcQTImYF3khbeWxhhi8Bcsv6O
hbWYJ5TBmxjBIFKfgcGYwnSgorBHEOJ2VzrG6urRKZn0RGXoxkeHjpxzSYiNtQhC
E0BQPZXkHNZm0ERH+i9IRKjKONVgAI9ye0vvqd+uXvrkrMvQnucxSl8GadZwDSdd
i42dPuxoii/dpS+231pREoLetbGqSlYnGGazlPVlXJTRt5Q9PSOxMjX0yjaYa4vH
i3vEFOUn/aWmGQW87BatMmrWsXoFhCHBI330QwSzyZ1qhQvrw8y69xvUfZk6TxGZ
U6zVlZ2a5Y99a8qvZTjkNi115z42KQuAUo99+kkXTrIgLZcBhjmkKoYPckCE5LrG
aDLBW9kCrWT6RU2e0o8l6O3GsiHqfYJFnD2CDiWDiidjSYFKAMM+bBq9x7C0WgkS
2RLrPb44UzM0sNaww/800O94+XN5PSPMXybw0C+DUbdkFnEk5hq/Bv/XpFYt6htr
OMLoElVBTWnN0epYWYUodgYsIYY+dOjLBJv+3lrIxwrFJAGn9B90LkxM/jpNM31L
KHUEcTEEtwNLrCecpE4a65QmOv+4/Y4tOurU6pG7WDiFC1MbOLDWCNdE9/jx+He+
+wAgimv+IrLOhfkGbb+UgXS7gbkFFywbQHL833qpCsvUWpUiXyr3Yn7rvHHfbXlT
VOIrnK+bpNkt1Pe0TldnKvKnWMtaf+LqunsSFdEmWas/HhMWoujJ0fXlyk5d6TSg
K9DI44aLqM+kAgOiYA2zk++NHA6cJWE+KrfMlBR1Sjfwzq4xwrzU4uZ4Jz3E80Lc
HCiABqcZxXjAU6gqzjC3uErgkIjYO4jPiZSkInxuZkqQkg+VNDd9g2/9OrC7OpUL
w48kZTJNyOkXdfO+bMBdF+duCNzqhw3YF3lOELtmaq9/LDzgg1h1IGH6GPqfk5hO
ljT1Rs0nn6ppKHlzq/kcZAEBvz/9JqxLvh0GT5sUl44YVwuhO0Joa2Ihmwx2EXMK
BLml+AB4MFw2ENl2rPhChWxwOINm5ABA1B2h3VKVOTdMTfVdxlb27Js7WIeQbX8S
/aMpaq79+ui4oxPoet4WRzVjGZyBYDynPvP021v9RSJf5m1+6gxAwEHHNlNIzdpb
zkRulrGX5AW4cqOLIiycXJlklu8M4+KA+j0iNQAGugQ0WKV1jTmnl00EbPcZGXGt
hQS1f1XDT+PLgEhU9XIV7kyGG14NQZwIuiqWhcY1HO6gwMSL6nlfjq/bgvqCax0o
CoLD+3og9dITGPhpleQAm5k/N68oEfJZhVuVjIvvJxe/HZSyKBu9xWkjKCQVd9kI
5sV7yXUn0n9AgQgp1osfXF4vpvCeRTWyrFyd8noP6MSAXb/Lbv0VSRGO+54lN+Fe
xAzx1re7ZXTcvsK6sIH4cseTMJlgGsI2/oQJ/0/eRXavNINldwduVSN1XMWrsvyE
cj5YeDJen//ceMFCE6Qc+rfHCLa7yqWk0B3WvSrItW7/sXzf8rUGzAIfUt/UO/HZ
JAn7rjzXYvv+QplQnLbkdI8uL6eTxMNZ1m1EzHYzdmUxusUmLep5nrRsGYCWi7Uc
KUp5sIVoIfESrfrEZW6MfgBT2cDpbNHZrEt8nPogjsW4+42iayC8b9ki8sc5CX6j
GXSHLn393B/94gOlINiBRgLcLbrFmTGp8P8ToKXZ/iXsaEHV42UXoNlrDhb03xan
3RStyGyHlD5ux5LnUIQ7gDGvhNwo0Qwhb1uUs1REYk1MDgXbgW54EQTc4pJEelnA
HmJy477JxrP00cCDzVZ8ykvERrT4YlyHK3iExvlpmU+XLuRx2e+bGRB3ed6I5kMP
Dh3Ytal3CAjMpj4/7C6FBkzum51DHTb6mWEF4w4ApxkaQWZPOuOSX36xHNHf3+i3
BoVlQILVyqgaBd3HwypcuPmhno3hfxvrL7HbLprOL0GfnnRlCqOxlgyDw2E2NK2o
Vr0Cx+4qZy68AuRNi2R4janc37R2DyO3W+jYyKtL0JOwrGhOgjMhQmYGxXFo2VVR
kHP1uRfvOWI2ZxXXuVQzo7H3RnhebAuVFLIM+IQPWuBqIHVh/rNFXbhe2N0iMnOn
xDMwjIx2wEoGqFZNNK2aGdS9kJdtUTyAX3UovM/hgTYStggAYUUx4vOEyb4pAakp
/QUMCiedqUrRvhyNi1xd2IkgEXX2gQDcXcCrv/CQMO4GeBD+ocWO3ozhVP/Rmv2S
OhNjNW1r4xakR43mKtmN9kMXxi/Su0LmPkPnPOtJDueLYtiGlYqeFVxCfmkm8oSc
NEhPVBLKL8H6hvZYOVtf2ehxd3l6nbWqjzVIqnCY1/4IDNUQvFihNa2L8ay4ziqE
mJ/uboOXCfoH0QP1pgiCJYYnaSXSRwVdeq7bl40HQvq35LO8XUMyub+XLvrKW13y
Xw+i8Tf7P8Vntc4USRUzZoTwCEfMtP0eKtyqjuFzTCkAzmLFlkc1bjxDDi+ZOSBr
TXo6wG5CAQhgwz5+LWsgFCpET1ouwj6I/fPmocW49DbGOmsohAEllOuIA+opaDuV
+Q4QpK+nijAm1XTQpPPlDCdVIVlAEBFmg7FH/WyG9UMMyaw+/4bcF9ldPRix52Z/
G3Z8lUrp1ex024ZB10yPJG4/ZxZENviyAnaqln7FKVh6FIQpcZjNpqYVHJnb7o55
/5joCBiQ5lr/qobxSjL9wFSh8eyMXZOOGteBJn1aK41oelsGfIEbxDbPVwwbleal
1m4bLi+wE0x4cuDjyBRzsTZCcdJPOFV4oq+wZYXr43eYqonn/AA8FbDiizje6EtO
3Wy13KrOwzJs25wzm86pHxYADv6YT/1OirZDGXw9vPIK3mDPhwBP9cICpxq7+rdM
3AWuhPXiITIDqv17vYCFiE4RsjJL9VwRCdoJKJrfm+PmxWwh9LHysvZvnGqU1PgD
8vFV3MJEJiy2Vau9FobZSjab+i6GsrWXQmsniiL/lbauBdm5CwyEPFDxdfopXK1g
p3dXUtoUJNuopDZOxSiaaZgoUivi4nxFqHZQXpIFbJ22u53U4CV1zfQstGAgfTxT
IiWvI3emKtaFRQCB7f875Gy9WoQxNsEpTY8GYYe/e3xLrXT2X7uygH3viXEKwQsi
W1mncWoqTpFMlyExsHXC7Jor/PBav200PaJugckZAKuH/5aV5mnoj6LM/Kd3XaHG
DPU+0bURqvBtc16FDN8qBPN2YkXIFoN/3ilOzmFp7B8h8axy6E/rfE0Npbjg4DLi
U/aMuz9ddQdmbhVRTSg8ZL4SZbhimOlsVTPqcu9qMGi2QR1MRGU/rcQW+QbwvWSd
Ic2QlKJNwO6HEgZjmLqbtpRE06RGp21Cv9of6aZ7nHK0MOkUALoQwmpBscJhxuwa
lJU6al1/paa5fRbL8/O3X3iTcmx/9rwkDROKy0ZwWuTQzod62jzTeYiPEHOlD3qJ
oYHb/nKDywUwKTXikzMILFsjvm46H0UqDemczB7xdlWLscufQFjeoJlOWhwPFiEd
31G4kDgUnIfd4InIt5R+HjoLPKj0ynhOqVdipA4+dgGdMwYINJK+ueisctp1mGJ3
fRV4gC+rCYtXWt8b83BNlkcJ43jpSna2/VI4cbaLL3iyHfxot9TwgSHH3KtSSPUK
W9V2VxWoz4uLr9qWtohdHB9r5wOymyT5DnKXHEeU7IbNya0v94jrm5tY7oHBDMBu
2rTPoCLEO9AGni20DtIZ47ogueBJvOIuxpWiZIMqtyNHh1K1Z2nbsOH96fwo19yU
l2q06aArcVeR6zHIih1AiNV2xpWWRdMt4jaYIOu2lD3PNuGKXjSV5BkStrr5TqjB
VDZMDyu/DhkMhZKILz+L3pXBmMUkiv4P1mZUw6RgjyZc0boWxsrHbODuMuv0bxm/
7KcB6X1/EF52X2Zf47S3b7zco7RxNfc2vvxd+sFSYonTBcMJpdJJ9Uv3C6qCeMUd
W9P5GaedK4VTgYW7jVAH/K3Z8zenNjDDevyQJlKU7iFTLwsftZJxryylxMw0ULmU
PdtQ4i+rwRkZb7hIEvdlMh7u9LinA29NZhMdem4ZZs1oI0Cdq7chLQtc6dhlfKiG
hQzQoxOJXlX2YHQZHXkSH7zUpMN9N5dBFXxMjnKQ84L0gttEbDr9+RQWJmLQ7VNn
ic3plTQRyWStUftbqf4BhRwigxQ8OLr4lR4rwpdg2qm/XRltW6gCLS2xgJLAryhq
w6IlgLSVvhxu3cZKboOR/EB2WjJ89TgXJl6ZXOvRCb7fnVbHasneXubGnxyuToPg
WeRK9KrBHxnLZIv5GwF+DJKRmOIePG7Fki/XxgzDlHCM1GMq3hmR8xAG/fo8FNZH
1IzQCdPku4sLxszhC0/L2QB1WyhNbiYaI8+nfXq/eZxCiE4LZau9ePtRKyFiVYzM
CLdhziao/fOFFqd4PHJJU0LthKxyb09qEljo5PMkN7r35Q7lK/CTLxdN4GaH34RI
6Sx9rPaycoD/0M0Y7uxOzBdS9aFdfguzhATxtjpCrXqwknLyga71oQgY2yPdnx+B
Ku4/MaTmtMnDLpW2YfMzfxzJ5TBPa+lG688xzsNfqA5glqSEIPTw1wQqSM9AqEBn
FBtJri8uZ+wZUkUMger/8yxnWVQGxAXKQzgjzE+4jsquV/Qo99vU5Cn6/xx8nMK/
1kQTIFSgwWN4XZypzQGH2P8MGgv9cksw1HBv86YH/QBOuc0MrbTliMPrsGhkN7By
TDTIB29iQxX91rUFHeYCPQzjik1+pQNXfAAj8F5dakCnbBazto2DbYiIXRPa1xTZ
/Ou26jtrixQKiCUWlWdgmKJS/FpbQ+wutxjn/eaCP2x5d5KUjKiUqhQlsBj5E/6Y
Ukvu3KcFGgAod9X/klz9QVS9OMlWwwFHVtFMqv0Jt4RMLxib5lqsumcz3Ya9TX6g
opWOfph+OYXeLayGa4YGevNuZFA+TPWh8gNha+tqovteJAAS4yoiPJBGlGZSP42K
8qdK/ijLDosKRV87nvqa5L23fGV+5VCGtFZEVi75FzIgNpaB+uR39r+O5RmCQjjd
9UTSdbRIVR12MaTyojT507TMU4E6e7yJjpLu0uj4igq10aTCpdSuQFqWLDBS3YIc
7U7MUq8DhGDGPJizjHPy0lp+mwbCPKQ7wid9x3tfAD+iBIobe4KX49AWlrcARajy
3jPldzUUubaXNPSw9A9VhZwFAuD0OCtVV/4N+WO23KXz/ay7sICiJMxuB9Q9rkfZ
O2s6aceqyu6h7rlHFuXrvD9PAWCmzYwxMPQMwHpnMJK4j4bJTcHpcOZxdeO73VYo
2Jh5ZB3wEZT67RcKOHJXuV75ccMh1xUDg72rzYS4aHEsCDe4wVNhcbsVRVKIrpl6
vt5LiL5M5wi5jHtf/UtiBeIGYUVIfeSvZmqql5NSqeLVvPhOxn/tos6mKIw1VG/V
LsC186hLTPxMNsaeLy15tMvU4ku/qNTPeFC/2+odF4Ews3nCD90oYDUfi9FHE/UO
WWhce/fJhrBr1dcHRT7uQw0FKmJGQTnjB/PaHcocSJPoC2L+fOaTYRotVJyQIO89
EZ1QfYavyANr9qGD1g4z7DP1Tjt5aw273bZAKngEubXLbedmdVdy9ry4tb+cx/Ki
w3HS5inz9QGxdJuxlYygAKJxalkWUEwMAxJOdzprKqtfopRLIOWlXFseumM6FDFM
cMBYYVAcXkBqNLCzZKbVip+JBX2hN6kngk/YQhjHgnPvFvGGWUPYPLsoiQDo99Lv
kAPhkqVpRb+PMxWc2YOudRtj/GHWjIGNWFlsuiXyJ6mHNI9UDH6q3l4hNzXE96gd
mBkNrv6MNlugFy3cqEeMhojX/cVMaoXQTZD1Gpp3TKGVYZDiSjcTuRHawJ5b/DeE
gWq0RPwzhgLrcmfnTpZ1mxXX4gcwlQAm0WIu2uA/Ov/64iV2ijImccgK1/A8rQMO
A8uqFRh/k+bHsmoCkAI8mm8UJz/R17UopgTRqmiCKW1eZjqWIA2U69dPThost/sN
1Cl7qaKVpSWWxG5o5TvXOpd0S0/Ayvso7TserAOxffVB9va4xteECQ/bNMj2ac9a
ppT+ooQ+7ugv9wxejuyARMU4cghy7r4916o5nMHpAFtGf+rIgCGWr4cqDiIuM15t
uRkSF9uqEZR+/skbEV9rKXXcZyilBCJ3wmz6ZQqJR1cVfb5hrZZslAYc+6O5wWkK
O9vjhDYrAEpkeKIx2lRMAE83qq3iWKO6cs4ohSxp1SdK7cTH5QF0bpjWelihz/W2
heIndnC9lMY+Rft4CeE+AvxjkZhJHpEn32HEN0LcBd6ZdEVDuMp8T2hh6PQgBBaA
0FvbceS7ty8j1G9lfZiTxGhqbB3wL/PVqjIsQ5Mlb7mOBA4MzAXNYBXhYgHHdT9e
LfGLj8P/ta+Hr6k2+Aw4os+CUTOwbZOvW7HIafLgwSTOEKlNLg0SSG0WVQWMoxoz
9K6jxO+z1U9qF0MQNK9cdWGHgSZao68oYwWUUdWxc2U2F8yOE+d3/s6S58n/JXxB
awT5ov7Zk6TA57xfnDtgniVJVYqWXqjP3weEoxhBks+i3hPCJ2i6Sn9k8jb25sUp
O8tkcaCnY9Taw6koJZD5sIzOAyMHNSWs4h7lzu7TYBOt9OzOh9x3hl5siEFaZ1xI
TF75g4+rS33v938C7sCsmvATHHPDbnYReiV6i9+7rdSZg7u3CuEjcAFXV3W+JdUt
nOwjYl+sHBUS1DjXug01KXSNlm6TOQpODnmPImDVeh6VArAnwQnaJ3T5UfaTOg/8
gIKzzC9UjL1n46uyVW4Lized5SVyVCkXEQ3RO5g12qaxzzCCm+I1IHV/Oz9TpKqe
CtP6GGTfP2Qb9+xMmPM3yIp9W4qyGeFmtCjPGHvgbL4er3bdiCNaNBPv7meY/geE
dyKH7WxvVReTF123zfMQafyX7JiMzzIo7SIGpP1DZ7ywyKxKlv8YhStA0hsWjzpo
kjKOAsx8SVHLAUeRFOq0191Yg+VoGm8e7PrYpUBAtVC5kyeqEL3QkqC279ShpZkE
lYrulNntcw9Ntai533XSOj23g2Tzp+dVUMyEpftqefsuba9Tg13/PtjDyK7WoH7Q
jSCe62P5kdkI7fqY0WmnqV2HZJvHUJzwdidMW6xgFYyZb6D8mRShWIkpwh00+mmS
nT6LFp4Pjgqe+JY3+8ZPxu781A1DrgWMi459Aod/0OHbbiVhoi7MUFEhwKUsUFiJ
eTActXAL1HxmzKo+PYwQbTLbj+uOJl+i4YMwoa0bMzHYIoEf73mfZ87aqUEB89V4
0r4hfXvKGvgOXcjkZX+b2xOI+9/Zp4DkkZoB1NRjEqLUY5K8s88MmO2kE4V6ScxZ
EyP4kntDBUUzPkHcXpb4VZ/Wm0snf7czuwSfpbXOBgVXWXOqI+KDvAeM/eFLJzbM
J81q26awOQsnD1XhnJz7N3XXNXy9wNfA5iWCcY9MwTxHs7OgPCiuh/IDQGkDiArd
TCoVilz7MX0uH5OLx2ZJCVjwHXbp61D5o6/Ke3CBs1WvI8Wes0KLE7uxHtjflYyr
TbnsIv7HLxYF7LCrpnjgsLmqICi4xHmwQoBQwLs4Ga9mqLZIYN0Jvxisu9/IE8Hz
jqNgCCsngx7pB1ONX2PWjbJM3PKwlH1/sSsezU0nc1pBJeXZvXalhv4KBKMbYLhk
rXClwFEpYh9BVMIv+0jnHZOQxSaqKynY7zR7zZ7iGRWnMkZMfTkUk3mQYc/P4mAh
7Bv4XnhVIPA3z5iidguldnrw72uiMYf5tLArMZ1zCMMufROwmywE27Taj5jGKkwt
Iw27673eWlgxsNvsZFl/t9v1/BtC0j+DCu0pETB11657m3EvNf6Sjc+oBS5nxj22
bbIW+cgJOivsmFCUHqpD0CJqiMFM1XSr9rQrfQwLvUrRc9UjGox+m8ArFYifIRCX
mm97jjHp8gSw4zyzUZniSk/j3eNxGVXzFM/vIYkrJpYSMuxYc80UILB0velltZMr
VnfuwiUGWoQYcj40pj5vNyAsB7bsP2NLnAExz4kPpjP1UpI1auSmw8nmh70hGzEn
aAY+klqRJfH9kXRirUK+EWqj3LjfqtXU7G+JlwmFvc0mCVBp7u1YrrQoEKlvOgiN
8Xw/r54x+FuaLu67MkXAZk+HPB4JMU2SK9uvuywhkPGphyux1LUHNbmyoJ4B558O
sNJr46tsX4V3qkOv/6gm6hgXbWzF2AHvPx8G5WOsvYSwFAHaXerW90DpieCvQVfK
TgBJ0r3CiUvA0Q87WQ8L2dD1N/gcv2XOkTSC7VDBYaNMayAWa/U4hnsx9VMoCRMP
iLFrm039+NxO52MHch4dPd6SGEOXhGvIfPxQlbPsFIY6XttMeK2I0Zv9mY0fhgbe
LrExdLdwPWwszzBagug+cQrFOpsH8+G68O+l264C5etmRzOmYY80pdWgnOqX/nUx
OxUAPSJVn//BGnL9t350YUIwCicpXQe+I1RttjEr1nq8Jv5wCdYP/sNLXPt2UYUu
tHtdo98V6nds+lm4A1zak6tuxiEoxRlzHGh1Ytb+D5gQrvMxX/ZaiWJHOf2Z6cuD
Aw8QtY47TITiIhnX45FcwDlXbl6CIFMX+DCOd1URdgmnnviu5Kf44SmcopbL+ZS5
rZ/PgUIVyTjG5Ue+OIGmR9dwXWuM+auTiFqCD6F2FuSV3fu57hxqsODqJJdJG1hI
TS81MwXFaTXwCPN80eLuh/zu1lAVnSS9r9dtvV/tccbllRxVy8mYVTLe50Z593q9
CE8M56UANWe1od5f64ze85fW07MRjKNDrWxSZHs2y80JfRcBgxBcWorAr2EopmuI
R/9+nUoOMl3Q2lDhF687iGaKigrj5Md2hCWgkdrOuPJFs53LgjQglIzl6nTjzTNR
GKdhzm8cOkxj9OjnUvJVgRxfTUWWyyZlDRsYRooKAWQns2+ARiXVgS02tYVJTR3m
K3kZOg9A8XW3nUqo36wPW9YE8C9Ym69K3TKFX6mX+KrP9fZpiSRyyiT9O9CDDBoS
HNDyHKitX7CQNK7WVxwGeuEHXGvg3DwxLazyz/0/HjFCgqcPrfelOpKHrbBCFAoi
bEzSpo3ePC3uXGhxyyykIhTtNZfgi2IO12eRfGnv3nSr3hnwN2T0ufFkDEFI2UVM
rGujMK2PPV1gHCZ1T3vZd2ZR5B9flJulJaK28gO+P8rHNMO0Rqz4vfdltWI9/Mqu
k42FL7rDgZTQBYLKImsp3CPW9md4YfKOOqUFOxdj7Timbgi31TCNgZFvXNWsYjcX
0iyz+2PEd9rpx7BaxvGORH5KMP9uQZTkiVS8Q8II2JcoJv3t2lFIEXnMGhIjo9L7
RTHXfeH2YBmEIWtC1TYHQUsFOTFuTAhZApOlVT5xDR9LMviF8KSa1hoVwCP9d6pJ
YnBfAYnEnjHHme6iPCqi7WaB2TUFzbA8Dy9hgIq/wrum2RNasgB5qCG5DO/Mjpob
hCmPNjIt3sevpgyttyb/QSTt+b6wgIkRl8ON1CZco/su7xhKdkZDM9yVVxUcprln
mibE3MaPqA/gK2fHYdcwXl/rEuKg+NhZzL0wfl4G1zyPPARKJcwsUQ2nv2Tje0nS
WOJBz34pAf2Ztcj9kZ2mJ2ZL067dVPB/P0z90CzgZRY64w68xLHvZumqU9BX0fKg
rYB0isLJ5dVYMm3Da/5RNzgcigLZu8q5pYV0V+9eKGT/3e2yF4NPYYGflXp2OYgt
MmZOINDCYd5BNOdEH+4EJCWY1SYjQpkZeFg+bNODpwObPVSgt+G4igwStcTc6G1t
ie30tm2KOfYM1qeEBKOXREi0tLPsLvkbEak5AXK0XCis/vTmDDVo/5LJmQhc64/z
clVR5s+J0dLC5BdoolNZ/fOFKQvsPDBja9o69zSGVR1mcDeA86Pv1hHNKcZe17a8
vPc7fE7XZ5yOZFPtHjKiGBWVvFRH1D8RE+gJa4cIsPwbJLJ1vQO9fjFCpII6QAUn
tOL8LqSe61cy2qb2fzXeeRdbRnSt3eXQsNtKlLjmxVUUxFKPZhwz9CZOYAsOL1x9
U+zSw7QVaoclMmXJIXbEfWeSveC9XeXGfQd/nn9Bx1jJmmx7oOGkAEr2q59x+0Tk
bN6BuPYWlKX3EtrkHKcIUK51CDTuMmM2OC7MYUfNly5ecO3aEEe1kxrz7tYHkAx2
dn2KvWLePJMWfiGP7UaMznM4V239WcpEgCtvDcNTYn4QAmDFAdP2g7BOuRXOQJrz
OPad+PhpEHgr5SvFWYTBaRzyrmIwJrstsZKLME58/q20m4UKiIhhJRycguV3yHKo
xK+1JSiH+w6HIY446TLWfdbFVohtR9li4uwRLVhA95n6NzDmdM2SiPs3dHH37s50
yWOTZc4cGHMXL0Ddc7VUNS3BGX+qlTQzkPTEqedGVXAANua6USF0f0F03lpQTYkY
nlcvXgv+3GNRA2IcewLyEqZM6u7GmD4rQUqYmAf8+6Gm2nj2e1Sc0RqyQihysX6s
DbXD0YuH+7qG6eorAmYDFHXJpomuxKSTnS4a78RNq+TkcIFoVIxpbOj+YLNhjo/N
UhVrqDtmyG0G018NRRtGd9U/HJtBtx91t9pbkfL/pe/JYfVV5daJgRkuze0XvzXE
nfHFKCgTNkqN4xrtZfhaA2X2II+YKkSOj4OKjb12QJ7omVYuypbQoGjAdM+SUclQ
mo+Bd6ChC9+HxAMMjLcd4MZRwggK2S/c2VOk3qJbx/htDoZRBFXvoBcvGC4O70sU
eOFB+tu4TWx4rbGziUAHNUeMWOpFjr3xDMR0g+vepPhVOvlYC3SnMI1KTUVdzw7a
EATuyt8imu/vcZCaUHT6leXduwfURHGFhLq/wffHIHSbi0+4eR7bF/KcWdFv79h+
TqoYQz76KAFlrrtKkMTbMXJcjrL8IfvxjTghj7hpI+r9XZ5uQlQgLiaER6oYJTvn
HBIvNLKCNnzBn1u1zdBu05yBsDYzQbxMI8kjg2qZkhVes5wO5rlVIfdRLClnVMct
50MTPDVkp+N0Ab7AhDw+H6FFABMeGUZQTLfqXB3U1n2G84/2Lr5GCK3wt9wb5MAA
ebp2LXeUPCNetA4EWsG86d178/uzYvyA0u0Xv4XFJbRKqM4O6Bhsl4QKSJL2JZOy
IB0o6m17HPtL+uHOL+h7LyHrKwDGAFR1tAY/XyczTvd6cSfefy92byhr8n+npTQX
2ME9D3Xnxk+voFSmbhin7cA4jxAS9ut+WTTvOTqSBkKFsUlxG3mTP/5ukSg0L52S
RbcTvgVtluJfVU1s+35483KBbHWDuzaKTGiR225bUK92U+jAVfudyA7FIgBtVIqH
RizG6FBGGW+FbSZwMrgoENTCnEhLz4Fy5TfqsDXWWOtgTZGWiZnG18XRCnw2qquP
MJxItfq979OanIwX8WconWp2GtN4hHK4cguoV+yhvcstHlPcEakYbGtrCN9UQrvi
JLGrN8lObgvmJ4ARPbIJBysQppt/MQodEO0ZNBa3IXBBtz1VgZWxfLSE3Cdf6BW6
YeqRXlyxNsugfHZB5v2vJjaYKmMevc8wWVbltxN6Q99YJCy08+ZFPP7UUR20EDsr
0+sUsCHoTK0AulQ1JbQrD19bSgo/XUD9rgdTVM/vQ93Wm6ZY44thxnB7xQYtsgJb
gNzcDKxjqSvIu4unaUmFVRYyNKaHCtCxYMizCOeS4sLcAYG4puRLytkzXjSthrVF
fpmC03M+3JfRS1Rer5i8Yiczmwf11kcEgxznX5Er6g1g50WPa4Set1ntOeBLbWXw
//fwLUJCLif+TnU7TgKzsctgsZis9pY5W3JzPoOCuVoyZRCERaHcSy5rmFzXu2ZH
SA0cI9zFDgE3bzM+5mwrojcvfGWunqJsq2VxJtKpPZksFvqn99dENl8BtnkTBa+d
M9aEyVHjLI1xaKLnixDBviRYFwR/TdC41Jnfw5CKjgVOOvgMkRCseKx8tT9Zj7AM
aDaBkqYQfIzYoGvWHIB1G1Dbnarp7DmLo9OuE/uDuXLjL27BxY1g9556jQxqFGkx
jQxpLj0yHfhUefPycYnWFbYCObr8m70zrwCsD6//HQHtTeeLCRCz5YiAJt4Z3386
BMWogMpG2lHdfoKk9zyM8Gqvt47h/WCZD7Fct+Cm0QnrmeZB6aTcyYVxIHnDeh4N
peB0Sj+SYOBxLoyt09oJyk1XlJyKNvANlY3jc783UO2hBJUMKOQ0CXyshauBbFSy
tQJETd6xyU/hXwifrZKWYkz605XSIULwiWSDNCW2vtB3Gs9aqN9LTzHLHNro7fik
Y+xzx7OQTO/D7/7NDk51P8U+t+wRumaJJ7ntYYTgOf0HgoGig9sk3ZyFf6+ci3Rz
1KytkUecZYJxTIA8QcN548Zk8IsrK5H6to6+7foHbAsmjEs90JFbgIz5EBWHErrm
SgaL6Y1H9+UJZcP+6SCxX4V+mbrLk666b78hvVOcq2uCiRtfcDQb0Oj6zxU6Bva6
l9GsYNSQXGoZyj8J5HgWfs5rj+2KP/f8sGtMM7DjDrV6XONzgCp/EnuxLhlfIcbT
rloPI9kdUf03IWgVldqQZNzErHsG/RsJmytSyPPMtuCjWzRAqzqYXVJIeprEwdrl
YUeLvKuD8w6DIIMnAaBJNmQfKdL09jHBoGy/vvI0CJ2sVnjiTixee9avLBWkevrO
AbGuW6TK8zpCxDnK8DINBvv2Bca4YmQu4NQghE0FQrDrNbav4aXuxDWGMaJMdKYV
4cG8KtAUIZRXveNrBhHUTR4VEYLoAytt6OU4HgHW5r5Z0KYIqDoVlzVnoQloFXdW
+DwLN+Flx2oVnYIaRo1ZV4Bd20Lp7GmzcIwB45RrpkP17oJR0MkfAO8wV7VK7Fha
hZ012PIkh/oIzeTFPPilkL+ixs+QhhHUjiZNKPF3/1EsN3DN7Mf/4gioDHsNxvmj
s7Xjn8M/4dN+dgRZ4S7uRtvIjzgj2GWfFhXoW8nNad05PRI/BWJISeWYACTWzs6I
SHkLfA8ce8X+/nLaV09OEd6lundagp/xHno4BLkH4lVQppHO+E958LoMdY6MywMm
JTfMBmlCmjMINVZb9T+UNhuMCnq0Ntn0JrAsAYFQnnbbjp7oCQir8/Fy3lSnwgfP
+mpD2uK2yceEQXNfBcOoz5Ijeg91j9fZf5zIB/cbxZ++sbcvEUyQf+eYDziOSzMS
aguq6cPb+BezbY16Rcnz5Kx1wd5ETLzItK3+gSYYmvcdXdqi4zhiLzQ9JiuNXy6u
wAwHxVMsG1OTcB3Z/Z/3hcLqL/Wf00Pv2M5mYMOTg9XtbN+YU3K/vrzBQbJ9WlIe
oQOjjry4uKVbywDQchm6WnBAjpII63wInjYPeeQMkvt8swibLrEBM/l9YK+9KWYY
kU3T77IsJuRDC0msmgLW8zTjAmEaZMMP6BxMXrUZD0xqX1m/1C+KbNm92k9H/qNn
OgNhWw7oiIvhzZ1xku+J4EHd6E7jLo1Dhd85Pzw3y9kvNDm0idY60eAhmMyTuq3u
HALpJ0XnCuQlgqbPpNW545qaComir9sYiCfWdicHIKqWXjSMx0j6OMQiy4nETjRI
y8DTvSCscCZ0d22nU4o5efJ2q7X+EKGDvGUV9r3HaXWqQvZE+Y+d6YMgM1Vmp2fh
cb9n12L7FTe6EjkaqPpHEzRFCIpe/+Jmb0KB6LLH5LLRfliIFkhE3M6aNsHlqIz4
LJDDbB1YUh+Oy2Uz3ay+g9WyVgJQyefNH+oTbhcNwE6uKxeJoY3JoJ2cSh7c9Qz9
19mfc+8QCNjJWQvEWUfjieDVpbPUTzPhvIOnJEgCkb/Al8sNbd56kdlXT+VAmN76
v6Ho1VzZJvYB/Lk+GFkUmQqgXopgPRGVJmBWPNCVn0L2pWaCoaayIm/raczw+gnL
20kw8cep4q+qLI+qoYhIHjeG6f3+hHe9UfrB/hE+aIY160p05j3A/zstoFsMOw0v
GUKpN/1agKGld2Twl906J5wBnwcs2hOlEWx09UUvmUgpyhvQkYKI6gIRsk0EeITf
CljGVbJ8rFqEXD5lAWmSG/Pke1j3H2qQAjyiIv9J1nEv2n3tja1P3BgQRl46081b
nokuPHEu8bDfUK5ndp52Za7OvTXqM3l+cGbEx0wvbZUQr4j42oXhyuVoS3lpdjTk
B5jnihauS15wgUqMvasN3yDbn09ug4FdukiCU1aRtK1JyA1S63WQGmK9Jm+Ugdwa
7erB4V4Mw6dupO+2kqb+LOj0AjfdcKtioASQRDuf16J04vgu+CiYNF2OYgiW4lmI
S2QFU7OoH6iIvpyMjRUVW7sNTCoDN65/SIWlWCapl7dbPhDtTMqha0x97otLtIbR
cTiu11SGjhqHTflfBFZ77t3jNXfIxjhWHhIM60PBryAf38Oy0mJlzfg78Sk8iBWO
7maTnch8NKQGn0MQ+PR+f5qOdTOqw8PA/ok+n1jnwJKHJ94f3Tvqg6idyFA+kn7p
qy4rGpOXu7EsVtBX9DDoB/paAFnehIel9n7BEq1M//gjk4U1HE2MDjLx+DBPJNJo
tRcxZYR81WXKu4E2fUZxmHyTj22MoQwebRsLd8oMZXOeniLPgpc5IxGlqoWCRjkq
LvVjuYs8F1DeX0ujnJWJdY+6lf/4baavEOYmBwLMT2hJQT4a43UfkHy7xax3linK
gF6ax3kQ5yxypdKyKizKNeof4WE6qjueurXuTIMf+CKSujKh0RiMcMGZfn0BWwwb
ZKcRBb2CN/+AxzksNgOI03mndL/CreASmfn7jqyNlrdlJ5uFgkDsFCqPdV4Guw+f
4KzJE2ghbaF1HBGo9ZdjXnNB/exZyxevwzzlCnLNy0ERkeIQPdk/FPdK50SvGHcs
r4KrBhlAEICr52q+A5AwqPP3C8hv6vG48oxVsJT9PEY1o2k3l7TO17FFVKPx/yS1
vyET0V645iCgIZ+Qpo50ppFIZ8s/JbRNgGq42VzviOMNxzRkxEUX8PhIkkuJ6n6a
TDIHjuWKKvQJOpFc0bnUEnlveChtdwtLPW2lA0ykpwttaaG7uZIZVpereUnOmTNn
rL7X5FdoRUgCDk+oUQfCM6zVx+7KxFTENBn/IMseewDFrYSIeC2WBrU5KsQVxoSP
Xogo9Oc2YU7RBlV/p4PlnEZWVCbx2flAx0wv0g7fw6gkMOp+DKek36+WNUjYwt7P
0B7zdpQaqWSdeBKFOtbk/3vYAXGdZeOoUqQPd5WxisQJU6kdHzvvissyblKTwztI
/gpVM1CVyscb3V2TqSVdssTh1v3DETGGYrehLSHCPLZIU13TZnou70QcY5XWVy5s
L38Yo2dd59VGs/JtyXAJR4fXImTAVNwSJXMlkifkBnU3TtLS//kXT9hKJQc2g00g
XlCVBl5aXWynxpe24IyVPD9iXKrOdJRkQPrk1/eGlNFqsT/v+VoGIWYybp+8mUGU
5l1pRUACsT1DLBdRYZJS7rZdSPQSq7aZT4uijffwYsak0NH8OHofQOTMIr1U0gYm
vot1jT1+3JJg/0l03xGuQysvDmkm6rCzQXH08DLpaBndVadlRLtjR2U9lF3wKasI
0nsZ29egtpUIhiWvNp5DwSrs+w0Cy/Qzt9uKFxwyZmbxM5DfDZbInQUVgIixlk+Y
Rs+cQsfOtir2U3vfWspi1AP9PmFebOkaq3P+GUSSdi78SX7fBKLbNCjNt+IUI+dX
nFsUj6CFibB1CVpSn0LSN9IUs8UjiPtIx58kTCOK5MuHePc/2geB5N0TwmajNFSR
pR89yQyPgBZ5GzKBvCmagF6NTZxOuOZUApA6fP3MZJWdMT7iNBPXdx/1z/1nyWT3
b1HTJl57dxWeTlrqHRToxWJa9P0kq9w1BCk+iH3vFjOa83boLZrchMudxZfUMTxa
Ox9IeL3aQNfbBBDNCfdimUkOs/BZVzAlbsMVKo9AfJFnbSysysPk0kiZ9f9EQVVQ
RL/dzKZ5o310xdeQQNGTdcILygTy4XAV6zPC6XJjvfX7GT4+kbW4qGDmFSr/o0SC
gETuFu3xbLJmErV31kmnM+dau/ynuhaxQkAa7IuVSLuaVrSMWkILSa2KhS9rpqRK
53YNT7dH4ncFsikOEzGSqtTrYqD0NDLinD2Ukl2LIEsxvh9uWpKg6T0SF74L3az6
52nbSjm5rO5OJl722hf9sgXb3txYbgeuFjOLwsXFux/DG33LL9q89v/n6nE3e8q5
1HU+0/6sEkRvQXnP5OHeRfDNksV8Gi+L/9Acvp6ajoRMFi96Iu4LIEjMBRpp3qg4
S6DeLIGRVr97xaXie0H6UhP1i2NUqJLgHOQu56GFv5ZP6cZK8EUg98ldxFlrB0N+
RFZlqZcWDqWnNBCrCHKeX+9vJjMegOpWboIuRvrQOaVrIDcnaZCNJ4RYvmDuWHRJ
u8icrVuFrcu/ywp5HspdKIQMjrnSuQH5o7nrWjsLpLFd98rntDkqNR/ua3djG5Bo
pzXh9wKUwpIjDh0vyPEnhE9pnF9uhgjaVkEUN43R4V/DaK/qexZNfixjXwsQ5StU
mzNZWZqXAILcACquTPxEyLn9plv0tWlboqDyWnV1bghm/qFG7CTmJigkLEKRUpWP
SLixV8Cy2QPlmDZl6QSZYwBeKS/op6DzFX+zjoKNP9Shy1R+GyLFH7sM8P6TbOL5
0qYCITqqPk5IhqDOu6+uSGpG68NflnMM5tJBBo7XVQqCUUTgx/K8LlmyIIZs6CHd
emkP7vhA28usB6SEx9J9bLDA0oDDEg4SrHc9aBDD+QE2BrCGeIJGCuIfUSl9iQyt
kq9G/bwwNpYRbfYQSf5uv2xHr4KE7/BNvVN80l51kCyH2WZiMXosBBgwY0PINKsn
feUVyQImXmtpqvlWgvMbxEO//yXpzdFlJLnPH6HH1K6SMtEDFuEunIcuFHpPI5AQ
qZ1/uK4KCaPaFEIUY8/mTAdwohn9Ar2Kz8P2RTAsajII3E0iSkQiKOvyI4/hE0JR
IMUVCq3gVC6DRmHYZDf2NJvuOOVigo5XvlKhNaofY1mpC9gSHd7c6+0t8/Q3I2Lq
Za19ZzDtGTF84TIunnatcdIj/jbc+zCoZBXiQLHmI+vQugzkbFe13JlOdMnmoiZK
yazT1HLHTRw6aZ+wovZoH7mvgVAPL5dFL0LjSRcdQrXpjeKnIzzK1yDNBrvB0GsM
0W8gCpcPB/LfRarWeE1KYgJorWdLb/DhqYXVAfOOylRvfgogsk04g8Ohsbc9SEw+
3Qlayp7N3HiHRhjcxGbUhoYiJUaQJyEaNMavieb9IfysMccCLNunt5/1WjX2PG5H
2ixzpag2mc0J6yeBpJKN7q6ExygVWk6TIK6FnUeBVVIz+VchERW+oe93X4pHCzCW
GmrzX4KctoHCDO2EQ7WzsBlP+MDVOgDUDKiISOsfDdRJ5vjZKjTCZcs8k6ifj7Vc
GYVuj3JuOdBssdNGRxfgu5N294hwbNcRphselUK8x6ba7q+6lcN+uqDUurWu5IZA
TUQzZ1KqEauVEnvQpJs4xQOBc+QZPXIbD6S3PQ1Dkp6NTZ11PjSeXCQF9XjjeCsY
hgsqNmuXKb+hqhU0PaBOTOsa54dW1UYtrzPiy9/ceK3yh2P+JXCXAWGqVpQXxzeQ
U+Pc7znjQ3/Lq2F47c+kJui9XQK1uSLM2w63e4E0zFSYyj26mVRpqB+AHNjL8R2p
DZfrVvaVWWzWm5nXcdfzfOEtHNrj9JTPrfLxnJXkxRe+7jV8MDDJxXEL0dPH+4A4
qPwEYIEQnvaBGslLv4CzvdTMVXAtJaqUd1CfyBS7760fYzKMrvSZaWx0CQUDrw9C
v6k634cboQewOoy4rHOykZ9odHgI6/c5q9/jlxlXVxQBzO5WWM2FjKx2lcICuAhv
zyV5WBK8B5dxc549syhJHKqabaaeREJbfReveuYwAKJxztxh+OFf8Pf00LQIezVt
i/Onak7BM1k+Rjm5nrsi+qVa/AFyUFfjqqgIE7oL55nNXuTh5JFP/QZ+cFnfqYRZ
+bYYOKpGlRNAjFtD0WS5ouymSQ2sSTdD64d4eVAoCA4GvM08g4Og8yGD3gSPF/gf
Jm08c0eGh8f+t7z751l4xQbxbL1kDLSe5ZcRMYpZt9uLVozxHrY0RzZrYbRS8g7g
dSfH9EJVEJW5ryBKiSNqvpj7ryDbPSX2a+qNsb5ePzd1C9KlF0+z49L+T8xqhZdW
vTmQg2LKe+bgLz8PnpZ34c2EyX22G5DS2RDABMt8TIVhU9bV8IwNxvuJBlzeMNu2
W+2qitOzCLeeidTu8X7DQWdQ0YhJ77VqtmeB9nVV/6vwErgXXe+JWpkgyCx0UqPZ
UZL5l5g7TTfloZJg44pB7RcBIytktBE7Ct0mhhX/tyKQtS5U7kjALg2us4hvNi1y
Zn4ewp0/2dpxWhvQ2zXFnYas0tpB3IBUJZwh7hTnFxLaNwHnVLJXBmLck6KtldLb
5BqWowCTfHNr0mZBBCUwCxvCde3/FA6KjFlQdIqkYrGEmjlog9Ro2TDC6sM4oS3J
SxtDWJ0tTR3sZScHS0KkLh2ueHE2apCyTA+4QGloDOaJZjHQ/8Hho/4krOgJS7HJ
L4jfZrphI6L1HdxYpbCNGRv4ZK6OPFTUWgNuNvdMY2/gwpOz/BjJfyPSwM243Ehw
5Ro31oyt80IAm9pAz3qWq5R5c3KyOPF7OU938qkEXF3rVU7XZncAWnPNO7gg/JPh
kpWvBZbvXAOVCuXxVQ1lxmhFeA2ikOBwHgY7996wJBFKUCn3UZ6T7RhClJJNOSF/
qh1QA4jFuE7/arYZqoR+CcQVkVMA4YP3U+IAB9Vh/WNrnxKICAudakcS4oi8Go1O
SPPZKxeDEles7Sn0hq/EFAGoO5dEQdknVWFBD9NgeF9LDwvlmOsUBy9xQGhlxhQA
bxlrtd4KYP+9yEd0DCT/A7R1tKXD2k7zvr2/JuE6p6sQQlC3FLdHHr8NfHYzJkyC
nrVPv1yfc0//0AUdqY1YLmVpwT85Dbujf+iOwtLBfSNd5k0V3fpeh9L0JvHvPD9E
rzRPh3gg7Rr++Qp2YJMeXII7KYdutaWTzPB8AlWux6p+SoDamPJUXUxhpQnHZsY0
tk7+gjN82tfvAjWYK5KPOvMxzl28CrSsUu2bpJJeTgCYkngpap4nxYWxO01GxK1F
NveACKe8bnLGV3fr5C91pLdlf2tOlBJNHsBupCcip8xPdADrLhYeSb1e7qOI8hft
o8AL1ECEry8Duuk7Knycl7MNWUvhDsrN1Ak1ubOAzkbW34GrOHxMUBfs8SeNmOmB
aYJcmsiOgna8WG8vC5pkQapFrd04Ip7BniH/TeixqDFugrbr4zb2C1lmi/pPlQ4Z
5pxlAdEXPhFnm5gF2xi8H/r65gIcTnQkdcjHXpVDE86FjhMlrsu7CfITk2SBPmru
chwuyvNp5YX4HFoJpA92pgdLgoyzPyzjdabqxKVj+2m8Vz4GO8v5LJK5XFs1pDdT
1gwxqgR1DsuMYHK1OPoi5vjmUYo6E0Tz/dwbF+Zx+k8DiLQDFqlRgitD1feZrRDA
hSo8l9RJgC8+WwTWT4no/XKA4gyQEYXVjxotZGupbPMrr7kO0B1Q3doISqmBQG7/
5LU7DLUhEuudB0HjQgQyeRKsTFSno2smctM0KWbYH4PiYyDs0TO6dnFql6dZBFGa
DU2y9szkViuP9nqI8X7UQqyl+F0OEv+K/dYY3ZmWgxNUkvMgV0pPNomjFeLlbBTI
CqIYuHfiOsPD7vKaHmPltmvc3iW3GFQefb4r5SO2bWvtHlmnz8VbR8dHcx0gVBN1
fN4DUte5kjX5lmXXJiwqvzfjBMhcHdJDuaYqiz7em+VGBbRdMoL5tnRSqOFIt2r6
zWoqosq8+xKj2n9t+KgwPPzW2Xx7ipQsIGq+xdbC2tGUSKc2o4Wbc02gCmJ7IxG5
beDgwayO4SY0l+3qNIsCIOuJshsuTw/AvTgpYfu1aj5QzP9HyzhP/VZCZIOI51D3
+Y0h6UWwQbB6o/Uh2hFsDgLuiX/lvGooXY8d2KngNm+b084Vly6CRrrcLuHmJJrB
HsKR97f9TxFs4p93NoPmrCoxSJ+leUdiVePhbzUDYTeYFHJZA8ocdZqBg3O60mJX
NWhgw048PcBVkLAi2fnSsoSa9W/Wl9T7PJYIIVvTtg6HlC/MiacKsSpTpSK4DqN1
6FOm9bSJWGamqOnPpRQIWggWmm5zhTlSWNiRkjoUou+IFklvkP7nvIbKrZMsijKI
cbZXvYnj7Oj9OokAbfhY6jRKR7MfdshybFBynfBm76OvaZHn9DLQsu5Pj/GBW9eC
lecw4TadI0KsmKk4LYPTk4zkk2ku43xUcTF6gUQMYIS4vXhvTBHDWCYq+Ru8DM/W
ua6KtCA2xZVTp9e9Kb/rems+mQMcx3bkVbtlB5Q4cTKBbUOlwEuGBWFRJc2gsfyv
n/ni0um4qthuHoZl7yK/DdeK//XYRbvsg/KEKs9ne6wuVNCm/y0jj/Za8FgjjRoz
SqAibvDQRO+7U4AvKuEaLwK2v7YPPaXk4OjMdmo0iw9SAUA6IT+jrAAm870JMvr0
AiNv3k6OMcf5PnvryAgG0zfzVG/GTrAQMUNJNq2hxqV/qQIEEEHlnr74rE06R1zu
0bjz0hLJvivyfXKi21WdWgLpPzDd+Lp7NispUArf7c3WBbJMWLoexKSuRXGaJGDR
pKckPNPMr/JT4PNPMtk57LX7eK/SLpQZhxdRxsapuzWLr9Fx/4Nd1wNn7gRgtczZ
HMWePm3yQkzvfAxvNKazkKw86/MoOi5IBJIxtYSGpReF93ENUpVzfR6V5wl0xCZp
DxjdKBvOMdrRJ7CGp+Ai6I3NBfaYYZaZU3KtJbdHeLHqu6GZOJYdSJryNwIbizj+
Q8ASPf/Jmz9H0jnaIeRYfCe4c59mczrNPUzkbaYWM+KnAKw4MNbI6dlEeyTFNRCE
kfefBKONUA1nbzjDew2LSb+EMaVsdcvc3TgtMnWFwZ9b/5oxH0B6C0BsTTsJA2o9
AUtU8DJoziN4EruMROxmVz66NNaDAxN97oCEoH/Xt51fU7upyUziSZrCig2f1k7B
qag9f7ZFJeoMT+U7rEydt3WF4zijQwOXKkwqGmrmRnxDAxQKOF44XuZMYeR3pWBq
sP+XJra+7kIxnowYRQ5toOuaYCjZDSvDTl2v+JbZ7VE2/WTDVCkrjo9yw1NS72CE
sIaCPtfu4IU2WSuog7BjqimspfQMOVnCvo3PUKux+6sLlKk4ionDOD57yj1X7KnI
lp95hN9dZI7tWIOmmQpa4VjSYUSjObgmwIeEN6vj2Q7z9kAU9S9cCN4xu+Rp/m7v
RiVS7zsJGrScyPGSshCE/CfYpjiVye38VfvObJwK7FbkkeT67LFbqkTq1XkC7Ns0
D9W2BgoTfdWr18IMGuz+/SLbyxIteo+Yivr4Wp16On0Nck11pmosTrBO2UTBkCGZ
d5GmxqRWbGogT7ZKrdrwiJlWbshyayrUwNqrxVr005lrODs3QkVY88Ma4rYSFk4x
Iw3lEh3HZbDs7Ejh6G13ANNT/2Eyzn/xfdkfNBTrjYc9DJJ9IgaBZ0CXfvzzArBT
qItj4ss0RNYsRJ/zEnP9IwIfLAKlXmRxigmXJK+XvD7Sq6B0PYK0wgMYv2IXsukd
Q93MfMrNG/kmO+cjsxvuL4CTUU/v5M45BJp0hMZw9rMFbRPQnl8BIx0FMmD8SFDI
OJXzNWTwMMN0kYiwTtMBt5JkCMUVU5zGHzaX/nT6+xtiQ0vkjQVVq1oDQitiySNS
DmDD1alXFfCh1iADrhD3CFzaUR9cZYy0tNjIWgv6wExg6Q+rqNgrgegWF7mL3jqS
pC44JJkz4Wul0/4VgQR02nRtm4JmP0rBbebeFgqaFbF40pjERsCn3gR3WmbPCiQn
iIMw2O7aiiE5Po8Mo8pGbxODt0xYUtnNd3kyd9QlX/rXG8q+UVwaVr8FWthF5YLh
ENJYXTA3FjXAGSp5iPdmfLumTr/HT8CXMCHW/1QfAfcvhrYD9Dw7VE6yxTUMxrJ5
uyQ3bjttRXjSPiJNmDXu9rb6eFKXttGrh71PdKfKqMkPSJP8ZTGFGjeqGaRETPe0
sDTkeVD64wPAAnJsodK3kj499U39vMhsEkspVakclZ3Ler2JQjCI0Fb+9PIG05NU
se3SLmCq/CcXHkQckiH4iQg7rlfKZk4NKz5QSANnbwB0Qr2k6zbXzpDI9vK5EDHy
6jCty1EgezdW8vDLJ22+2f1l1kAWHkzdnPmE3df+58EHSogdycDuf6tyJCpKb/Vs
s6TyraRLNqgJbIDaJiYUipxzZPZiK4gQmC2o/muoDsbPJ7XvdU+LJvMeCTCOLY8V
6zTcmLXLVV6sXKz6g3xAHjJ+Dl94OEYrc+iQY3UkgMWP1zm4fGGDntFA1t+U7d0T
O8Uj/bcyOxbA8afVnnw7ZlU8bBBYLFXT3ffDF2FfgLnZGSC9SH/4q/lDL6XWIoer
srxjCMHYtevrwsBpaoSsM2LkCYXOXhtXNtJLE/k2Ta41wWEmO3zIT9AvRUz8rDy2
GSv0shWUm9YrhgbnEOYA6LGgKethbw3IFTmG8b8qsO2aXg68zYpk86gMHqUUHyQ2
Qz8CCOr4MYXX43JbWsCgEPbHzzcvFeaHcFsZi8KFpiiSJP6Jy6HMgVHo/unl+b60
LgleXe2rOqMYbCwcOhSdoZceyea3G18MlxBE8K+bp3yztUP9YtKtbAs34ITCMqQn
gn+XBPZImeUs5if72YKhSRxrBRMeCgu34RXnhml4M8s2s/MzKO5yfkHDNy2m74ky
fjTRRBx5IlzDl9wteokeCZegLCG6aCVOTseitLLKoVAaUr4gPk0qrAVWIwa0VGUJ
u7it07uT81KjhILwrtz9RGU9Rnmft41rcRw6emTAMxJLu7jhdJz8hb3OYWdP1DLJ
D4oWsysqfTyOEHDOZM3DgZ9YOB8P3cpSqoIrT8dBydkYfVGcrd+aBHL65QrYfpsA
ONPuUQdvEcpHfewAT/nG0sT893qKgTPZnvHTfWPaOAFflg6K5oEgZjL41cwabGTL
UkN8V5T+m5K7boW0J+MA+eZUmBztJN6/pGGiuL6N7Eft1UGzbp73E4z+CJk0pRev
h4yKrV8aD7vMJ3S8/3YC5sTmDHEcDLJpTl+GUol2UpiqYy22mtrwfEgpf03NfQ+U
Cxz94hyEsjyQanaDDkggtXYCZmrzn77Vr661PVBxkYFh/kmfq9zz6iwQejySjfTn
xMdlUE1FoXlVtDhfzq4KPI78YLYUPwsRKo9/P4nLO7fxNXGb15s0Pwqq7BNMDSz4
xx8S+N7UgD/1yDqqvkKmwg==
`protect END_PROTECTED
