`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5m1ImEuhLrtjbRmhTPOI26bU+QKZAVS3V/E5uLH+mAwqeXAU9/NRcRqJoiI3ODB
KFq1f/19Ju2f6RersvRexuk4KplJ0lDqYOLQbiNyNxAICYc3SvBJccl1trZq0hWo
mVWOCSm/+t+tKOAXQ4jF7RhCjc0pONk8/WgKM5/txFrCNCoyeqd+Xr8UQcrjJLor
2XPUHKlbtJlhD6J/41k0cmuFA28BFXTtDRQ5lRguJws18WGz22LxRS/SFvf6DxGN
gg0WbRKNgvLVrbVMjIWXENczaVyL1Hfy8sipEOby8mLH+3u7MCTSThQGE099UB4b
o3S150O40d92HDHzJTYj+oDSTUkvkqy6MA+LxBB15nSwR7szBVnKMvPPSjQbLaqx
CiBFyJ+8Xm2GccyH4nkxQ0zdVzthbwZTv50G6yFG6xyHCxcMk4jHp8lfapSWluFB
WlqGcXnokX6u+qKuKfM9rjywIgSwQaXwubclSzx4LZ7HPdfCzAwlq9EFnQC4JcTS
mNvdsCx6HQEe/2Juqr0OyCqxyiVJnHRerzp0HoOMAe8L2Yjdez1SbK7aJ5u7+1jJ
m12k7ezM5qM9zVcxwxTuvrnqIDFxtDez7mUu0lIRVzL7oCBXgeXm8CU9EHs2BHXl
mpvYZP6iUQYNxr1XzNYnk4zxHvuBoywiG398smvRW9eW8B/aNKybuHDRQE5VoVZt
hVK+8grg4Rtqda1yIPJsPK63xzcuvB2Ue+9Ue/tn4psm/u1G/QDGVspg0/uKL73u
x9keFiA72bFQ0NJTHzrM9uzTck1V/+BUnlufFmyp6lmW/iwNwd6GSJ7tCrZuKB9o
Hxb13+Rt+sqMVr4vH0UL8EeQTQWrhZT4wszt53RNiyG9Qo/vDGHK3zJzBSLgrzjS
OwJ34pmen4z0Lz+rQBfqtp6oMtG5kAzwnDHQWA0HChzCv6eX1bm03ziNhQSrUEZM
YBCNKQ5msYxhwYOtGPCDi5H6FW4gFfc40lULnKNrr3v+RqWcpSWV9K+P06RzSJij
f7GuYs2d3qeKKEg01m80Qd1CFZWvrtly5jojRR77j5tPQDTkmmTD+RWgt2m1a+ER
q+oWerM5ByHpl9Mr1ygHmBmpFIoPd1I1J9umCocVJD7RiqQOahBq1WanIpBZgeXO
wz6U+vKV/bga1TKv6O+tkHOTDISsLSzZbAPHBnYZYzX66keRPb55sBAQ87x9Zy9j
2ODglesxLeI+sI8bub3AjXmO1E2tQ8sXMc74SXkM8yOG9vb5mNpy7epuV+Pde3Ke
7gDCfthEmkxdIAPGNYVDsThxm1SrU97eu1LTtMDO8hvbv8c2tLwbRNE+NjWwhvd/
SucErgY1yoayefPQb4/bZ/6hH1ACxs1OZy9dh6on0PjRyliFAOEO9vv8wk4UNyK0
MugzzvrgyVWTIa9fcyCogCKTJKz1eE3T0ijGdiwr+cJylUvQKSb7ClvLlaAycoqg
K23371sveBv62y30YQ4D3d7OW37ubNifrKkbgiFUYQRhZ8EhbQopylxWDDAluKTW
fmapgLx1Q3w2NJ6KltdtbtLigtHK8uUyrSGYsNWhycvjFc+D9FL9wHKo/otgJR2P
8VvyPqCzXhmh4LK2L73Sr2soPjcKgJbUiEgLxpPdVytBJrSFfMmvVo8TAEwbsZu/
dzXg+Ye3ri8rUIdQ122sLD6c+eHqqn2lyzFhScVdziOaFmKYZd5oM3Yu6biTh5S9
P6/YrNZeS8rw9KZgUnCZjuqnLjX6LnENlmGtPUyRDCb5FT4iW+qLm6hpfEJoF09L
yh9Bz7mxkLcKXzBhG3WhV/CCIo7AQalN6NNJtKX8zRoAsw6aSTfmAkX52EERxH//
Dh8zO+XJLBosOKkBf6QqtwE7eU7t4LkIuv7D/BCS5R019vyRrnqrIY2P3Ds8JwMj
yBfhmNMBS97nDs+yRfO+8rOLrLDDokHE6OMJ9ktH+OqsbXb3IgM0Dj6t9pUv2tHA
l8KM/6/3gsv2S0AqVwdIR/1MA4HkSqWTpIdrJc6ldV/FCF5M3jdiAZECYjQVNHqP
fam6xUE/0C31nM+osQURGz/m474Xh90dZLZnSdaP9A4huxNUYqD6hKt0tmOGBXqE
ysV5QOcRIh38qYsSwLmyqbyorVWwqZN/VL4qKrhUo9c6aVGNzYhaNB8/HVRSWyyU
LKYlDRH8noN7Cahq3dMT1fpiRr/MCWXmOg+bJ81175uNhiYo1zowKp5GNsRrQja8
lglQlZJX+6EafJPO/PhTPkCGcEFq3e0rFw7Bw+arXmJVOtod/Os731gN3fF/0egg
+ddjo83qNQXi6esvKExGxcQbehT6NnRketIPBeKcHIBd5nFnlp0BzmKTmQs3rSZL
jHcXUVnS5eF5cfKHK2uiMCfWRljV1+/SyKxV6TDemXaYZDt0GAX8B3RDBVAqsVyh
XelSDhwReyMldu6tOIwbw6TZi8d3lnGNoYIJyeN0bQ262bn6jVsL7qOVwjq6RqjN
Q7jjU4DSv0e0/vAnvRN1qJbrA66hNvTghvLbG+ma6+kXwZmbMxrwZdow5Znlp5YO
DgRXOG47U6EEGQ2IKt5lUbd0XH79EjIKzr502qVZ9CjqLrT+GA5JAJCtpoDVP7yL
4GKFwG0A33SA2dMCuMUNCHi7yU1VFUkXjweW/Rr8PQ9ZqANkSfMBIzQe9NeYoWwc
8SI6CK3Vv/DHyLzKl4GXO0Ix6O3WGEczBAic3e9M2vkAP22YKms2N7uhQMGPV59X
xCT++UlPXtcqCRPyWs9U/swnBI8Bz3lGSMR3OuDXrQtvF3CpiO9hd57jjaMuWhh9
lpliM8Qu5WiHgzYdv0fJThUZmB/3vWIQ/Pa6m0JUecyv7fin3fNhcBawuYqEcTMM
scVNHb8HI9R4FcyF1quowNUPyvo0stOGQQG8weD9i/LDKvI1SQvIjkRZ6Jn8LXKB
ixm6JVY+tSEGDlMdgcLa827tuUfPyWtD1bDHIEGgSjkq3yULbHKoqPXF4TQFBDVV
Gja+AMA2MJkElMw7d3FhYCVus9NmOi9dArPj0YNywJqIy9ntesbjnWZo2dY+/S85
0U8CR6N4xYL8opE7s7GHK7QQuYIqkG+J0lcRvTJh40iqxX5nObQuEJGETxxBPjZb
3FsnHrFurCjEVBl0rQwn1WLJfitXFEUUkcPyaNGHSFiqNccAbFs34xLIZb7fb3Zc
AoBWmBgkjQKgXWe+M0cpx/8Cz5mKZ3Mdk+0E6dfUTFSdyvK6tJ+pXNNBrbK6NC3o
N0tdlGx5o433SV+dnGxJfZU1S8AaMhCwU9yYwiYbsQRDLrxUww8TFL5ZgyeRSF3P
utLp3IC9HW9c+1dh1nzNjjEIgMW+16e1wUq4W2FVHP+kqtbP/2tPoZMJZlQ/Npi+
JQbZQsy70eMiaddCTbPl1lAguJuGuafVPG1620enhZS1wTlt8MrpHe9zq31SBepk
0LLNUt6tQwa9ntCZHp0Jv1nQLY72v21Fce6uafZHN1Q4L/DRGusedIrKTBELRNf2
baVONSXNbkcgodtAXH3Opwxc3IWOSDcwypIRhJ8h93OjVGWORpIErbA+A214cmGB
tiU7e7IsH/BWN41ZU2ekByK1E+wgxJDGc2WDLnVE5fThBl5M7tBYcfC895G435bB
WOlOm69FppA84rlppQgx5AApBgXT1yFKh2a8bN/lV3YBhGQRLMxGwgp+h8hPAOjR
F2NrWE7/lWaCCeokMZG5Q78o7DuM5QwuCRr42Gn4nKnGwG32aeAUB6FezHOo/IUw
IqWxByyqISb6LC6sJdAhZHqYjQowyXSdXcGFgQ03DVm16EZ4i3w8sPW8NG3+IhBz
oRPk/MSvHnS1KBu1+4asjl0l30cdzgeBowH9pnW2UAvWX7GjQHYHkxF0749BjPyl
S4+/NwWD49vsT5X8jBMaVXYiUJi4fJr2AcgoPDBcT1yA+999sAG+bcv5CVYnh53/
KWvl1jNsWaj7rmLX+LVujKoVw6s2nMfSF6OR9Xs2EUuELOZjDZHhVssjzu8UxZPL
uZ3m/dmnIUbZ5OgLRlguXCUAjB4N9All4bW0qKHT4rik5KiNLE2rp7YoQPd0lpYM
+1kHOALZGaj5B8JCZkrjj8juHU3nGa8j4jngRBg05ykuQpj25VGX27HTlGHvAYHf
jAE2OTqRYgsoKbyL9smosNMLOhK+dmNuGOsxxoij20Wx1Dffp6TaXhKyj0lSAsNf
ArjKUQVG8YbyH9sD0EYCja58Pa2efPA3+6BHuL8er1Ey47zeqTnpOIeOw3LS8hFn
vAN5ytFXpIJROWDk/dyFyznne2M9yBd0UMqty1CQQUryvNuYFCDYw3CQ6/8IRt5h
tSSs5NRPq0QFaQwJIjaORTqNIFwlwWdDGIsx+aGi7pTIxl2kahs0FolXlnL363IZ
pOZOzNs0FMHdLEflNkDTtrN26kIcpkVhM9W04gs5yQHqVIxIiwx4XBGsO39dgU6G
f6mL+U+BW0UE4vGwT9WY+fPp3MNcBBLpot34FmPn5UGVxNA4uBoevKLNn188u4ik
3vEK768eaXYtIXpPUwkgf3dhm8fgu+QSMZN5cdHXARpeASPjD9/JDrdB6sW1dYG4
tLRNVsgYJPAfWHeGm53bS733tIgTp1g3Uj+RQtcRSlUO/VZqq+D79K/0OBzoWCTz
GOFM0mBqh/zpOA1o8GqSXzaiFGIFVKdIY78ZDQSbJDGtXr6z91wRQzTf0w10ZCQb
/UsmILLPOK3EERDR7gF+uh7v0OWKKRz0ns4pqDuuImCk9542bCfWDvJSzqU8nyVt
ZOwJjX5EmyHUDp50GpPWXx1689oXpjUVxrBkvh3+CCNekS+mbnKKnBBR4mLwCT25
CMplMEFsVFP+c7VZuNbyMCO3DtVIYhacS82fBudHuiccpQJec2QYVpnSRaI9r6ZH
GP1zjAFLWXFeKwCZltmHWpnzS9uNdY5mPfQ5MueEBw22FNm7xIrkdD7NhG1Qq0k4
j9E8KShsVdrP6NB9P+z5OV2m2Hh622Dsn89LIsJpGq1YtRpCKFn8uA/515yKfmCs
PBmuSjOWEh0/hYxVbmMqstu7azdX6Mq5inhMasHpkKF8bxSicHo6kVs4dbb39DY5
GkHDdAg71/0vRq69GgKP2ilaGrdInhql+O+NxMk9I4r6dajOuuA+LhLjTWiOdk5h
YQ6aGxP/c2jkRLw+czVCdcoXi3nR5c4BsRq3DWBooe0S3+80H25Qb1DtBR5EAwc4
/b08Ya04ENnE5l/R0oNHQYmtcfaEJscDEvCiIo/WJe8uKvlZOLUO8cJE8PWZx41p
Jl6IKVddZRUU6+fMKDSYI1QNyc0BeZHz9JiiVssrdgzDmjwAiFpu7IgfGwydhNki
RnOewqw9g+M1P3xgnVf+TI+7rA9s5OSsvYd+kl8kJRBRd48kzqvW/8UstOij++8n
cCd0SlDH+rK1J9yYsc3bAvNJL2/B3HIdDxGlt0l5+CpGleZIuXQFhPeyt1YhQ2Z4
JxURjKQfZ/yjPFS1A9WkF3+XKw/NtiILv9UIjt2gm0vz+RD7Al3Tq7dWCgazkEwA
5mUwPHSUDZZpA9JuAjIus/eHEEvqVy+TDeQ3VEgfwvOoVUZNKtZCzDeUlquXtEQq
KHOtH+4yJW6V+cyjus7gugGSCRm2jOi5S9c8OOpQQgY1rR5uD2vDgURTPhfAIY+q
OZ3UR7iRLjS9+jeSNDwPwa9nzOXTtQ3CnEV0mY9CgufRwQdWtGbC+YzZ7b0Kacnj
Clo6O90UmPu2auRkPUehlu3E6rfAA+7joP0U2WV39rAQ7HIADDhInBnG7Ezvj6zb
POC8SGXXU6yE+IyxJUs0BXc9celW1L35pXOPEzGJkqyosoeGBpPlwDL3JBRJnJ7P
S5nMFFqcNXDbwMvSi5AhnueyC34DMYyKn2CfG8/k7V4Bz1rILA1UNCzZDNm27aaN
3wviwdQaHcUMyesfA19a8aOAU4C/+WpEgXqrFQnpBFwvy9Voc9ahJnh1yHyDc95b
nIDojTurXaewItvJjHOttXI/bSTVl167SfIbhRKo6AJ7QhaDiVAV7TbyeKf99ZB0
tXx9vC+btaWJirP5BviIFttiF+lF8FSy1//0Wv3n+CvVfJfsa4LEiAlp3SeWVrUt
7gsR+5Hsmgxrrjy+fKff3Xzuf3vNk89msTQ0g2DrujHhjgKy8CBlY2XzuWIZe53X
unVBQ7njX23cVZTrtVQvE2tAhzlmTGZz6koUqi8STyRfz1Zcd1byokUT/sT9rgcV
YzEPP8sebYqQFS6mnNtclLXSMSFcbpRjtT8XKJ6RcOGEfcRkc3tRybwdPy6iZGMD
0B/LJ3Ba3X7/gnTb+Z94QFqECZNMZhRrhAVEE+vdk+KjWOepqAmy4o7XSL4psm8B
p50KEIdfGfebxV55lLCWzbZ2rOaGhOoP3XCBTmdG7HeoHL+SdCi8l7aVy0fpYEKO
GzUrLM7fmwJD5JZ0cVW0hfsUpjTB2zquMt0CCUbRKvdkElAWPn61irpyoTnIfo3+
bl5L7oIedtOJJdF2Vpgs3XWF3S8fbniFOk2x6jriwH/4Kd1KEziTQllQVtG8HjC8
qYd+aDSuzeHzBer8DGFHmNGxt34mhP7xmIXoY+P2XLYzroJyzBW6g13aoPAHQsaQ
uMg/Uz8gi/vl4TSYxZev1xj5gWpXO8uMNDthLsEG5Nhll58zwncn0WfuHMsEVNML
Pzye68zUyOzTNhsveyQ024xyf9a75snK+ryDnYWdSoAW/UJnCdO2Ad96Idb+szG4
ctmlcVR+6tKg8oJYtCXPh2IAZ0p1J82o10luarve1hSvVLdFdMENT9D1Bbf0vjZg
8PBysAf5fw4Ul4Zs07OjQ1yqaocL3cqBf2g1UAsUJC8M00tZuDM1f+y5cQeoPjJx
IvW7nYqKyi4Q+nS8MNx9Ll4w3tsb+3g8WrwUCtJIuYfYXv/xcrcLwFXir+pP7Fv7
XMOkilMTSbQ8+g7zGa/ef43EcElLVEfB5lGr719QoT+K6ODw1FasZ2zFrlMQxTXS
4NUZiH6iiO4Dw5CannNojMcYq6VYU5CCvWgU40SltbuvhroLivCVIyAXLncDikrr
jz/hSHNRUzGIzeuje2QhVA2ErbngCuWFigAdUtu0mjRnIIENhNfawtjUzZt8t19a
9SUg6M/MpYN4Bvd0WDRljTkSi1ba73y2kKyvEgJDyz4kKU3lyIPmkAUlFHgfPExe
DBttlU22FgAeZwgCMgvob5XBj5uiJkT6p3abruM6qdE4e38CEoHCzkD8kMJOoE1U
zqptCY4HvdxJQB+EeiJ9J6DIwSP5DHMinXrf82hFVuZ6ZU0rqjCb5KoUD9WCtxHA
62U6gQKWSJotWaAwFgCRehh9UnGF8OXAifEuNJe2hNZ4QP/7PyaAGNiRAcXQzSX3
bHxzN43/26HAzSvNy4yc71Hc7ZtAwLWtzXetth/1TWLs8WCGcNTza7Pexr1iNa8x
2NTeVjH6cTyjev+NmjxV2Ai7hSGjoV5g8RO4gR7XMgXFrQUMKPudl9khfvKcPUAc
qv40J+ZO+itsy3A7X5IVDzOgeUjwPZt41D7en+4GQhGNPMwfseFrHFdYw59scos1
3rAF51/Qnc55FX49i8ACl4xKWYAJU367HEyHgBM+Q8bHeuSA5ktsxWp169Q/gcyG
1Fa59ZgZcK8WnX+kAXnI3hpjA2p7p3jNch0oVnujzILqzbiyjFiGOloK4K6DQ08e
Hnty7sWqnsX9mVcXwUG75cWQUCsecsUktAR2Hwy8sBl2RKlRmcO3r6x8WpXx6Jr5
sV+waStxLeyq/VGlJcski65CEu7PeTFSkom0HWV7yzQENhsy4qjJceYhI/gK3uEY
k/kaskWqHESXSPGJsP5jJ9xcdBszLjJedpGL5b9BHnJL9GFEM0K6V1fETJKN7l4D
Bsku+qPgtS2JxjKr1LbdF9kYIaKQFdc7eiGRxwEsPVY4PcraL8Pt/c9oo97Iib6Y
NIEgt6tTo9iaBBrtXo1T8ISVRaj2wfFGc/WRb8YeK1CpQzPNlalRVID6HvhITW2v
vvRtNqwXWP5CDyD/tkMvmYnIe7Sc1ZuW8ESbOLCMjJ3ufrYxHvmKRaZGaJZl2HAH
nfRLBcRftSApOtDC9uKd+5Lrz/RH7yMq6jsseA0g9i/JxvvCetV3jdX+tKbDPYZ8
i3N5Ifk9bNQR9g32V/zBeb6v1Dwadg7DRBk9me5beuu72l4yHltwWGS5JOPHbYYt
U+kFB1yPB3bSaTngJRGvWqNtD/iUXS8WQpWAVosdolBiAI+mWznu0NyeXnrkHMJp
byoebvsJb/3rQ4jVBvCzR6yZ3yR/+v2wSvSLxvDP5YU2Hn0hmcNbZv798qJj/H02
mzEHjqQx1yNiqA7/KliEm5ggO76MmxC9phnPbdXYP/MUx6pyXlVgGSNF0PVFiv9q
qGnIMuRCBeoXLM/OawsHa+kd4sNh9ohhXo9OhNxVba11MrcW7ne84KFwyZ1qpjZJ
eDvlZsn2FWstoq1Em4Nhx/NjN+Ji+uA712HxzJop7iz2W2CWA4vpWbwDM9dFFhXo
scCb4jJWvLGIpZq4kjMsScdaM+K5gHP9ZwjBqvD2BE0Rj3ghRTFInUPNyVO61y69
SETt42l9QXserk/f3867/pcADgp5gf1tm68joIcwc7lg9AkMxt45cZq8I6PPI/iS
ojH5n7y3R4fQ9UfghlOjO0hyq3xQRPws61vicK1mDPDbJhOP/EDeu2DNnM7nuONI
gCU+hcSpVr/cueQwQCvdQEL5JnNs/vrstewvBmE74mB+1n89MXNFd8ExnSEIcK8v
CBS1Wf5Yb02uax9rikkGZCZwJ5vGNz5tD+oorjn9XB7z/vwt/MqQguDttiPDKOjr
c54iBk3/toVXpK5DFL6g7wzpUCsV1pN6OSGrUhCSJW6YHeqjb5utz+iblTsiHSi4
YqtalLN9Q4ZRqDZjol7cPHgsWSzDuZP9TpLqIE/Xhv6SI2tDHa+AVuNGUbw7a3tK
icXYVVGMctXr422pmYzAztspIrhtZsVMcX3fFuNkYYjvfkjquwaKSX9RrNeilEjp
nRjFYzarHDOshhm2qFhLIv4sXuIi5IqZSiIrrdtgnrMYU/1At9SfRZgju8jmIA+S
W1SLpka7KvuRvk69v+BQGFDY2hlOxahhTg3uQafong63nvw8Bi7/I/B9Fs8MCV//
pGOrJSwIRCED0csqLhE9Kho6ByP3bChZrKZ1GFpUhSceLWEmq5s6QIAzbC8J77ZB
/ZTn1sWfqy6osz7mSV0JMKVtq0Y6wJAvKv+X0YRIZmmjJ70YIdOF0WFcihdSyLxP
cTsGNPCLbZ8UJcA+2ch3Fzlf+cqMLqgK2QCEdZQx3kBS6+k6tRvSEeYDI9h+JoWd
PJNVzd5VqIHn0PCC0j8txSi1bpalZ08TiT1Y83xzEc1iPr6d7ZCgQGgK3RdEhiYY
sp6jQXsnw6otrj3CI/QEEgdk1GPqpS4EKTynfCOc28p6vfW5K+FUHRhtTAJEbacO
+WVmAeMbEphNWJoTuAZpGZBKdjtihga2m6GqY3b/nj0aNkUqDAaykCKbbp8gP5Si
yvoH8mRLWlHEzMDDhkfvK03rCr2F3fg44HkmEB5jorAU7488ZRvsDTVQJDyQWt1v
T8XstCCb0FyWN4Ol03BWAEqJk4EzX6+MgTM0ZQgGlF047w+SJO4YEqBDJOe3E0Pu
txLxfFQCHD/wM+HyqKEUtm6+YoMItLuvnB13uq1yH3iMK+FGTsLjAYX12bmAtYWd
htW7jH4XpBvTkK3qBo8yMwCSY+Wr+1+wOJNMo9Fqib9kL2kQPzAAMZoTrouBkBW2
CZlI1A3hQM8dB02ZcRVZMWcILZTYWvvzHo+RoRMsWkPYhe/I58sbrdqAxtiviurI
FXLaceROb6i4MohZmo60FiZFV6Vqhm92apo3FZVi+hjPIQjsoh4qsMm0xVldQzwW
YKiMVjKORJQdrIsPaKKYPP7xoJxeuQwqgQbH09ZYI7EjY0GPXTSijlVMQpH4yS6X
RI3U/cOH0RzNA+ln1OfM28ahrgt8gzERxwPNfLOnJtqKhn6W6aTOLWHoeUNYHkw6
dJIWgyMszt0wcXQ4FGmyOBWBgOy/yEJphoZcQEWiFCRBk+C6bz8FsffLiSzc1/fM
1oIkX1eJ7Pi9oMTcruZBbmuvCTJHi3z/FwNmvq92F7XztwfRoSjPpQhftTimcItM
mEhq5gz7MXne7VspIV4VWfvBzvxvrWdzgZlMZwaGLaKSyQXo8H3AhyqiU1J8iia0
Mxi2ZxsFr1LbIpjCYQunBJrRC1PvWIpn4Y/PLbLCY6FVSfvTNOk7z90Ah04B6ZtQ
pRHI/pBIiDcOOkKzs4wHlgWu3y5z+C7l8is+sws8mFdnDextsAiWCxO0tog90niW
8/359paZFqMQnks8qOe/JJmcAkY73OF4VgDqeR5pJoyz0h0sReNvos+WK6NuKIg6
3P7c10F5dYrhpyRuny9ntP6QvQA9k7TsEqPzYSafZ4wBTTL4MODPjaqumlrM8ueZ
Ss/KCULhgmsn+dRYUxPGYxyDy2NnBV3G5QV1gSRzm4p3IAf1RwqJN8H4FPmh9N0l
HX/ug3RHpkeKLQFCctKYXv9R7c/T4dumhY0o5k8s3YwK914Rdf5e11iI0dOJ/7Vl
1wLaZm3pGmSYb3ytYhuDuxvDm4MeuBZk4N5IOzF1eV5r/U00pgtp56dB15fljs7K
ZGn3nqC72r/eT/OipUcPVdov83q4niKGy7eh2MZOx7qlSKpuFTjQi/bt/E2vfWRx
tFqEVuo8LmylxooeRggLhb68vuKTy1XEH0cizEX+6FRZgUKqEk9cjCZTiYBKAPHv
XkmIupXVUbFbEHaTCIk3J66KAHoOGjGFP86LyQmfei+nKsGVkDk+qBqx4W/fQrtd
N/aB8hDPIHiaNIGFwDG4SYPJrjIwlweEo6L6PW+tPVteUPRqY3cNkPKn3syZizYX
WNBEa/gezBk8ojuWSc1Mqld7C4j+CEDb1AJ0bVrvaXd8TwElXV/h+Y/+LgHrCgw4
pj7i3Bzvv9EMhA2ib40wRLCH9FCn1VleZsNqALVOg7tIWbk76f0822sYcFTIENf8
LzxMmaUeJcsmpfN3KRRrp7zbylDtbhCW5Zm7MPXJ5UMYrJyHjUy0XCL34Zyik60e
rhbX8IYXJxjw90QJ5D9nDj+G7cLZNo5sIS19hOjtluyj0ZYE1s1frSiWt8KFqkrc
BYHExcLrdNE5/yYlPvWhgESPsKOWOgSOX0G4LnEbiuJ7tLXD/qs9y0kqnjiagZaP
myh7fnfX2ev3yyVC/V6yNe3rJ6kGTwF6ngiGpQEsu8daVL1xX0AN06uAmI/kXDMQ
cI0lwj2YWoZNI9cgvMn4VKXT/5bqY78QdAvGQd0eSVtMeCBV+MAaDcJ+jYuIZdkR
eqfvGWShNXXkbLVVz0L3r9IA+ktTohB+NIztDfPxFE7C1cmHGQnN5JuxOni66ntI
YzK/SC6+KBIeKpZtzUcEE6ShxOgJDMFRzrwFMCcpquNz3a3fWmuyR3RAtZ4dnLnU
3RlZ/cTxhQZdTyLhmLBwnJI18ye/b9JfvX8rCJSNZo+pe9oLgACcAyAeA5syif/q
IiNEtZ519QwD7jEohK059YycujgCG9A2FRZ3IytH/tqXakUkQMzNd71KfjaekBP+
NqHp/SzFamO2J1OEiNA6oKR0S4RqrogdmEfBvxdZjwcIegAtVOpY01MDll9Pe4zF
0rBZJN3EBgMdfHcBsrLn71dOUMEHTgJSTfE89Fpxxdbrlb//k6IszzGRO80ZNqhB
w8x34sHnkv8NQa2QZSlDc8fs2EOic0s2yvQNj89HMUrrjr8TRoqRBN6COvZXr4et
AxCCasxT1tLU0c0o0YPKGQzxVbVPfuL+ctl5FTKkT4svYcaZ/fox+IYik4FLpVIq
ZELVGGXUaglyCm/s+8+oViWCmYcuko05PRMQU0dki2RfGFDf7TYFS6y059qm30cg
64rBr3uwd41GCag9JnQwBF1GYjqqKabXx9mjHCAvOMclwT+/3eOc35SafP3cNAE5
e61dVe70g56mabaoy2/5XVRsVKvPeSNadbaAXDoVkAUFfkrjEAidJvF0+DweLf1n
fXh3ZCeIsjP9gxsq6FcZOsK0UlchIQvS9ii66OqL0gVckU8oDuhL8FTipKl0AK7X
hqAlMtTKud55HATzdyiE5EEao42yGIa17gbbKE+9c3OOeH+dTyCwobye4417+g6U
pLEBDE/TdbImo+p0q2/h3AIrwJOLd5w8Lohmc+Ld+FC33gpFgz/0slY3F5nHfKi0
QKdbpXH2t7tDiB9I/3yaZ7BtRZqXUvQOUGWgx7qT0BZI/Hu8X/c/WkJ2Qimyh400
X3O9/qv60+GPEbFraBNog0KHiavZuwIi9NO+nGxGWAx8mCt6kB+gw7jmmDbO8OcK
l+i1AywMv8vMjJJWIUpxmgfTVcltk6L09O0cxO5qP5Dk5Ur4dLUl02BOmlAjZPvU
hN6cN/QVFKQWFA4fv0194DYVespkR8nkXVmD3AtP/jKXkhSrhBLOXxDqCqANYTkV
Bf8O9SinEUbMf4WIHoNRdLM8ejlI2yIWh0kii03yeu4y+pvllWayCa2rNHlSI+3n
9va7Lk4dgSzvLIKAhbA2pk1iUhHEkL1w1MjvuUb5iowE/3urXIFrTAoDkqO8s0zt
aKmriCvMxqnUiNFhXaKdotCUXiA2RTEsrEJNXMjxtZRK4Jq3GU7M/fuWMoStjS5+
W2CqotBvn+Ejeu/3D3CJFCKDDvTKNfPR+zbsaqbNelxUHAlECHUx+isaBpFVHc0m
Inlz6LMVY0zm+CMEyGTROZLk+rbhCcGLt9Haynd9oDINK5dDJFkjm/uka/5lHpM7
3/lGy0jLmj82bAzu9JGJfsorj8HdolqQOcXDRa/coDI/uEuyNESLRB8mn5uNDKkE
k4JFnABSa9vXsf2w155vWs/gjGwf9SFIPk08boH1rYAK9M8lNFMGW5iKXtcHah4I
BHIGwk8/S0cYEa37Y9Wj337014kB6SASHr/+RUm/NskH0Rktoo6u4wZyhfJmtG1d
my+QLJZ4tVE4ATg0Ox4GqITjEFazjHjZICx6SMami3Sj3l00Yk6dBIaQ+Qr8cdVU
jQi5t7wq7OSjXus7AazcFqlDdI9FQ9uSCVPf0zBeqCkp7OCX9uuN+DaoJKhCmKgO
FhbkwgDcunxqWeeEwdX6qNwkrDKkGppvdN4/Yee3NlxNrvd7xY8MvJ2XnUJ2F24a
R1DdsJZEnYDIKDiWH6VtY6ublY/EPdsT91Vm1gGsA5yZAjdENv+iybGsPkW0WkwP
Rwo8KMNERExjWgmbbJXBjRPQr8tRWudhDapjqnBfFkhTt+L1iLC4aqWctD75RvnJ
n820RcEmNaNhqLTdYk4exAc+hUktJzXkG/jF+w9di8Ehj/d2udqvjeV4yTe6LDoJ
xrGX+7LWG6uoYyAIsDBTc9ctXsZk6CCn/ZO9wsIOlOY/VwA+LLD4hdqooRV7Y/sd
3G71R4hvOqcc3JT6fme+7lo04E/jXlR4hnfMw7SCoZho5FJ8N9wjFKhMN+TjByYD
F0nzFNyXl0HxGmImsDWxSlhpY9/wPWvrqZM3SMOIVXUEnWrPomixIc64ia0vEmbz
Mr6VZt0ReVlrL9MgHT+7VEY+wKboUH4Z3H/DrjFi1OZCNYx342U2GfhgfPH4YDmB
iOAHJP646sb/JePUx/eqJgSVc8ibQ7dRt6WJvMecSKM56aIvewCsHlA8drDkftk9
vKe0vfUO4pP8E0VdBg4Cd8Yvlu4Fipmh17/VdLwuBbTrIOCyw8ue2sCgQUKrklet
Wre3d6BdK0UV01Tx1mi5KodzYMXEKtSon9NQjMatbZnp42QRQpxsIIn+xtfmDnJE
KiegmabU0e17mKBo1xg4eWF81SkVB4cYFcLNilJ7++6dOvFaTL4DYU52aiLx350J
MkhDUKoWCLpbElJUDVIS1UebWqO3KrBNNDCsx0gzgOn1lT44QfgNM2VHjq9FH86z
OL7Ov5hrjNMbEdmz/vhLT4s4Xi7mhEOsS0sC9Nx7iVWG8qaQep67uh18c8SmbNW8
21WZ8zqihJll00HMF/jvDLYtYYoFCohLY9jqp40LvrQ7bh5l8/i8meKV3GdZpAJS
0JgPk3VleCmAKJwdEeNfRHI7KFATd1bvL6qli8/d5uuNyI4OdJau18Tgs3mfdz2K
BvKULH/59xYPbNi/IYEebfi9t0h9KCR7sFCZPyZObTcibRgVxd25xVQB/95qwONo
dPJ2aJUkEYzfhWP5AUUYbR/62PamTTpnsWfDWE0S6TRUO0Fi6zZlYCGq7zrtR5p4
Y+694Ykkz2YuTthvQ/XkbBQk9axTlLHRl19XFVhEE/hXMUL8+Zz8kCN/+T1WPsJC
vl66hsuTQMrwy9ZzlWx8M24sCNCPjb59mD5xjIAJwdGk68peZDpoCgn53mo728ql
dg6BaD3zdc5gISpb7HwqBVtWbeRhWA0Gh+F+zrk5XaT8LPBfpfz+HHocN3AU8Rz8
3d+e97Tavz7fl0Ur7a8XVnjOlRVcippeqvawz+SyzY0Bsn2w9287Dei/63rAyurF
qSsDDGzF45UuAyrYv/255tReD+yVRPgKoSUbIERzbmVOmqWF6KE43B61IGgngFy6
YFRz+8Aph60kZfqqwKyAj0y+dUB655tyaPJ2saiM1DbTn2BfOLZKtTlBKbt8zCUb
zovVYluIILfM8jcPwdfo+uJzji0ZPUDiYrf7qySmVK69JPV0ou1crCHcK2ZFV+My
au6tfcQEoafCDa37P4YfjbfcY0XlDiqzIcadD9QgUj7YIYUBy2Lz3Ufd3LfVZ9Rs
DSTZFGB/Eq9juzDTBnO/jc0JJ010EUYbsy2CN9KRloATOftWXp63tFRUjoK43YKw
YHja8535Gm8eaQS9RHWSHS+ya5CsIoLzgEvWCQzCJv0bXiBBsjKkDgIo7lqfIOMB
Pml9t2ABVv953O1L0QTSrHnBkmYc6SuBUQLpF7Pwn/VPlzL8qhVY0NqUJAEQYYWQ
6fvTGCXTI2FL7NrWzQdp3qpIPR2XlwRwJhe858yquz2IPJcB1mPWtGM23HmTW0T9
boMasFfXSORT9ChRwWV3zMPdAnrdCKstbzUaGhcXIJYRtpUly6hsnFZqfAeOdaLI
NxFXfCsSu9/uVfs3bLQ6/65WFg0ouxyem/ekQCfEaz1unsnv0NwvvuYp2OoVO+oy
T+UrExKrcZt7fYnhlPi16EWpLS+xNWjiKt7KtgRjz7RpfQ23eUsm9giFzryLJtvK
Bk2hUw0oZdIA45asuosp0E8XCMz73znH/Mscj5D7W+IQce1MPHFinf428f/4jrHM
2IZ7D+R6rvMDusqGitZtx/tfz40PmfuNVsrz08/xdFNpYRYiks/i+UXmauUBSKN9
f3PJSwD2DvSQDLKW9f8ICDnZL3jMGMc+KXvlrOHmcN4UxSQPrRmMaMzQwf1anRBT
nY3CT8ZsYAs8gX4p2bPC7TVYMJI2sZOqtgAzLqjkzCKxj46bW8aSwH5uprXt3ZYH
Wou1H05eBdcGoHXUC3snSDI5/hIe9s9sVeJMr3YCtWrEWvyQLX4mDZwT3uC4JrD/
FlvJwUAcmEzriFX5VannMvjLUcr64r0yRN4YDIlV0SY4jsFhn76Um2xzgSP1pZ2H
0nn41teIY1g/yV+05U6wTh1XwPqmllPv0NX+T4h++tlAR+RvgWSWESRQU//+RD8B
Wm2AkJpLKGk5Q77Y0OVNu+wayPUcigdXb80oCn3booNBcvm12zHxWMSlRwNiyd1S
5sD+akSzyO0ByHBTqr26uXyiK/33i11qSB24PdTW8ZoOHRdlhW6urLt0vhvwXwfT
r1vLkdn4Oi3Lq5PMch5cdP43OqTOHlIJXZu4OnAUxYFHnZziMcSI706c7JYRoARE
Ft5pj6IJ7mJY6hmQSULedIhF96CsFiIWONyIsnPTXOkQvGa3G10Mlgr/l8BTEJ1R
/Z4mh29M3kHmjSCmaf/FVqBhIgjFZIRMVAws4LUaoXJwgWpADgJ6ScQDzkWBOl36
CVpk35rztSeF6t9inrfzQtF4evzpJbJTZ3Kcv9upQJT3TMJLKeZXTzd2G7V+hqBj
K7IQwANnauy+ZdCoTTRSWoBiDWgpA+bnh86QdJGetICfVpd6bUfgHic/omKRvhVN
uylXkjPGa9Vd85vwnHzjlnvramUxm762JrbQh23WngYnnGiwMXcsFzfAM1YdwjSz
d1nnsiIm4/3/ZgSsFkWybpf2JB5/f+xhvno/2slTgn7cexnBNjAr8XeTpo/Rb/Nd
Cto7lw5kN1tuauqkK19dzWVZerqVHVmr1DzcK5z0Zz2ahuWbhosy4xhtQp4Fo7i8
I5/3MNoOoKLIvdMNf1LiVYUwWO/HX5fArTgjPzZaFGER5lvwFNzHupRpzU1B9xJa
C18eTIrbPoZctxY5KZ3Xo8Gjo8bX8HJeOpl5pJaF1kCNlQEh92zQVJswipoA/xY6
9F5Jqukui3UI/IalezxHzFhiC/sDSmbgzxv+ZEiaDYA8T/kcdFtXqZZDHZE2OXbc
ybH63YNZqqNcTolXA1nALdkUyiDDW88jptC8j4DKY+fYGtrP5ZC7L1POQ47uHtUb
8IVenCO3ncihByUQ7RZ9HnN4rX/tuiSGT+XcbPU9VAYjBzHoCfTK9r4EpI2frJ5W
anj7XMuGAuUAnrjwnoGkKS0ffvird02yA0Cq0DVJRZJHDs5Jwbtvo2B2CMxPMuvX
0KNbWDSz7BYNA+qhRWlmxVEzG1YHu7LgzlEEiACbpt2XlK4GD8/YEqvoQMeAecLE
ZxHmHx9VflQeWsmoAyF3DrI3O3PJUeeuI2knQ90R5akGp3shTsKY657IjMEj/Qk5
GLMykQ1uMKsnw6lX09bcDde9MZG2jB7YVI/KIjvgJYytSoIiRCHncYInVEu53TOy
nh1Nkpjstwf95qH0d5QlG4LkSp5OWaDlFqZm023fm/ifEpoZf2IQV/OV/EDb+S6m
5cY6EtGcF1Wirj0HB/4lwzDHFVRWSjEzF1YEzfYJHFxt4TuxOaFLq++vfxEMX5e/
0HTSVVqNniYK8tXvm2ellQeYqEebMlU4w6GlfHru1K3SbnQTVngt6JkW5TSBKu8Q
6QV9aixTagAX5/7ZGvJi3kl/E3QXrpgPlNB1LqTRsF1xj4dpDJHY6ilAtsSQ8l0S
aT6mAAPPOaXcCZF0AtyzlLZbWypRDxM8/KWWD0aDYiHiw8CJteS+UZ0FCasdh9dO
quMYA2mEJo8Fytb7HRrFs+C4sqiZliwDql3JrpFBkegrgqFcfp8hn0QFuDpNFNVC
ZKXZ/rX3QmekiJJkj1v0H3lXWxlWGT09JljxkdHQXCm/wrAELQPymubjjYR9/x3U
gr/ob9lyFvzQ4qwtF2Vcq7cEbUY0HmNEt1N68wkKGAbkZvXHPhKPIiUsUyskoX73
g9PD9wKZfx5NSWpu/tdooX541shlZONvnao/ggAMup8gDmm6xrJtutom0yHIKsqc
HF6lBc7Jsenuk6jP6cbfpSAY5Gm0E5QwvLSRm0MH107ajdhkvg6Qzw6bAJS5qbMK
iGy+2dlHuk/bESO+iPp/Af99vUXXWme0wAkMxx/Ms8LFp1pC5P4H4WGY9FaqtBhO
R85jO33ahjfoc6CfJ5DypQoLtICxU9QIm0/7J3u3rONdUDcxUSbSRvav6K6X4Ul/
3elxL7zFVxyc/DHaTYB3yfvA4Mb+Dknkc9ZLVozAoSCXbzF+y5neqTnys2uv11Ot
07TIqpyu+emxK5CNHVimXi+SVpoXdU1fHIN6kZGdjsCXAkHBTB/PdnkPvJ6x/yaj
ohGIbopEVCjV+dOBzXyDubxNLUpui5QIju7+/hDDcbDKU4HGP2OJloVy99kwHvu7
HotEP/t2SCS1hy/kLg/oX3MdYbiGjm2Ei9U2G15+ChlQPTpYT6pVJXK7oEWj6s3H
q3dc5fng1U4yqDj5Z67LkCMZqZav3vPdEDQXtCHLFiVqrlTE2QBHtLzRNYVYXT51
05q1J6Ry4QlrrT5K4OCSjsZV3cWl9Nr/9IfOoIQZMnbbFEQlvvUnVTxnEsBkMcwo
M+i+aV5NSKDZ7BWHdvGXnJQWBdEi1BYjHdhSVrz24azjgLF7ITF8l1M46xZ9/zQ+
lqwTIxEIrdrNFTOU8lcBVM1dTYi4e3mhosf9TZFeUTg6fYcmQWeXqc/Vf1+u+Y6w
EQeNYbJ+HOQ5+Zt8KPnrwiPcrIkCFwRkQsfV7TIHsPb/CGH+KElSUNXntzs7HK+5
HWOQVmNoVR57WiSVbDS/ygKp6+w7iFHJdaDWY8J3hnCRlhDrKJ3rH2J6V8ZinIm0
tLNbW0gUCqSWN8l0vRaNk8j2uFx64UuO+tJWEE+leL0Vc/ard1p6o44Wb1XIDKFE
7eAuM3SRl3R5EhySt+6xLSL2Rj2DjGn3n1TIhdjG9g7NuTcMSe/eg0Ig92DdwDBE
dEb4L+3IcL8yW2aIspgWp8A6ajjXo+psixHpQkMP2iJRrlfwN5YrLZj/hMMSBeF+
Bd3PSBDNURUuSx68Nuw4NbJeAqH+jP4aQgY/YXcT1IN0bKvHYFuOmp6jPU69XTyt
vAV0OsIxd1vb8jNw9XOqu+v2we5xrmRXOmecY5dp4zx0SHa9p/d0BWIrmbbHnXjS
AdRCDb8DDpAYnzs5d5Xu2UF/N8KYynFP4Cu2oYORjeMx2zpToWynvUrSs1JEAVQn
IOMawGcTQgeGZbarO9Ym9gqQ2pKy07EZjAOzkVBjFr5y+A8CGjvtl7VO3V9LLuSM
UYiiH19OiK6i6u2lU+B7EOt0WmhZ6v0z37YOl/Spz6aumUfAV18gdamda9ynboet
yD/wxu2O37v1Cge1T0GTFMiRonf3s3Dl5p+m3Oy7e5IPd7xolvSK1od7fslLji9a
TczULWjQMWP9Ov911oGctKPLP+gEHnG0Ldza3mQ1etCzkJrzTpk//+CDxQHZZnyh
/c3nYNLUhYPmECJ6tNU4RIFuhgnu/MS6P+byBSbaKQ8P6wJX1MPs1Zz4WwzxDK9I
kvHqrOk3YDgvOiQREOnuiRkuzEFIg2Zxms0HUsKxpE6hHJRwbkEnz9m5wHf1KLzB
44yd3pHG6l635pbLYYOqJ4lA7YZmiofbDNwnUe8xDSJHWL60/7DnJMrRRrVCr35Z
kKskSIm4/gweBXKsTZEEiaOVJRUfQHPzV/ILKPKY9i4sQOv/vZpDW/FSP4equFKL
3BuWzv8uimTyk6V1tsWugVdChrGpsqkbqKwowQwd/q9czyvYQx6G57LRxMNw973W
9uyG8yWaiZZh5ChFxeDTYDj8ZXoSFgIS/eQERenpGNsUElTya66qjYZb9O8ufK6t
EwdoEy4N0EFYL5bIHACWJHCDKx5ep8wBPFpYZysqA6V3Zk9KLP1NXKKghajKEaC5
ksLDKqkpm8zXD6kBuy8YfM3V98fG/DZD3S57U4uetgp5sYVgkVndGoWxJPgYFKi1
P2nAhTaeGCqBpTfwHp48VWju4BNcc46TFDj4Q95kg7+4O33wNSg/WRyEgqJV51ci
WeR7LymoZg0JzqxREahBcuDU8c+gwSuCEAW97vCj1LqsxL3LuaJHuj9AmTHBqdeK
0fV6ItOJf67MdU7jMneYs0gqOBwDXZijB24o6JVYMpaF/HnlRLCdwsubsOpzQpIZ
YqgcbHUvXBnHu9GXNkeN0fSu85IQXsloTlD/Zhdc5mAtOMRecJGxfU40QfoUa2D2
QLA0P4+B7PuM4PExqJk0Ue+ZsPhM6QvVuleuYxRzExcwDR6gJQrdAxv5bCqL7YWw
gbJ3iGPTG5gDCX5DqG3/GRph9FfDcqBdYS+x7321FmXIBVZDjkKAZcTkxzY9PsTn
6AZbjIA2ILAz9BqQ9Uo373QOiPYudAmx27lfg3gCNMHgdQlspNr52AMyrqF9e+qd
Nmcf6ydTnTQmiT8ylXjS228Ie3uAV7IJ4qbBm41VBRcLO8MFz3tU+yW3CQQO+Ezo
0IOwDbfNB6VywV8S4SYU1eDNQ+yUed7Mvh75zTYzQW0Luzo7Kd6GLzIAUatgFlo8
7a/bzDNqv6pgPzplASVz4xWK1VTq9Vl2IVMcIvNaVZKC5bWs0BbalzWS1wYyuLTq
TVCRuJlBoc51lPTHUQ4jpcbsXwRLUiL9NYMI4U+NxxBhHVqFa6k51FwqjCpfzm11
gIHV/GrylrQU+oo388Xab1YmId4oMi21YfXtGBivdDhuS+vx1wwWWS3yDnqtsrxp
9czzjcP0A6ug4A55Kz6uJsG1lm0qm1vobzq7n1fEpDjVBIhp/3GwoKXn8C4OlXM3
at1jVEvunW9GxGsBemChrYpOgVuhD5NkismWuwDbUHg10W3PAJ8yzzgfX89Ncfr0
vr63uLJuZNys7dWT+D1ajJffSHdfgdqzILrYdbZRLWQAfkplbPMEXS+jFjOLSwmF
agUHNHTVh4Wo3o2pGFxs9hFPdhaIjfZXztdKQPMfUHaVhd40Fc1RDo0rxtXLhJ9q
ddW0Z9/KG3QTbbI1f7yZ/JUKuuwiyCxKSSQpQBPTBZ18XFIFbnbpMX9mfKx8v8pm
MEryuX8nvGAddsiz0hNdCWi3HdaHQ68vRpDgdjhtfovGrlqaz3+uQZITIb0Cwpf2
L3155MnOO8xpB002p2ZGgRhDDdCrpJJ6cGUdEczw3qaiusSaUYKaqRU6xbEzSwi1
mDxaZSJ/KH/G4H1ImcPOmunT0SxpjDfaVJfetg0MgaA08ivrMzeVTq7b2aBVY3p4
32g17vrYVVJQPktgoKc2KZZe4aLRA9bujCUaKmCuXdiCKwAiTMW7sUFFa0nFxzXg
B4kyriU2nyQXUIdZSJcaczPi9tsClYKj1N5CyxN9Wc4FCXMdu8U7pCNyJgMe/cEo
7Ja55a17kEBDaV6Kh3R3H7XMVTkxCuKa1abzF7ranH7TahsOfS0pOvNzwkbNo17l
BDzKVEJ9tmJOiSUZbvuAD6lWqaUwG/t03/Kr68QjrU26nUcqXjqWL5kY2yHAueKr
+7B97aZGSMflm+7i6s6I2WLqSK7huzsbcsNFaiteqGYuhMwcqRuDWz9cUOKfr2jm
8mR7C1FHVltdqNqZcnVKNUzG/mi8Qe7q9ppj+7OTJryJUb+qgpwg2/XDsdU+vyFf
BN2pHHy4v4qOQ6wCcTywg7Buv6eDQo30mc++OaSa1Iwvv1eARKX1ap/uCY433DI8
WCHqpErMjs5NCAQB5aSohVMSlALOTfm8GfQN5kQt84+zdj6iY7p4Uc2IPTHpNO2e
1/jTQMFiYsc2GD+PEYohtyQknOxugDcleXV3ZG15CZCGtSbHVgs67P39EeHopavI
fPea/+7j4ztfANsRleXb/K1nnKOhLP6j5SJ+x9xSpSEVGbQxCCE6bXHzbT8EmyR0
1w+LciveDs6SE/OPXMsgGHOjoclrekAEGWiZERsZ0E7wPy3DNFE0q8cFZfDTbBSW
wrxkSw3x+iG+ajs6QEHCOXnQZdjS71bBwOCIXTm/04S9LS2QyO0PHxTfAoAOWHMa
XJl6F4QC3mMABlgK1zfQk//UiTg7yuETe/OrKQNMQ+JFzq0Kfbrc/Ow3KAqC0ti8
5fd4rycpyHf9KRkqJmcTNM+SNOuR/3RPM6hH8XgnqHgvlTgPnc3unuL9XuV5PeL7
HinsLhl9Sivohtra5mIp/BN37wGZPSBGvclhaY0nMhA/aeolZFGQzG/Pn86OihGP
MkvKrhKwyxLqRskeTcYNy2KsJVJ6oDrP0QWo2pEvu0APt2aEWqS3IYDYy4Sh6I9V
VC9Y8wb+6IqLEwQFkgLYcUhzem0Hn86y7qUw1GmsE7aP5Y6QoVHEuGG0c57/f40e
/D67dSZWlwxr68vl0arfo1i6IxxkaZRxePnGZBgAnrycn2qcyFsOiUn5WjyLvgcf
34mvjDPhX8FBKXVHhQvuANQQCN1dFt9M3hX8s1PZDV1l3OPJtuTFg2SedxgAoOcD
86J6dz587KSWUJgCHeG03cVodQAhubvyiOVTBgUIZK0vHB6nG3ArsA8cKzKhNst7
VI6elKTxQApEDvn0wuAsWvMCKX1/Qzmu56d5K5uqpoFM2UvirBUvrUoS1g3Az3qL
iwGLmpvuOnsKz39v+ArKXOuMgwPwj2/MzFQULzLkwF8zY9FqocOmLFjb9gCXdBhq
jIKowUYrJPi2SdIO/bAnYhb4fUUi/4vg7fpLzn8cOdVNauMCA6Jr/1BOp8aD7Ffd
r/IZsWPBbOOxGgcMdQX8HFdjMhQXnW4rJuPn+fh+zGbdB8ljP6Km0vA+CJgI7HMA
Mbl3M/DroVHWzJAvaHl1g5Cw7Gh3WfmYUq8thHcHIfxYYwoJmsDG4c9Iek886Ryj
mnxZO0xih0zMFawuPBb79ASIA+JNb8rQMOeV58VqeoH23Kxr3OyDpHwBNhuzw++r
+CGq8An3nwMfXYsjmeG6FP/9qu9fjcHe9//IG8FtJ/bucfP5K83+J48+lO7L13FS
V/gSMBs9kJr0f5W0J741GjGs5eoObS3+njV5vAn6S53Lj07qm9wusgkPBbRSK8q9
KLzFo9JKLpnHpi48rzts636/0QfaUXLze/HEWf+0blzUlIlf/tS+ZsKAfuWDOJ0l
/+YfQ/6IIokpRgVTHPDhR2sX58Y6yAJaeFAQOQfmwQRqNlyTz44EAWGt0TV5shEJ
aOHMyKf7MdbDKpUX0SkDediiexsNmreSYlClnSomNFiOSgxW8xK3KBereC+t5tJO
eCEusfykZxCM7nCIMiSnPErZf59mGO/wJygyS6EeqaZDq9Lrj4UDOSlTMZTEyXxM
6fZo+WXVl9lC6gxeLnUkNGz9Hw+v+yVQRMqTeQdFj4P2g1nt8v479XUvqwbQMsoD
GGMi0n+sl1brCMJ0z6aLhy0IIVkvIloarpJgRvDQNO5I6yhWMGHd1x8mnTH2S8vw
KfkMKIGFMuF1Vs+RgoTSlAbvnbPyxOsogBadvG5VCnmoNJzf0lx8DHSEPRMIA1Gm
06AyIC1MNjkLXAcKN4skhx74RGBkNUAbMmfC5YGFSfkAUUDNCpl1Je+hMGPbpX5W
3irorCB3nm4rrNQw2iYjGokgmULAEJqknG+TUE5IW7HmlQ4O8injkH2MZoy/D579
Fg1L4J5dHvNTh6Ja3hGszhIfV231ntDLA7pBdkR9QUtbYCxoJxJijpR+jwzoZH8t
qrsvAd+hG0//54dLLd0XZ/bTKIDcZbrPNDaXtk22tFEkfZ6eGp82oLNaVK/PQZIE
SLEy6uNT2ErO3vnKTUdF+0uleAWToIPixnTy5vLQgc8C80q4HVA5KgkCgC6yU/Nn
wyd3Gwnl54T3NoVmXBMj1+JUQt3T/RUHOEEPWNRuyOCtLcGI+NleQYxEtC1/hmDl
+4IvtQBh+SQKl0OQUexZ9yoQ/TCZuPvf67Ux7YyYvja27vKDiMr8N7L9OIyY1X0O
4LbbzVcNVKz+diRqr17d4SDPLpHc73o6d16awmF/EwTh8qrO8FrmFKmr+BsZQFBo
nx0tReswsP2dDybGNnlOzmLkNptedUY9k8J+S+u/Qs7/ejPHeBtShRhS/MJvh54l
7eSY5KLOI1RBD5upzZ1e13GJm66Ri6uKvOWdNTpk4uFIseDaDvd9q3ztAkaBInxq
eDxvBVDir4PCDKtTwf/F5vireGKKXEnnfxyIiuYT4xuWNMsxvrlhL+Dxplz/sWmn
k+rnJFNsCGXWVogxgep/3UdYXplZj1XTEcd9i2iMfmL/1aFE5W2z+5l0q272Z3t8
1da5z+RSDfr4LHPz0pZn/HGefym7Jgl+nV5Ya+UQ1rke6erK6lnmRklrl5Dt/BFl
MftdPFKZHHlqCAXbDFlfCEQJYW7A4tculcXn3Op7sLDP3d6l5J9Hd+I15/zby2gi
cRvAFLcZeNCagsCOIYdTyUl8TpPpZGhR92Y/22CalVQzU5y92iG4QHGsqKip112c
kr6tO8rPIOqucReoKfEkZ7bzxJENU+snePISBV1F8WAPDlAIJ5y9XoCzSatpe10d
75iyasEnMcOeMqf7xJCcPe5VrlRzguee9eTae6Ma6D3sZc2Pag5lxhW3YSD9Dfkk
gar6Wb1h+pMSieDmHdCZAhZOaMinyxGmNKmG6Ar95n6GHT4zyc4HnhwnL5NQuOFP
YNyQ7EXF8x8HXxQ8TT7vU4aiiYvxjojYcSDAhza5y7+t2+s9RsZ+mPEAsVIHGyHn
qpeNjP9NkedvHKCE+thlTH1XpeLgF5qDIADuprNG5wWisgI3NviV8d3Lnikqi7WD
w0jggWLc4SFcAhtXJ/421Bah/jt6WiJQOwFDevsttBvVdbp3ZkFIQV16NrIvDoV8
T7+wcRJtv2xm1788hkHMRtf4YsoPc26oeAj65upI1dd6cJM3lwdW4Dg8JkVnehXm
cZhAvb4IqUpoK4XHG60Tkw6plvjONDrHKXjEYwkWWMZzDIw6LicP9wRPn0GgmzKV
X945lubch1QaRIla4dy4Lo3vgvppzeZEftA+cSiy6NqHVBml2BnKBOHqO49mBOTf
AmUmeWppUwhcU5prsNBt8ROIVuL25/m1HGmX+enMabxVVeE6pnrbIIYcbWJ32sxG
ikzp4qsnuJWMklC2w/A+2RKPDH4JPhomXgIMOqdU7A0b5GsA9oTmJ+2xoE28rsFX
a4P3I9yczwuGBx+vv3k1wV3wjKumdMYuXzV5HIw5sh6MNanJWBq3T5zam/SQFTM9
saF21Hn6eoEQ578j2ZaKMhabJJQhKvp7j2MjHFvI4e684JeUVJa5PzpJcsYoK4d+
pD3dGIFw1ooJ3zWk5evfQ7s9cx2IXgvkm1Q602fY4F57EPWIbHXy159zdXTFtY02
HH5JqK6amhFgn2zkQCFfOlyf2BZMkUt08HPbmxZb5lTFNz8n51ZpGF7gGXOUVeeU
9IG0Rgu5ErdlXaxrW8+x1wUSfgiYCb2coFoRrokowBOSkncdJwqhOC7CJP9Qu/Q3
s3y2I0c+1MPr2AKD7AcTdUmjp7TH5RrY51ozn3JU4NkE2giee6RsM1pQlwQ0En3m
40bkVAtAhHZv/2zP0KLMQ3g+xWlKTUYs3ESkOUCd1h/SFQF6t/uPgbCFGifhcvUj
r5Hdx2fRmPk37RQMi54Ff621OSAH3G8GuVVVhgGH2o8E5rVX5VjfrsPquzfl9EyI
QrJtYxPh9CDrIdDEb8PL1xWABuI3ySf2rs+uXoGL8pinJwwcZhWYisENP9TdwGO4
hbiVRBdFMyXrG3tHwhHmJmqm8cVXQIyHGOhUIrCrPZ8msIjYcPa363PXXhZrFNma
3C2uOp+Hb76Y1o9fXy9VUpOIl0q+m+U1/JMEzJEkDQepld+KRfdOVHYk/IFecZqU
gLm642JP6cN6554SDSmDtXR9ufz45KkZHdm1NlXIfKjOWDUA8kC/93QwCeA45Nyo
DKi0VJ30RoQydyYvDsxVb80C0+MEJp9j+6S95V0Crx+i5baqha2/oJvCWhJJI9Jx
50h5Ir85OozmaRU11t9og/AhkiIXtV+ND+fQDw/90lhMi3hvcC+EyEe+Li289dBD
iQWpp1tuHPciV7tBDOUcZnP/k3mabRGZXf3JaT6pYkmHKzmgYahJh5HIjLOhKdhd
l4f85/WmPlxs5Nhe/U6tv0IwxKrGo7XBYzqOFfAjmNH+2vBxk7xX6e1Ljnx3HD8B
CTItu9Lkh947zjXEdtkMlbNChVOV4YmxbGp64RxbIgDPcVTmYADktbS+9yMmV7Ol
Snwlxyas/k9OkFWeNqUIgOtGVkVLNPwggK5fnhYrwWwMiVy2lYEhPDYQI22XshQo
rxEG+z0SXK7qxIB7Z2aM9LnrCnuamH53rZ242Rum82inHOvg2BWipKdSRl+hGehR
3Qi6aH2QvwdIo/snzRsOj2SIQn/Exm7mebyGZIV1gUhOM64L3UhiMLzx2v/fOE5T
ZdkqjCtvoYgtuTt06jUp2K9YLAze3S0d/7N4wc7qIakGyOhRfRbOfZZ3rt/byl/2
Y8Xft9BYIZB0RAvtJ54EUZoJSO6fFGjq+RGcSozfRDdB2J/sLMTYMHvWB1NYEV3G
nwRPHrbOTaDHHHrkP4D7sGIhpTSehP+2T9d5uGS1e4ujxLkf1sZqHBESUTM+x0Qt
Z5Bbks5qt8JdPuv6d9TifZoR2E8qu5hn0/Y/pbfjXxkoJimQa0HPIMBNdzvXH/cc
KsbNF2nIMupX2w26vzZ9rG5CWrIGxGZ7y8hf3kfPlFBOeM0++f0DjANAdAW1OyzJ
cNI6CieccFYE2P3/UKtOX6mytC8gk+YqgRr/Jll3jGf1HXAG3O0/SkyA7mMIqX/4
8reA/D9qbh59hWSqzD1lB2EBr4yekrSjl6+N88xzp3W9UAhgxhsIIUwa9SVsQB6L
B4o9ewpi5poXqXx4+LX4xi/rSrO3sB2EPdaHhr3Q9EbVdpVkeGvvlYCxy8khvNQV
KC5H5zB4OC+alsfUalxyOnNZFazyhWKeTo08zZLQ16CvdRpgEgwBv0IsgnDJkDhO
8/RFC0KJnCjnBbVon8+9H0pTvhvqJLmIxUuKjlAoWwtoKjY+IKjj7K6JTI5rs7QX
VSrw6+T0dzDf90iraQicXBta4vnE35Y+I+lnIUQixwkN7qpH8DVgMhzig9ktxBxi
RID+453b9PXrY5cyIkQ7RRvNhfqf//b1NUX/Kd9AZA8f9nbndbmchkPi5viZNcdj
uU1vpPb+ZWsnBHlm62aRuGG+c8X04gO0TJnxciki1yFwZS7BkL5lEO7uKYbelTJL
Mtp/bPuFr0t0Zl9SMok5PXkW6/1xCvlsb6RVCU7tCua3EdazAj+sIiuk5/+e9vBB
gBmaH4ZywZpznIBYk2OgTf6WvMo7OykN31otEnJAJPjyVILturDUiDVvlZVtU0O5
jZ1sBpvrKi1Z5u+G5iiYK7yoEBjUlgiiN51GMHjWrl7sXnIozGnWnmchfw33gYe3
3qdw3nhjv1v7O1uM7yUKk36b9BGHue0I/BzQnKIjy7zJZQg1c1EFXRqIenE7c9GD
11rtaeEqPdzsRrjKuthVH3VKNHNgew5UmSVbnsQ5Nok9SIORBJqHf6cFJQh2qaNY
RiArtCylxoLl2t2RblyJ4oFdUPQ3LDtfKpZD6Lcf0tDyaBhGjQ/8rY3mFqztguCz
VWEYUKdWlSxJ9G3Qe+Wj+gn+kvv8jlDDvFOzaRZ5J25Nz18wSluZ48az7rE7TPGE
B1S+b8sPC0t7DduuqS19SPfYHSpsZ5bz307+HVbQBini1WmT0KhTSF08usaTvNVf
V0kn6nk8WYM7DhGaZpXsV+7yFm1mYS4fKzgqvIVD6SEMbs0AHnGI4DvQWl/meW91
kAfI4QBi4+hlivDRFMUrC5Jpr8WIxzUIIBEDCDFcSap5BY/wvCHkky9zUYxInfeR
jFVm+C7+hqzwoWJwYNxNXH7T+O3vtt6O7KlsrWXaUJJJUMqeGdd2wHNoA7w9m2tZ
oDROe6JjpugM7Wgav7ep+rjwcoZ/fbYqtDSJt7R3/gTGwv25ySgCNoJh1h7Mgi4z
uYUxgk/JAWwcd0ZkfOjFpo+ygqFJEPNJpBQGGB3i0ta21x8g4oxIM/FcxE3/b5e1
3xpAwfmmM2K4bLjYGAoQWH4G47KXYviPuMxZ/6UHzA0VDj21aTzBbbBh98/UjeiQ
wQ7BbxyjuYmIiU0MUFinP3XBtcF7kgOlsNIdMQ55D1i0Z4sseGG1WSdguyCW4u+L
GsipZiuzUV/BN2Fyc8D3177cW490mFGn2mBTh5lIj9zuyx7Op6JhrE7Hs2uehUFX
AWF9QsV6cboyv1kiH0anmgNbI4/Cq4j3eTH4Q/djwv4f9v47nJvVgDIsYaTWEV8X
vmpmInPkiIJdxG/MQ2VR0aO4JeHuwydO2/t2clvhzLTMV29z6bueRGEl/c3SjAYu
HXWQvwZJ+Tanmhy0UOW/5mzTEg6x9rJCOvZmQBNWjvqY2qAtrOn0hsAMPqyyXjWD
JGcWDUdDJYqRNva+JZWWTPk8v3Q6db17ZiXRbYo2q98QiHtWxNqqFTfbhmiaPtz0
3+5Er4bHhMipUzKgvKVdvyX7q9Nd3PJxGCnJqKWMPbVB+OZNX4+eoLSIfjKn9PeU
24zt9GicsKgBO5fPpG0IkehMu2RDEdxsQd/pLm7Nws/+fBNlCFcgjg8mQAjvuTj9
lbWgpQLhkM+G+gb0CExpckJd6/q/XEnGLzr8UM4lie6RjNf0swI9iunwdV4GbIpw
4ItNbDNCclhoo0yBvVlR6dT6YIdl3VQRgjXUMAn0xfVT+fpXzEFgUkn7sQUwzCjG
4n54bjBmppsWLjFyrp6QE+K/5x1FgkLju7COefJBTJRrDc4nuNkc1AJ/cWBfU75U
funkhY/mNX7w2YxeGeEiBYSu8smajW8QiEhsLntgcmnLhwvQwtNSlufoF58aaXkP
AlEkuaPs2evDpSx7Vzk1XY3dxzM61hnszHLGNOYwFci3xYeHWdjbCoJqrAnDmSVL
7KqiZsrnTrWE3rAzjpzUIHMD02y43IfNNEgYy8VXJuI4ticJRSrmLbvdcm45NW7a
w2W9/a5uJwpNgN4fCbWLTYHIdMBmmT2nftrehLMf1C8Znx2XuqDw8Vzl7vZbhKgc
HeiPMHpeq3BoY+uI0gVfEIilVfiOREeQDgDoxV30RCinH2JsZRtFbdXoOJsyqNtG
Lvs28LUfxayPqnrxtTPovgCwfo2A19GWqsQ8noBJbHiRTAcyijTtz0zSsfiBs7Lm
MQrywgnbJcsu39UO57ATZ0N18Nlpdhs6iG8vPeGygUr5v/exIq2Uie2SeBY0QEM7
lUad9qk+Tm4ssXirxHMchAtvsmgyAekrd36YTcwxRSA8YecAh/pB2sPYRLIPQk/y
qNscEiAvHTlQnxF6gC9rcDBbR+6Kha9TE+NsJiU3V99Xa8chMiZcSv6fMbMNYnbc
CMNYZ1creqcGxxO+xDHWyWHfIt4+0wk6VKyKJHYZPDkGm2vP9rTRygpUDtRW9rZs
ftWLzhwaJ6w7olIYwG6/WCaAmvTTMNOpnL+BMyU6va6dX5lLlbpottyoU1i3nGhk
ZI49h3DEW3eonSaGZ+FUPqkUTH2yRDHf3r6OnCbe0CoyFyNTSLoQNxuL18yN5nxM
IDec0g1Vi+bmec86C4whSqwKJcmKVi7R5P7+CE3jnbfUxZvcflLswkrxxIFGeTip
bJ5fSICzyLwCk0wMI+bvhZzrutNCFAOwRFqA9Evk5diDLJmzpp5fSCrrhibEseC2
DlnNKmz539UIhpKljzX/HPVq2YSzMsE39n0UPyp0ZgAlbnP+QN/toVixcng92y2K
E3Z44EJHRx0P+JuUiXixJ96xnylUTOv5AgYJsqAJ1yLE2moZvTzoq0DRdG1LBfK7
uYYkA68fV3Zx/3EXChDCnQ3/BWas8PnK3HEhTilMb8Yjvf4Ch3Ed4biZuaPNMgSH
y2t6XQs7zfBmNIn//D9COzwE84wpw4fimDThXSF8Wd6OQHr1ueRvYc8dm3Lap+hO
VXnkDMirx6AKWrwIdYQjuNPGKbLKLRx+TDeUnc97s7ZFNgvC0pgPYWuulEKvfgxd
x4DKWdN8A/C9pXvO85+u2Pkgh6EVr88PL0IyZUz7bN04r+6SS+W+HXdrYDq7OVde
+pbQAKxdwWV/gzSIVAighIxyTqj6fdwSup2TAHyRhcCbmvzrHo0ulLsHMSlbDmLt
OaGYKJD07HOt/RcDn0P0DZqalKn23jAorhUOntf8hRZEn6Iby28iihw3frgvkjDs
gQTLD/xcm2uDnzQR3Pf2jHG+GXfKm/vz25OfixixFE/n2Ba2tHiLtHwIHbK2mDRo
22bW++k88XXQZJzSkxCbr0Zk8mN7KQJ2fa7lUClkRj7u/lqikPwnosvSKYTgo3JA
MdAiYvzKylUbSV44hEkUxManOyG6hCTwT+9Zx+OnuKHvCUxLj7IL6+QtCD2Hm17/
0yLWnNfQSMkrzsqHSQ4pxZXExaBoKZQGqKdGDiXatBpDmaoDRZ6EYWCM4/SdkT9r
npaYy+QeBkpM5qkxzAcA6K1cAfspuaL7Yg4x+HakrVNGF53QeNB3eF2zqubCMQGw
3DS6vc4PcuH9hSq5iRanHHIpiIvU3laBuVZ9jCVNQkwvn3loFrA9geMIsOgC/JT7
wpEpU7+jZ1Pu1+IZen9DIC6krZSIl7dyzsyFR0J7RDxclEFDqcvxCNpdFP6R70ZZ
kkkdwbZG0L7j9ST0Y53zC+fOGdY6Ce4cTRTYgrH1osv0aoVRA40xdKQrD/8mylCT
hGdF/+3X0l+5WHAai7OfKAm8EZl4izJHTfSw2eAwzhAB1+MbhBmHfZ6o9+at1Nht
admcsSyzrHJPy1rqb91bDmviyMukLAhoqkz3grYVcNzM084OuxVuQmpBNE6A00Kb
PqTlSsZBeIW6/NRce9uIohtEHKu1a2buOAcK1nlBXC0FsiZlOBMRHt5SwByxCo5s
c49G7cTY2mdEFiMEC62SJ7cSiKTI0rFRZXplgjgyKHztklKeCSomuU9Ql8nbGHHW
HvEf6fJrqRKOeQJf3L1hyJJSoFcqvHkS4U/AGdez/hRlnuqJm7usq5yP98CTsnVo
rr9kBuleREBTDajQ/O5wt2Uam72tAX/PEBLVReFjS2qxwykkplFyaDjDwUk0xpjv
uQSlmseAqUqNyQjPLY2FP9xvf4e1KLbLtRPv0TOf8bmZ6g0wXuW0LWOW8golxOQr
PbUXjPI/pL/znzv15fKHcYxLLU2k8vjxZ/MCSluZuUdTaIUj9O4JIFiT/kQXit+y
7B/F5BDjb9nmvWabnLZ75pRiLfTefi12eTkSmdC9kWV6up3cDHC9Q90f6tOTeI9J
jUOq4ofqa2D/PLoT6gG6ROWBFNgJVXwX1MfsAawiUdf5KalSlMvvN4bGD/YGQ3qN
e07eG3+RGVP1rSPzzwYYyDqWkFIc2iFRON6UEoIS07S+AtMdEe0UeizlIkP44m8Z
mFBW3Uxiqb8qyE8ESMTXOzQkNvSzgbrVoi44BBYXrRMv7C1xeWrCg0RR4LHQA330
JVUu1lZgenXv87aNHmpcCuPMdCTPuqLZJ98c58nepxfUL0NdBOsFHBgWrhAy6ISn
uCbn8XDIaG08Lgu0aGjupPngM8CK2/GoNcmkPgja7PTAsC4Pcdp1nrM3K0Aufj6s
T+zUP//XeWs33Fh/1ps6JsrhACUx0UXN4diuefKjaiFjjpnoYnRAjTM2fCRyjMUC
tMuU0lxwBm78Maa3UGv7g/OcxC+t8Jd0IJ2T5OWMUomels//gvSr61myH4u0Qo/i
dSf+15wYNx9sLIFc6RxIjjZfxxQJqdn05xx/En9UobFdHRUot5ULbXCXLXw3+Wbu
JhrfEThXF+hl9bJMwmaj3EYaEL5W+gxR3ZMPdmjXpcN0VM0mYSf/pj9qgeXJWmvQ
0tI1d3OfeypO2BducLslgMyfIoEy2aMhk0kwq6iIpGyfRGsfrKv03N+ezU8ChaMA
1XIfyDflYBciU+dBkvAbq4dRjqzLYpKsyibuS/qxHeP/Ybnhu2lTu8A1bhSyPb0M
RcjnTHi0AvvDXchH7rRozrM35aJGFCZLMIJuct33Yu4+BRIjbqMMblDVeVClFw3l
HlevToMJmrwLlHDAQRHyauU7WlCdAaswybEMGty1oZoicdDK1mAM8y0Q0ezsqY8I
qiX38ySJRTEmqSt4Rh3IhBCYugHc2DkrD7ojTfEAqpIrXUqdcaBNsiJBGFJJkFlv
uwMsMWF+1uYdeFfz5s5ruq9s1jrpO3jSvTTOHnB7QEL8/it63YjNphcaMgsnfhVd
X51LAbyRjQ5xYyN52xwM8Q1ogTSyTFHzpdBf+balJfEjjF4yxEoAbdA3CQX/fx+4
UbKVwNpKSphg+9fi4Bz+T7sqQeEwPCJKwVL+tkQtaon20OK4k5GSPE4qrF3mzFqW
kuLl8dKv0Rft8/qTLcDF95X7p4jRE6EcG8eVJW6zIYA03Fyj1Md1wTnk0Z0RU/1C
CgoPtMPX6CaTbH2RH4xZZBTMewA9VUetwpyNTU7jKL/17+KKGXqXm5qSgCdlM7+E
Gd88JR9If6ie9+vN0CTxP0EqJYTUPUUj41AbZvgMDMs=
`protect END_PROTECTED
