`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Azogln31o3jepIFfTUT6qrDLQCy7r1HqYf1WNPxBTXb+I9z7dEexsDJsaLCmdrZ8
DzW5xbUM8Q3KQqgKZ6zOZ213rreIt2RSM7C+W4uuyTgPnSTeVO3k8VQdRcoxMkrv
OQOo1OMe6JwjE4WzlSZD3snNy3jCOSGXILA0C05XCqUrljk7U66dzjUGsjOcS7wU
vOLsu+UctHV7AF7Va5Mg7cuDIlQrZDTU8i7/VVXsCYxKopG2jnflOlw6aGQNV8FO
O17FX2+MEneMOc2dOPwNzLcOwaaT6bGwE6RuQvUzGE1A1xLF0KW6UHSqoAiNNcBD
H7A1JiRax4A3bdj0I5498Dl/KDRzAHKOz0bGMMZJN1VMj/Yykc85kS6qY9JFF9Pr
tgW8spsw7NoggFq96Qsf837SNE4poP2S1CTrhVnXxN5nQWzDTu1ui+ssU31cIJiw
BdoaOPOaxz51sNivhDmKjA==
`protect END_PROTECTED
