`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dhl8p7hpwM9gdeoXTOHAsKX4Cq52jzwV/lK0vBHlZMem1E7X0f8s75OyL9lvD8FA
4A0Pe8PaxVjpLcRLbcZ6LFyc0oY6IhIYmnyzel/O5vb8JkAFi4zuXlcOCdhkDKqv
F0rQ8f9cnedB6urR2HOgdGpnbQhCNRyUH6FJsrTEnsv1KgabJmIGRvbG5aggFzjO
nsCpbJMLUvmnO9SSHvPw2oHE7o+nYeLFxva3GdFzmBqtH4y8VY3vIB5klo4IgZAX
C3GrL/cPzoTIuP/Sf6HIkzJsZ/xwYjAJy3RRDN62xO8TFlOdqdOmRzwl1vIoGy0o
bc2EIllliBM+WkSXfoXhQPStu4dLw0bNhuinvuy5kJNjqzZLvhJoTTNuMRGIHe6n
lfqnIQZncuc5NrHy96lu3msLT7PYglneSAHgxJ4ye5j4m976BjoTsd6f3d8AnCWG
02K/sypWgZDB2RtzLthURXDamvkRK/+opGxfD3t40BRQ4kJzaK2TuAfW7JTxzpQ+
q3VXAqq+T+7BgwlMObD5/+gQao4Fm8KMxZUkJ2Z0LSqjh6CBCP4nzHO1aSRYhp+i
TJIiot6ycIeEQLSf6dEp/VcTwW9C9p892Q0GSXJt9G0YBaH248y/StSie6iium5P
sDidhoR/dwU5+UPciMZog7+n3ljKhwAZfY0NIQiJpS3SoHfSBg2ap/r/Qjdf5jQ8
b5mf4M1b6HGW+A57I/z9R7k4AkGj0QJ0b++mshifQWyEjkBgEZ8U7W9AtMBu160L
mMjzgcQLraI+0c9NiFSjGWitA/UPixtK2uNRQhm73qV/ZZzmoCHBfZWk9slDtp+P
WXCBomfGo0yFNmJ7VKQaZW2A0ylQpMmM5wDd4b3twNqO1Y4kWyokfnB1TFXEDt0T
0jYd00UdR9pKyPwRNhKSBBl7ZeLzH6BakWRnoaibYVeRccABkMppr1uH+DIvlplg
CvoD2Yh5/DjrrlWHNT07wRkh3MsLWrZvu5GRJjxCQAkK9oKHBAZyZy04FvMrfwUI
SRx9Dr4XHIn6XNU5OaKpBMFJakAN5ajvFzRr7CtKUMEdhxitKkkMGe4OreJQEL8m
DB02w8p8lDUUlLMikpqYdg3r2cDO4I0M8FxJnhskx5ADq2smVpfV9+COytFdcdJL
vCvaAHkRjyGhFYPq3BuyiZ4brwBxxxL2u/FItB5FIPVDyGwC8F9wIlUmL4c2CXwT
PGUJ5bmlPJ6uScNEzeiSvIYYIwuznrovn6KcYmShQEGCLuDyIWH6vE9Oyclsnd2A
wudnu6pvI8hprgMNknIGwQ+5ciebRtd0WlgQRnGSWTKn4rXNSiYxi3L6lxi8tFDm
tGebG4rdDOtrQqxt98tSn0I48T2o3s2ikm3Il6nNoKtmTe6tmR6ML4ymKEUkng3L
NBspb+BKqqBf2rAAwol3qohrcIsjrVvRugcYWRbeZR6ItZTvPFhechqidbU6sMwA
2v+JOqnic4O/CJxCPLOmegtgIlFN+gzPyhM6Z/S/7n+mFo8oKyXnABl10ao5sTZI
DDBACmvNysRjWjcpfngzgScNWnk84ecKF0diN7wCB2AmJWJXAc3py5kfAEcH1ljP
YXzRRyeDiDWMapspB8N3lmvHVn6DDOCWvxxkk4LPi9J6ybBF1t667USQSjGaWbeD
+Q+RJWT9NSvsTbQplDRaQIpBXwPouTOTwSqzh+OUoGEB/ss6INl/AFhE+pwAgQ6t
g3kFdg1oID3GzNK+SC5kcEOkCW44DCmivphHNtYKP68Nq4hASshBbDICMH4XnVAc
afNQlZznkEigLwlQOxIqraoj8680hUA1N81HqpBuvSDZxtjlqnOXuk4VdGcpORIc
Ks3TWHVU8VM1jI6qUTxHWl9JpNB6leM45/WV5zWH9v6YEAPpZe04rXiHPsjElNKF
7S2r8bTgq4cfoKYKlhKGtyb0OUt0jdKRcTn77m0eWUd7cEH0sWp2k5uVkMPqixRg
ile7OOLVJdZZDK8fVz0330sGdIz6F4g4vaCMlldXetkedFkjGoOnvAWrgxl4S5/T
4StWXy1k+Wlncr8IPkoTHOfTttlkBvmk0WGvrBfM2KDrvhXSFZy8tSrsCtrK0iOm
qp4JT3QKyomPmB0Fat2n0rd0jccy69CvOAYNrfyDdG5gNWnWNDi0ngntfNYRfbkq
V242YtxTShM7xdbvVCKG4xPxuWMJaHH20S7npz85iZ48XvVYXiqMNXu9zjj2UqpT
q6lS2fE6/Lx5LZI2IKjh94S8jCcR6I/BpY8AfdjDjAjhSBjaA7ldfip/mkMYxWYJ
VKtxTgVUpw8VkJlGaEoitKZNDhnQ7T6kt7bTYXBO3Fzg46tp06VrQwSDPK4KUGUz
PkaUMF82G13i5+IciTYlI1Y/AIaUqis7btatB+t9d717v5AgerOkB+/ZKNWPIRvy
1U2PSx32FkdHr7ys7LdAk6r8CH+VIw2fKAsuqumn1chrfiAi/JplJVKdtJaJ62NS
4R/D66O8SUDeQ0bvZSFphY5EhTOlzuq/YinWhLOct+8=
`protect END_PROTECTED
