`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQZBc9R1URzKQx38G3uoIXAgtchKRKTxiqYymF0+bgi42D21dx/97qMLxpyx8Ufm
jKRgz7zi+1fINl2LYcne+JBo+z7vSaeJnu3isJIRYw8YRzAhC6b0bNOUReuy2V9l
DBaxiaYO9nmRKvmGOoLCOePssX+bdyOFuZjGbEyM690vJ5vLinN5DWnGngHxjN9L
IqZzLGnFhIqAE6/arA/zSH9Q20H2gwYIlnP6jbCWoNV8y4PAdE2uZL+aSghlmjwU
6U+EkbQhQb6h9MRcBomoXp+BCYZuPVsW5VHhainXl5PCjeyEpvCywF/uYtuAgJex
U2BjxnjgvyGEgU904dZZGLSS1FzU51ZUzndQtdnTyyopR9UzW4Nwtye/i92GTlLM
nO6FoEdhq/BEJheyjWjF9BucO0Thev//FjyS14BkFAg0MjfGA5zI9qRgebUNflX4
y8JUFHmfNswGlFsdD7bBu+6sQIuIR+iMqp/bjWxs7OW5JfOZ+UWCvwtQMd7Hi+o8
OaF2q/58G2CLUpK6rC/0WbySYlpTiyDsGx/8szCk6LKMPmNugdjmZHpdG6WcrSpT
ZjOuwvsXYhNi0f13Y2JLr8ttUj78MGLFmnyPaqufgBGXLIJpY8qeOkb6gKaHEowI
05Rk+3BfNplglokpsx8OjYDf3/UhMnZqPSJ9CBWlaMD2LVhKjTtEOmpT3Al6bUX8
1mQ/hrkEFF5+KsnzVpMsWWf4xwz+S+lG8txxx8Xkr6kYDCQgpJxXmTyaO4Z2btKS
YIMOESdQEe+/mU12ehM+/Yg1Hv9OfbfyEmRAjOIHsgC7LDUJaoVTtxIBFOl3BIBp
0GM8rQblXnoMP+J8svhA/sYObAjUHzek/zs5d0Ggu/c7lE6o5l740u+EZTRr0JfS
sNQhlZFY+lky8oJUHQKYRVXqjxRywILt2FjH0oWbVE5XDDA5he5kHvnqgkkyWsgQ
fSmWPUpxttjIlg5giKnyrcuF3gqzwO4QTsLirkoXe0MDkjVVTk0xhvo2fr+egAyy
TYgYuvXKCqSjjEdfRvciIxG9hY4eZus24UwQczlwNIpjGmM5N8qmiVQxNTekoKD6
ZGsS9LoNd+mGVCq1RxeM5MmAXQyWYSE82ialoVR44LHDqo/nHvcmOIhhAI7QA9SJ
sED+SqyiNITXlFD0zxo9PkKu1U/MG8sNYBS+qmrnGYxC0I7hMRIs1AFC0a0TkH/J
GiG8sGlyiHds3GykmYLSmQSCu5o9YZ+6HAaAJMyI63NhZYSJzmUzq7XJllOY1E3f
vISGxGWx3UzJ1WQO4bo9wywFSGWBxP2jAl2LFe9vuqAjq/gMyYDKeSoLHbSDx6wb
MTDviGg8jvnqeZIpsN1x8/cIkg6RVXnM6st9yHYexyLVpkFs95srFAESzJFaBja6
JgBLQ4IX7kvPTe52uoENDBBkSR4XOs9pRqXvdRaXtPNConslV3NIz0H933bCpu9O
+egLJLeH+B6c6ks+SR7ldfqNwLwd4Vx1TIe2z+BJghsl5qrEaH46kB9lNBtXel/M
+iedQRHRUQXYvpFQUpdDDYjN0Ibyb7RG09ffo/efcBV/Fc+Bz6M/Sci5chHRIzJQ
Gc/R3jufx95SOdyxiYrjNb7YrTWsurMVh6NJiFVvwiZvUOWQlQaXcvFshzVXTr7a
v2AenULoo2te2cFIOeiKzA==
`protect END_PROTECTED
