`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hI7k5X/aM87fpngABuKwTD/1ebPa+eFAAVWioKHc3d4+LRM5gJ7cOurFABEkgi9J
dASq3wqidBu7pE6Y1Zvolnj0IrqfvfHCCVgCKRas5vEOHkpsBRC2dTWuNcxc32Kr
LLUYx62mZ78tgr3Y+MM22kvrPX602u/cJ2rUx1AaguuipKk2Vq69muaCRPRv5/mb
lnmvoTnAfYp82ElN6ib7tY8WFJVE7WF0Ij3Iay6+CN/B99WYPJ9ld/Cweja2BKak
uKruqf/WEFOq9LXJ6z7N7raJ6ykF0vD5lmOiDl+58gPUpaJKNmzG1m03te6oEBty
8D8nGe/QR5FNxmEAhWJSQFWeO7pEdRshCfTIMHplvR543uQwaSnXcnOgyejyZGdR
Zrn6quM1BUa57pbDMqzkiYidVrUViC9255oO866YjERL9SIkz5IHeKjbXVrvN/LW
WAg/ZSNpEG0y7SpeEfc1J0s6Lou2HE+ByqnWufyxw9SfcHa54ghQDxRYjhWwLwhz
d7a7uGxmnKhg33Sf+nvhFvAHs5NDJLjI+drWzN/3E+UTqPLNk63okZenzbSflpcK
fCnUhgOMRzfD77C55t2yxgpaAXz2o6iaWPZGj0QOiotDql9F/vgnBV5zumhuxanI
rD6XLhzMXt8sRxHd56od5xU+WJKQc4TsJfheCcycI6gcJrQ24YdrQGB/G7M5u6uY
jvNuJvzGCq31s1G6XWWrmNNUWYK/2BUdBXxjhWtB9+b0iXW5GlbatkDxA4PFHqml
PKpFsjxvmGs90E4TuHvcaZ3T0+/mW1I8HCu7c24yBdWDyatVda+oH9F2WMWe6H+U
4rYsszLFCt+yzN9I55W3Cj2ROSL+0d0IkbMOucL4aDkSECOAjLSIsXTfOdCLT9HL
/1fPbM1pBGBDh8nlPHgI0wU4b9Szop7O5Ln3Uzv2dWrWuEYRjPbGYgP9FdS1UTle
FM4Mm4zRDS6CXsMqgE4JriTkU/78LBcOqkB/ImDqsyZ5WKbWdFveDOD0OCmHGzfI
n34trgOq8BJpZU6nzuxLGOj22Fyb18duNQ4IO0AMgmw/VwxK4Yb1xoTR+zXdg0yE
8qzYXgazZDdI9zZUYmBU6s00GElrNUovwKMtKH4o1d0Tfa734MBbUsxAR3R7ddS1
waC4RJqBsLFDQ/mEgHIcFp/PWhnxSluSenEg+YK0035CBfllPupzb9tRPQ/WrLf3
HLEuU5RWAXJ+pNzoRGpUb9ujrJSW7PzlqCkx/62ke8Ai0jq9PYk9ns5mm1gPLVZO
RdpLwzN0yhGbItrInROdLGkcHjjamiR0a0u38osXmpuxR3yukHR/JOTzQGJ0TaGH
1N7l5P3ccSKPnsduxvrHLxXJUWGSVnTawluHpy6k9EYxzQKi7DMz7hFGOsn/RsLa
06XTb/lpreOH4Oz3Mgyc0xm/LuLPPip2aoMBn/RY1MBaR166XPzbuR5dMlrj4HBv
/06KBBnAREo9wcVPaYAaMijo0x1H4+2gyWjJjmoqSS0Sd6bL+EAEvI/7akCbgNS+
SccGH8RYnQWrsxrdqVOTvhU2Za5WfdgIkw5lrrcxmoBTkYYIcXcoWG3R5/e4xBgV
xbEok9aAKO0yQOdqHlFM1qMNXUXSdG0XyAWaKHKoNtAu05CKEkBJYqK9fTX+foZq
nW/IPOB73IfzkWCVokQW6wP1Ok/pZJoR0Y8c19+3vBHSWHw1qzrxF21sByBnaJk1
JQwAOJrGd/xYg4FVKyzS8vRl7cmh8PkpmZ216jvfBbAi6HgtO4gw2vyiKcQGbQXv
LBfdL87EyDGIYH37AnriSikh0tv4XITBpvV7IkJ+i7/rSSaUVZ9tJC8PTGeQBM8w
vzpPV+YKpBjAR8M8A4ye8RNBrtJiywiQtFvyuTwzu3JVn7UnDq3i2YbO3C21ZjwR
GQrs56aT1OKl/PX1yPZ4AiCuGp0T9tAQZrGTJhLmB2cqQq8fIPr/alHCV83Pyog+
3GkIn0B6IyoNqjHAkBXC10dxRHO+j0kbH8aIvFb6IrwY2k75024c5LP9qP30PTPV
D6e2BKV6MpiIwMOMJl9oI6b46zz93lIQVweIC2iBmOTYUsoU18/B/6DgKgLxGEFH
9SBYQlD+677nfA43/9k7lsAWD/P32ozyEnoMI7aqo3LfNSIW/mGxU/Oio+7adqxL
Y7QcYfbjIWagvnR4ctJpBctoKrVA0SuFMEmF0rYjSZ4pKiV+n/EPDveLuQBIHpy3
HD/MlfAJw8nwe/AoYhGcBtq4uTYAN63qh4IRtHa3ohTAZTxq+hrNibzWFQF/tAgR
I5GfASJgF6LlJEaFhyiXyoFLe7oNdoELIg9T3M21Zcq5+LT/gtez6iJ+KvXPlDMP
RH01AXJ5UNUBF7xOvD6tfSekeqmMBdxM9FKWBJ80K7ay/fY0QUSRxYmrrZGAt6Q+
P6RiB0X067+djLLCEnDTG3DzUhDqaV3njnaquBQHkd4epoQUfzJqSF9g57HrLnfa
phfrmCG/uyijqURQpmytqNVqGJjMy1uNXvlctmWaoXDssCY+zMqMheY3ZhsU8/dl
nKHtTJDZGrVZB8hGDCoPp+Bku59UVsJ4En8NFwCPVQZYDof2XkI8cMVF6e0j/xvx
5WPm+L9pzIZN+PuQ2+DFpBrOVnjsxwBAXLCZiNPhNafisIqQ6oyayhU3X3Y5kfb0
dCIsCabOyH+tXsYwcAfolAJ5V1yM8Q68SaJiURKje47lXdK2uGffc5lgbeKT990u
5XlruJFFw0rGwNSb6969gh7qmXOfNQAoWMr3GkmVJpTxzQduuFfsn7/XEx73Sbb5
hKDJCgv7e9h6AdA5CukmBrd/i8oUQcoaV7Slrl3QxXqLjVOJi09+YZcbJYBl1Og2
0gGcYKlSowKY2vyuPkOYpEpRKwqUyNbSm1fw11FjlqXrkMT5tvDWNlDg4JdcEzb/
3RvkrfCHSs4aG0BwTqrQqTB0h+w+sffcJMZ5WAhTNfehvSRMhIq/NvstYZOaUYYI
KhK8PzWphSjAGDGdJY15VldXcx5pa6Lq5YVtoWcVOkd8eoMNHnH3YqFyNXS4Hyim
RBXGmneDmXfkftg2+GBfDvFtE8dEaAQRhWEVAeHRC08zcZyqi1n9YB5pM6K/maRu
3F97mxC5txKWOTfwwjgYs5ENmVS2hA2GAF/TdlfPm6Zi7b6z2nQW25zfngiLT20D
YZ+Hq6yFp0sQ5XTLUCuSS02hho3P81tFgrGIH/JExwVO4BeFInm0ZBIrU4ST+Qnn
EgEUiANXB3HGC0I+VpEoSCWpl04OtC3DhC0GHqo5lea+UJIQ+WqwfRLxPb8qlkd0
eKej52jDzT3rOXIyUsSgJEd1N21ioqtSFsjOFrx/uUwDqn4j8Dw7WykpVkeiLGY5
ikHSP9xVb16qQ7VyHk6guyo/PynWAiz3SJbbM5lb4OXRBqxEP9FT7k4kz+vOvQbE
QRzSH2q7OCFIELm2gTzfcw9J/eY34J7xB4INk0Ygd49Tv0ZWFxQN4OEccKd8kQ4/
8zgdOPwPeTRizLVY/r7C528AdVT5uzq+sgit7B3hzwNC6DGAPLwRcmYIgAO3tDz9
WxQDsR3R79yEsDFaXKQbpyO/1HjQKm6kurPqWp9VBmvcI3L/q2m8NWyRiSKTvgrD
KY9vSH8NZFL97JNte3+gfrXedYvJPnrljEGf5j84RdXfXIHyK7z4JzLfUJq4qzLb
UWwiOQWvCU9IgEkDDDAOQcxg+klrkSqOJSNpwKrqwT/G5fH2lQEWqkIPyPm8+s86
3fKgZGgJXvNZnBb3qUX8SzuPfS+FQxWQVvCgCmRRdFUsjla2JMCikZ6SYcn1tAF5
AlIGv2pTSj40svgoStodqoRN4vUQwE/uCwLN4fsXDMu/srwBg0IC1AO1hAfq9Gr1
MC4eXpiOAZ1IB+GHor4fF3DXXav7JtyuwP8TMkcKsf3YqedbWXpCRcB233/QUIQw
Sd7vGhjySwajTPMyjLlhn1UTL63ZUqNXl11dSM3SQgX6TID1KQpKyCn2g5hOqH4k
ZSgqZCBKEIb7nMixhmsTARG08P2gkrv+fnL1onT2sTwXtWPHSahyVvMv5rtRom8p
5TZHCvG70PmCjRukfYXQxkqtEWc91njlGGITEZke5CLSr1EZCJcoPAXatAnAXjji
dPY2lDF3Ujq4cC/xWHdY9yCI8pc8XgCLqgGMeypeCuH0fkt6nk8EY/Nvme8xGSfE
dq2Y1dwFU6pEScZ6ylr1ntGdKHSxheOY6CvGgclROkfHSQHPTspFfUgLay9Oq1M5
6CY5LoxgfRO4CffpLCxgz2DeTvjNIP2Vtiofn/Nj3jnlgUD5kcGIg5SmFcPvuZpZ
pbIolKnZewR1eIiQQSXK37vWTD2MZfDFprUZU8HLcqeJywRmaqJP5RM0a07DJILk
SwSuP1IHTXWDampCq/a5k3drnQZ82LAtoJ8eCSJjBAgOOAOmjVCrpiUtVR1Gl54F
ehrc7B77pGO9OKjSmCIeRQhNYF6CwWk55FgdYuM93KP2TnU3heVAta2opN6oRybV
9lR3Uj5c59S5SiPykiHiJjCi6GCgLH7JGguJ8WEufJFssCiqQqVkfUiDncsfOg6a
UkRSYh9VZm6VuHsu1Zbk0uz1qUeuo94bPmMR4u3G/R9Ar8NDV5QVXqdDA3ceySCs
TyAVsE2ED8G8Y73ruTCZd+4JEcZ5ExKrm/WVrm2SIJkgffscl0PtR7eHPQ5+kq6E
YvJUJ3dWPAZ5iElJ9pZFi5Uqj+nMSW9eU0Q7GQnztyLtv7Mo9UM/aYGvGO/Zn5j1
L7sAv/BZiHTIkRfuD6+bJX+5qQrrY693YyR4PmayV9dKhqnQH6P0n5Hw0mAGe4aq
rxRHvYD6KBdRTxj8t1dDLgOxn9twCDXoXqPPZcqVKg2MLmk3+QQEohyYsvPkqslo
VoDO7b9ySwA5zSAJrfSD8+K8r7saxGHgTJBlemxM5OZfvbq5I6W4OijRzNfu23Ov
tupI5xHtMfoEkcoxGwuaBa14toBytcdi8j2Eab8y8FR70LtTka4UVUB/E5CXlWhd
rdG78xzzYwloMcmgRiYJ0zTInn1XPbgboo6Okybh8OhC2NX6wpINqPzf4vKyIriE
oQN0qYOFjQ7GQLGLYkB9hFKe6iH8EBvPvryYRkpabiwE0IZyrlGPZATRQb/Fj3Sp
0CougLa84+UEYqxHPXTZKOJI84k2sEzmcQbJMTqHi5axsN8TNteMTYt7PT9I1Kvf
Z01r+Ir8alW8lWiEOi+q4qzR49uFSWJwIykEi0MhEK1z6nMVUZE8NtMj1t0Rn6U1
p6qiQSS7htqIHwkVPxMBYFGGwSyuPp94Xp0X8LA/K65SxOqV2FdW2zuhIfuyi/Gx
sV4zTlEllnY4Js2Xa5H1v0zEYzAztVXhlH2ZdxmDaEM+r/FxMyKd7F1cOiubm7zn
L2IrcdihCzSKou+SNYri0FBw7vPWKhKBLfQ3r4d+2Rqa9jPA2CBLBNnvwCoeBiso
kGV2xocHlLcsW5oJEnmLgKD+wDvqa7zw2oxbZYkx6UG8IqFjR6/wNfg5/YQukhyY
ZkXZtpR7SjD3PAZ0huZA7C2hDRIUplyhs9VHEmfdvk3tDEPcZVThlKnj9nLQiKn1
RiiBgaP7o1X8WouMRdkEROSFc1VXnBotmizsDfdQSQpwzU9xgQf7Mnfj/3WlgIJE
QU2MQER6yP4O5Bu7DLUYFd5Qexh8yYmv39TC72BgbQA+x6+5Zx6LVyo1mGISrQw9
RAsulUhpDL1ZSrENeUqHGZQivVBm7t5/USgezDeQaWM/Ta3WC7WY7z4KD6j4s9ip
VgBZFXbt6CuY5JB8ZcR5cWb1DdrtJtRIUMmRYpfmXwA00tkZhE0lUftytNS4gl2I
+xTHtigYWNJau9mA8nrNcFEEu51fmPAqPVQ5nn31UQOL43xNCEqXiFpo5ONOBARf
i6JZVRtZ0fuEHvtuqtQYe73T+EPp6S0/K9B5UHP+dqLjym8j9nv3goiBVf6xEu9l
Y30qvve0qt1YwKcOpOK5WdLDGnVv/qGKjywIjKRVa0J0q+H33BCsZh2IbfgydnQX
4U7L47UP3xXSW+UEDESinM1JslW4GHma8irzHuA0Ve5iL6VVAJzomOoEbveQfAfu
Yi8I4B/Ahasf2pMxfwIBL0NKEwgDuS5+6YVgM3Km2jlHLMU5Aj3SKhCFBw+jIwGO
zgzi1njmxEdyzTfFtxn2+OxTy0hw2MQf76IY6OcQXF8KQWBHdUUzUzleshuBiJnK
l+kEFK9kRoScgwRrVH0pSpg+Baa/R3b+sUHD/Qt2TrB1Q6rAw7bbeA1JEHb5Dzly
bDpXtwLHINDGoR5603VH8wgHoXBXIBIx48uBUdiN15mcVo3qcYc8UGEf/8BZEY+I
YoyrA8Fa1GCt6KgwQhiANTL24u82+dvIUf+oIC1Jv8/rgjNqyNMQs+OZCVCuiThz
WdnApUgRcAUAf5i4o7PYVhWpte6X0K1UP2iXGb4XRL3VaDseabP59zQiD27A64bF
VliFMG6s5H6wK9AgB6ZuLGXHhWJM5d4b7EHWuKa+uw6wy7HToc9pnJl0QNMd2yFP
o4h8C/2IlKKq4tgy249li8NWeAgfQXbYi2DqAORYs5P0t8qejp4Nzl46WTqNroYF
Gyxjw7ey07fOgSJHjk3rpRjQol6i91M17csqNIM7wRU0ofmoDiEkDRd9YgwOV3NR
9E9DprMIbkdYDJ0IGz+YyV9fVst//Wrs0B2O/KPi+9bFu/KTx0oGNNB2ImixPKra
+pMUIRrktyZk1MjAC4mqAOR1faNea/wb2GtafNEJUhIzr4MOwwFhaoq9hlT8gtH8
0RAwUlnVSUXBPNuhI/GJZ77VtY8odpecopo1xYXejtyucOb1DYBARSqGSZh21yQC
WWqpij6SnbInPelgmu5c+p50MK2auhW8QLiiCIwS8eN72Q8gsAtx6dOoRs+gAMVH
SjSGI/sz4/qO45cUGBpiA+j5hNIxmf+riyYHvhQhOtiUnUXbWsDw3xkXN5CILSTY
nPpD2FY8D/VJUnLcI5vHtW8JZ1Ya6sFgvr5T5ISX6Ar9iDzR9Q2QBi6qSWIyx9Q/
ZKYjjzQku8/paicn2uHX7PSAGnz2H/9nl0W1SKX407LnxYtHSl2O78hspvfF3SyC
btnqaQbDBt7+2bYLEHe66aznLSqGJpOzWOEB/AxrVAoqu3c+vFG0inQDm9YSeC/H
gRJcTJoaDA+wSsogoG7dX4HsLPGckTPHYrprBuACWVzB9RSKBcJXlRbZSPO/lEsN
AADsI573jmIYUhGLswxCBA3NwrSAvkxjvXHLhpqbUD4Z6WhimawmJd56LISsOf/Q
8PORCpGRoe50g3Tryjq/FsLFErajsE2emk8sEFUgH5azdVSz588uysLhhxFE/f0x
neGaQfZ864csSVCmIZOcABNwOtFJ6DDrC9RMLdVLnORLC5JMuOppobvvsCEcUb/x
bg9DWrGaKE5icYUbzZXQ+wblPQvbO7h0Uxqnwhw9AdG619GRWjSQzTt7wSJTsdi4
sfhO6buSm0BHCtYvNCLVL4XhhWKPMIy9JJfGG1KmTLCiJMXOuWKLKleC+8yHtHHK
mjKl2F4nHqEKnQpTMvtsJLb9z5nwKb2NqsIcEJFiquUBeWqetlctqczTnzLo8uGj
66pTW4nwBHbJok1cXPL36LM+LSisXZ9y1VMe7pAZKeIZh41Uw9aLs+LRxrmTyMO1
0t9W+BVxvEIxRWQy8jIgelFV4oNq/W0oeHP/0mgCQ1OcVRL/slGugz0vke+wHOSZ
67l64V7hB1JG4v8SzhJQ8FFx/+yAe0EZvv4LDclI6o3QAMsHmRkRt8i8n7cK0NZD
MPATx/HkFA7cv3H2a3kSvGgx/mPgvHCgSH1TDJaPRCb4TdfJFvT86iNAhMEUkNyp
OYu4Th5qdUVMirPNnE7fFvv0v5RxKeCO2uz3yc/YPsDkE4W49bxDDS1BJsC6MW3e
BenWQdbAqI1S66iLshDi4P9o9WxrHwdj8CHHePTkugCVQAFGHl1XMhPZP4wW0aLJ
Jp97jpahPDNmb6XQ811QzqX7nwGKqV/F+rSaSZ5njb9mZ40sYyxREEQKawUQ/MI+
iwx1QmNr9ZVzZgZHxjaZm07KthSrIerjZVtIWtYgeKUMomRNMV15Rs69jlDYkjd/
H+qAm5yVmYTIiJClS1prWMtRDxNpm0Mi0yu5YR2/XbMV38t0SJvZl4Z9R7lVRR0c
uQ1MGkhGNyY32i7tu7IHvoVt2D+wYtUQ5hyc918J4mvQR/dzi5MqMtggNtXaoqNl
8F1gIgSFM+YzUL2Ho0ayGDwSqXxUC31TwE00xFA7vTWmc6LIWHPtfZf2qzdavw6e
bJbYeMPFCyig3U0IJ05Yz5bKijexJIWg4xYWYT6Vq5V1AJps+B+4sJf26HMT97tL
ddMW+i08tK/3+2UuNP2LpBP3JSxM88lHYzJgj0gFJPmK8r6rlhFiLJcfCWp7pjyP
0gg1cMZkVjlKPc2M6lRFkcwW3xmkU+vtpY8xj59g3xdC0HO0Nj9yPgAD8+F6r+Ml
62t/zPu2g8ykleEkJ1tfSVMudi6ujFlPKhViqc5X2IlPeO9XOIBf1ZLrNHkmb2p3
yzsUUjRNE8JAw/ODflG3BQXicsWPkl+6KZoiHd9JXyLQOO8iY8Hc7R8SHwo8/bu/
ZnoGRQHV5T5kisxp13zEb+Sq4TqC6cu9zRLFgd1SzoNBJP1+Q6J7yGxYbRoCyEgV
dCncJHTKwVcfWDdABD6AyALDO+ygoqMvvltk1MnRSiWE2gjbcn7u3cXzJKRezxSl
K4CM22uRmh7psHLONludY+fsoIVCT8njRkCUqw5cKdhgpYDMW4nlCJ0fcozdt4Im
wecrhRJJR01JYfRQT7dCo+1IBsSZ9/sVfvfD4Op4OiZGKkrCoe90v7zzCuqPiCyR
4ZZcui6JKV75Z66t2Lz+Fo6IIkYf5QfC/UVRDxkcYJ+Sky1Y9iehrdKW7LSCWQri
e4AUhlSCUXP4gbVMPRVAIiJ6YZQRJ/VTZCOhg0/vf8lr+Qlj9FC80dJugNEdZrul
FgiTFBSIdlXLHCnt7tAg352fGqu+T0TH19QLhu9cwni4P3e/60xVZmj8iEFL0pR9
NSnepfDYAMTF1OIg8FzZ0VsnYEAx7ZeD1H99D6XQZ1F9Ud8BuDcK6Qjncdbo8m85
IGOpK4EBVBhdai3kJOfte3aG4Hxowo4aLyM3d52OValGl7iu9cL4V5LD9qXv7n+0
NvW/HZJNsZompBN5rmYVmtQvun8Fw8BQG/NSBae8Pz3b5GgqTOHLdgT3jDuio5E0
J3OFEfFx9Kmf9QOEa7TSYgTKpcy3hnbGnHWsMLPembaScrv7O2maA0vFK6syVX8/
AR5nYN+zrQsToumnMounjxdUtTpxshOkHDJO0CjHiGAqXh/SPs1eEqQ2fhEXtpMv
K/FJ7kXJabRyRhtzgaqLoM3AaS+QOVsQdQC4vGIMPAYIjsaqPHMdxdxRhLP44v+q
kbjU9e1rrAHPRaTk3pHcXj3xLy0EE7vT+YH4xqfoecG2Kh96tNUpt5FRz7ghDdDk
l1qQqSARo+Ngg13/8czBxdvTrwXSLuttTNJRPlobZed2wjelQoCbB7YJi+kX6eqP
0pBg9g+Xey8aLxxMCdq84ZAbwBRpvPxeEYb4iCQ0LxnKdmUVgZQ+R31oEpxdMRSr
/xyY7VzGd1vhnRp+u9YhlJVD3f6yKwOtPqpDnRtBGm51p+wRsGUbXHUNIdZCzS5r
20WecH2keC2dwLm/G6CmeEpl16MzEt2jmnJxiifoc/ADAr87MC82jUiORIkVNz3K
RU7q/L/rXBY8L+5SI8jc6nzSI8K9oszurary8Dcjgx/ZZuXC4r3v2Py9VjJ88Jck
C3Qwj6ifQKyeWaacoU4698uBxEE6M5SZqcA3Lc8SfLSDb9dEjPgiIlkbX1+t35rn
RMRjFh6M5DR+bQHjFck2UqK0ojUcnzKIzVKmeK8ozo4nVLfKHLijtBc3sYLYqoUd
k4XeEqnPD1UHWGFgplE2r5gWRv77zANOWwdZLO0UC7tsmKPhUz9O//6sj/yeP21K
5zs57skVVhRxkfntWogvuKzWJQxPXOfPFjTPYOMdP/eBaQi1uwA/F7Ck0tTfh7sh
+6D3xeh4pDvfqgkziI0AqfhpO2kdBKBTaJpVyzdjFi/ioi+UOXwdbBAuiLAI5B7L
A96t6WeoeR73CRtyF41fuxzYAROOVRv3NIslQhu0404wNQzJEWx/GqaSFJ/WKTGo
lyvZpetl/ptxEmIjrcVCLFbok5GC4mXqQTEL0i8u+Rd5KtUHxIqOcWq9Er63REGm
jhdvfkuCRTxAwLaplyiu7xgJEyVVhlttNHz0wz9fgiH0oDIujWGid+NnoIlEcLSP
GU4NvO6ag6hzmmcdXxLlrcoeq3ONmhZiWEiHshFoEiWXYVuvTa3CCX9rM4gYG3Fi
/o9BlM58uxsmtSMuoNGIiy5r3BZPnSBclMhX4tOMiAoU52+GJQluP8l++E9hMl37
va1GKgXrH9LmwBBDQn0RXZt1rdxtL6DgjNxylsmJ9dMitVLEQROAmKQq1SXWTnPj
eud9pz6EdyXDP5WMmnLvRiybSAEOcEtzKKtbXTqazUmJsVvEaComqpSQYVrt43Fu
g49QLq5bxFijNQ/isuFJaPFGI0jToZ+RgGAllCVX4HVW33B6/JBYHKXlon0zPSau
W1saz1/JsSPkTe/nSygd98gJnRRKJZKQ/zeKy8CZLG3LcFPuj5Le9+9V0VupRhUc
EgdRp40MykooyCF9hI0/vEPU7Lphn2ZBhBBwp396zMXaY63P7cs+HX3PjUg+k5XZ
DVWg+9BgBGUbt3UE3egXBFgw7qhyVc2swqajHidjPt5UfJwsl9YQup0Wsk3AfSyD
ONMIjWjHDwUD9f4+LDdPB0IMJ3r2rgKeH5MGrg6eeBdI2W1lLCdnpljCwBcw0yI6
7s4VOWWf+tDnMgUVPVkT2WBl9cMrlrYYsLQqC9lJhyQrwEpoGGJnwB4uaHXYzQ6q
Bfgdd9y4hMBayyDPw58Gg8LGRpGY0nkoknZCEzDjP8O3r0B0TbwRC+Hq08BkSnw9
eu7AgA1vqKTP9m7bt2So6yFETdYlQr8ZAn+iKVhKH4703imzTt/lBY0ciWo0a0j/
xHYxmPYE1HAQSeJx7HNAvgLIuMiPjr2NjYqn2gNkHHd+EoQUxyalIpvhQaCSXJwk
AHMONLKqcteSLiQkuYshIgafLBFQV4Xrz9AirwRNOR+BRyvNZ9pZj7YP3iHyuzlj
sBvCU7b8R6Bh3oYHNPWkkMmb7b/oQGx2VVOvmidQ//j9psemrQRLkDiQdM86SR3/
faJV1gCVULEiCf+1xBIj3l6eueTd2IlC0L7A93uGNsrcQboBJ/QNZMLVqFkIPBUf
7dqngA5igBPiRjSULdJzN3nDp2gSAfgeiso76a+MIiZhHkC7bM7gcSDmbNIpwijy
4qGjgtD6uryM7tjkSxpx7CWnkCGDH1EDCRoyZk9ABaL94naVeODZuE0QT0jOO9b2
4Rgt4JxxKNkM683XoPOMbucUevKRn4EhNhZZjHrPGFSej+/uMUJ/fxxCO0lTVoBu
CLF/VG5dLKpMFkyHfYtDVaLMTe0JqrvQw6jU74oqF4W2Vb3iY3jn1k+IZ+eGMZwi
QyYD1TeqB92+AnLsmKJNAylA4KtwoGdoJHhQk096bFYRhZnJkYV0pybPWol3qt7o
X5FjnH6QfUIIUP6tKBIa6J3KIwq//yAIKw0rkgzabmLtO2fYr17T1sIglO7tkQFm
03H/xK1Kw30YvW2+VRcCXPiUXeFOCJkhkcNtucuG0V79be6rWkWS3aJLsTo4vs/+
P5biTolkAYu92krjspzjHogWuXN2pFf0IxIj7jEUzpOz9L9n7hNNTA4K/+2qPxN+
g39nO5UshMd/Ph3tBxu2BNxDeLTgV/967Xu2zIyS2MzyVYQKkznmbs0dZlIFLheP
t137NJVOpxHNl2f9VgTx8XKZ95wI247SyMRKYT0Xv5Xus37biCsrkUD223QNbTqC
2JOaNLs5eb1cdvEhnXnO1KPDdYHxZBdiyxP1tQvS1L7zxlIe/jvc7AArbrd997vr
d2xCe5Hu5flXxxO1WteIO9Uqk6qulUMjNMEaOq6sEv5M9wA8ATVNzRejqs6Hl7FY
kA1fIrL7hwWF1q/QaX4qJgIsWPqwB09VKkdgPyE81rr8TzrMu7RDJDSQvzWv0t6Z
vQmS8kkznT4PL0lTqTnONnCmz0P7e/+MSg7hIJF3zDdPfNOqKIcCt9dbnNnr8ptI
mSKDmlY4lGMbKuEmdmtzXdP3/sucN6XdtsXNtuUrxXpGJxReS94aMeinUE0T468M
FZwFP2AE6RQa6Zv6MdkxHdqjAluRILarEEd8Sot5Mr9zmCp8BrO86pYwLGUtonfl
5VRCTmPvDjDrpQtO4IJ+Gq75jPqNp/RGWrs6o+OSYuITLMRDYciOg56+mVYzvuED
Lj+PQ7Z3/4v+cf9tNzkRIWR54bP4Dp2/JPvHq83G3GB11DX6FEhf1hgmxWXJdI0r
mXywgC93JfChkdx1jvX56fznc07hvsvAexNplIQihx/WQUBLIyNW62YCxCagctKN
35fJ9ogrSq8CH75z9hAIayyqJMAK4Dj1URSO3MS2HXHSs5BirzAIZ0cN5gptGNbq
iowr1oihjZAq/D0qvKFnTuvDrpkICCIFEhgWNAaJhqii9RUhEP8oqXDwFlFzGw+H
037/H8+baMYh1YYuqJawbl/ay/abbEQvhY4wADtRmZHGSmcOA3aMyxBODmFdiFDg
SPjTSYnqQmonzA6qPkY58Wgpq5PnJnYLsimF/Ii9VdVSomci+9HLLj7LT9hyCRfN
shcdv6zVPrzMMGR/ZrMAeQUPxdGYTrIz+uFOmk88T3CZbkTQ3UPaiIcKLdq3ZmJD
/qL1BIv7lct9aWE7FGaNa9Fo94yYVIhu2biiGV+9Ec/RBA9akzwALBfVfPZsfp3r
xSd4xWsh3xcFx8rhe8SulObflecDsfVj+TRZPgqJbyM1WXi/QL88yYTYPdOngfMO
RlZG9MqzUcqxTjnpWj9lbYLNPOxtI+1v9SNlmoAjZisHTu7Nan/DSYDMi3nAnp0w
ICoYz7ntGYPCZUxGLBX2UIVBqmyFKeUtsTYYY6DZt9flLRQjc8e1de/geOKlwUq5
CkXt/9Z67/0WhAMcVBFqxh7V2roY1tZAMQnmuHDiWrQc81UI0ENzSxc8bzezntNd
JmuUNpmwCKkIwUR/K/1UEGjgTo3rjNGU8UfkB+Cjg+dbZyfYiv6QMhD41F8TjldF
6BuSnOLtAV42+T8OTVNH0hPA0UwpsqbJAoGR3qyOAtEl9t6DACqiBpSc4fTVamUI
C/VkhcRCxFt5w4+3FfohfmvtYRPN4GShPEh+TeF8p6Jp0KUMqQV0yQYiCsL5eO2w
JqyOgCtffT8AOtSQ8jtbMBbxOXLdBmuMXvx1VGexKAB2xoP26FNM7nDbU7+Hrq/7
JBf4AhoMA/TdzEHN8ec+s7kHiTDoST8+QbQSwoZ/ATics0EBaK0UVyxkgnIlk8cV
zz9GJLkqKL6/JuXEA1JdOadSfR1s4vimcrspd4/HV4gyw6Z/glw7YpRaEj3iMu0v
WHdR+XQ7LOPrwQtFzjp0pLeCVWezkBvpp4spKbAV1hgbSWt8lapsmrBHAS8aB6Zg
/hCTU26/ia6O8Ij/PAcqP2B3JA0hYTNtpRK5eKV3hC2msC+Eo05cVVR+siupYrlu
yZls60lUwQ1iVHHLf0XaaWo8EPIb0ubt1KV+ne7B2lgsnX7WVzJj1+X/EAxKjpht
DlyOEQSvU5IV0JPX9icHjskJJ59V2u4gX3c6e7ENDW8l0Z8eCukYUQMcuSV1uEmf
uN8ugFQTRx9doUaDiEY5wz5nLARUs5BT1Uvx+cD6BaCpAOtFhyaVmyyudhw8zwCo
8hlFx/novrbjxpExXvr7lk5OqpGVLwfGCnYR9ooG9zJxjemGDRbnca8mepcuURfV
XCJzlJyfD/rB/bZFE9qe0nhG8bt4cc5fNvIvN6oOyuNNrF9PHafV9ForSDmcIWgB
5w+c2PW1lzEg0CdWHY+A2qb9tFWGYBIqxWhUrAg0Pi/1jmWKtzFddL3ThpcAwBYu
qOhTKgl0KJ0k18lZgQ/H7LP4TrJkiIkUqi6EbnQLbKRcH3IiSIlsLYcStL1JQH+M
B2cIC+q80bDat3NV7iMsoO4P/ZC5m3mA7p+iPh4ZiKZpiAbV4In1VJOPbZhN/mHJ
+TU5Cypr1Xslpis6ubhybMoqCOeukZaxdlLqvLoI83GRttBU0Wx9/wYX7/0wjFmi
ZzbEFuuuRqAR2SFXWB+1BzAjtvlZxZgG/3VFH3pqlp93LDEYW1p2GkBT8+o+dzSP
IAHs3h7cjxlMN5DZdVBVDX7iQ8kkO5X11pcJMzvBAOCcdqyvXCqU82X+Ny4iWlyP
QWZ7JQMYOdCcE6FwXHEVKzlHx/wB6ION5NdY4v7Z2Pni47uAXA/lbFQLQn0oAv8x
GBvhxtkSnwTPWbTdfooeVjfmha4Xjie0YrE5061FZeX6Qm4QPfUxLbUKiC1eIlAy
/+Y3hJ7gjNlagJevE15MwcgRGb91IwOoncoxCrOQiSyDIf/1kjo4sT2RXmiG9Vzj
3r6ml9i0Dkr+AfKsUsYYYjssoTVu5nnlqSeaiNv2MaxMrCidSjlPwpQ4H+0tyM3T
mvTk4FYKmRpyunmE4u02hK0bspTJ3oo8CvGjN2BV929lb041dMEOSzwpY2Pa5mMp
ARJEtYThFovAcBM6NeXb/5t8JddulBLj28H3wvWZ3glcJ/McYgaYob0q+NbbzBTD
/n2fv/vsh+IYE9Ha1q7dhaDH2K3ZwBpDCp4VwmSkE0j9mKgv/NQAE+EtdpcxVXg3
DoU0pOz1UX3kWIMRruNFSnPY7KZmm7JIYY2h70kqeZFRLTiJzIa8Vv3Ad/ScB2Bz
y4aPbeHh2K/wqtdO3ZknXDR9ivKUuVrkPerCEnOqCpO2+wFhhiTUf1N06GP4Qb2w
K9z03qGQGXJiGBWPHZWMOtQ1ypL8Oj+6kHD7wbVfa66ngJUt/noWrMlEQIgohz6J
FycCUGCVBVcvfZtDA7S9Pn2onVEtEa/6wPW7DAK8wb1OF28KpkHjZUzGQW3yoJIl
dXy0W7KwpQodDbBS84mArhqoRYnrmuGoL5GWymRWHJRwTxDK9n3lfAbnpROaiw/R
WSmQgb40i5ncD0fc2mxVNMVM79oS73XPu7oGcrh/S9+9rCfOxMuvC80cUyUOZT3T
QWq/4CuMWhvGMZjLj3S66X/PPiM7ZBRbh2EMD6qFaU46AxqQ9k5hdKoCG+P4ByDf
9HdMmc9GVwOD1z7NpFP/OTbze4B++nf56UWESVgUMdNsEUwJCvuwr3/d9knbLKZh
6Y9ljUggm9bsGHT96GUl74mWRjkFOR1pSr14yN4DGe9wgd+dghvnZssuXiNY1+Bi
OTt4UVp3lFEkhS5yhzDMvCMt39cGNiwnlaKFOPxHIVCuftVV2MLHXsVk17ayA5LY
fpKaWlk9K3dZ0YaTVJ5bIVrd4/bpIytfYCEUgOcCQQk+jTxTb+Bqllpw7OInj0hc
303gnDeDApWv+1QDukDq2g+iZmydln6LskjQ+bFl6ZfK574afgylLshfzKdrkKZc
jfBchYcp6T0NVIJFSpkKsKqsXe1bqq1HGCvcqzKV4APalEfPqeO7GHFDYqrto+h+
sf6GbDJej+it/jwjGO1kbWxc/o6m893c0T6byjEjCDHXeACAstAv8grF3dZQbBXf
33Kg5ioszDThr4PxAUWL6xzq+z2ONCBsEw3FnKf0z3lei498R4tZSymE8VojA5b6
+e/Lffc1UAIf2EZiGBe8OglEKWmiTQ7dI7ffw2lOBhXewQ8YRRxqjgCDRZBmOVTm
g1iAr+K/MEa1P33n4/zHep5DVrK4G8KP3+GxDkxbpzQ55VuflOg/8r233OMB4yDq
cLI6mPkcOYRF4399BFfInUHl0DeKNy8F4Z7t16ERDL+tMobtPkmombmc+fWKmDCP
RPywSBMnwf8c2ncRx9vpCkcN0FDmD0wv3pn+IHbkKhSfHodRcHPq2NIE9ROWnzKC
ck+j0SMUvFDml+NYy15IEYJe5vJAJjzc/kBBEdN/P/IhXQ2h6QA9biBBZvY/T0Bt
Z+jlJXOWMtvAksGKhDnVtlJOkb6YCro9gz/420GR6izlMh04fEw5TMTLr/EyceEO
oAPpuxmqZtIJ5Z5qNG8jiUDoal3KwqX5b+THn8HrXCh35Irmo0qvEeg9WV6QQg0i
PUn4c23nyaamPRiZP0JgAQQeR3KrmrRx0PImdD741CSyjlm5ANOM34DEB1gFXHO7
dukFCGvnN77aB5xqXcUe3zCOI6xS0rVvjxM4nNyCWqbPm7JygGWOX7GpnW2EHaT9
NT1VOGLbHBSC4iAXODhdVLtq+hlXz3+VoWxYRrJ3vv/bAeZL3EyIS56DuL3BU3vN
55FFwpndAuV+tw2I9VVnPfz2LKDKNP/wu/oU3N6LFPRxqiQumLBsIrWeMOXDZYfN
ZbtY67l8z0ArfNSgulh/SunizgEK6fHoi+yBbRpQFzpEAky/mJoL0uO1tYjBwrnV
hnQ64axbiHobMIBJLGOT6NsepkOUJbY1foyxnxmFqfX2N60wD4V3ueKIzSTpdidd
G+sWuIv2vEF6AR5HxJ6FzynvO5Pf3cOY2GLoRn/SbZ7OXeUukpUlVzPBwCkhkEnt
NsV8nI26Lz6qAtEg7ws3ZLoeZtoutO5fVtGIEVTGMF7VaLGDa8ynqWfEqT+lqy7L
jvlu/ehbcztXDvhyhVB3NosuikwGuYdIk91fAc5tzgIVSlOEJzqVUggN4MxpjKMo
mbfGrlY9hQ53H9XQESNhodPveoWBI9ct1/xpXaZq2XDS/GeXkvPzvV2ycNa1+V7o
c/77PgFw+f5DdAcrkiChLw8/gg0TeJQ0SlgHh5bUtAeFj7NUaBBkrX92WtST4Pn3
tDSkzkL2aV2JcgKnmzVoY+Hr8ho9AVTKNXrm6Emqt2s1zeVp4OPWwzFKuCzrt40b
cE6N7+6QLo+SUAFuj5/0Cd0GTJ+CpqBrJiI6ycRholkGpW0wEB/zUHqBCadPQ79t
wf9waZUDfHQrxHAIIms+lIH44AgxFtBcojyyx2YvBzVjAgSo7MXdoGEummTTX5zs
2zBOBLM8YsAXm42X4FKksPA3rk0vxyWbcU2Dal/gOwgnL83YjI6YX3ROqDVwARMI
gjRHMkAjIo5/jwK0lMIjd5O028FXwuDgo0zvwrqOFJWpT7dhuUmALhbg4qmWNoDb
+1jdf2ihFUpSy6V0c4uaxFvUGiDn+vPUsnSiK6rg/ErvEQ4oiPs5FDgIwK01vmeE
Ruv6tELK+YHYybJYnfDcBBelU5kLSfSzxCI4Ch+Mu/1I01JYWfZlvmDtUj21neiM
FGAv5CycnTi990ee2o1ndLQEnrZillhzwPQNPVq/hEPA9hnQa8cEJFJoaZBe26Nf
1HGQhDbkp4RHicAxbmgSaQ9qImjQjvSWxXwXef59qxesveQ2BMxQzieTItlKmkSH
X1SewWEG4X6tJKjfBLl25dTaKHmvpmxRgywCX3quIWxhfkS1U7YjMCWF+4tn7s5T
q52X/7KN9E4ccSq0+VBK+pRkiHZr3BiaePflkbs0FLl1yCf2NcuT/Ty8sywg7gK+
ghyVqS/rY5bPMWQI61e2QVZhuz9NmxqiQT7orWd1GDi/Lfdcpf8ZU6Jx9eQIwzHx
shbDuFGVwvwFmjbWoWmQ9bwOKSrv3Vo+Y11apkSbJZxw+zrs5D53Ma56xKL7RBdV
7pjPcS8TqRdrnON4YXwXU5eRwF1CHucOpIxAlT+hluwIsvpokn25ABU04wPaxyAI
/LXNfZpLuJ4ioVlAZMaGebZcw4ERuf/s7DqJszATAXmbD/v5jytIPoR+BNoj8xJ5
b9oEPgY9bC+8ZLxxtWekE7l2X/0Iap+v19oHUBwWUKtwKEDEdykeZvlDT+krVoeN
eDKi8buJzRL6TDVoqxd0c/hwZcWgiSMs4e8/gSwU7C0n8gIMzYE3q17ED92zrjuI
ROlnkjlnFHeHefJROVcASasrRjoBPizeO2XDOCHAOqtR7E17ZlfgXZ6wqPMH+y6n
8FbendyahKxHbQNQOpqUvj9guw6C6eOaRTEfnfaF6KNMESY+aTzkZoaIlx9O/nFL
3FnCXQkYI1MnZIgDTfNQ+HQIN3jp+RpeBQsOnOaU82tkYfG7zaJUgWiLi/cBW+11
APthu3IBlTeooN/xk1GGSwxuxuUQL+YwDh2lQqv+0AIBlq0FyJYYhMUpyIFjiMjJ
MrqJRCSMc7/rfFNIisT5aOp8PRqG649FzYJcjuQHBwGShGaY2LtVIwX6m5usprU3
XZKjWFuHFFOW5841jfjKeXrWrIlsdanfYWVHZKIiJ03c8xdMZS9J93voCreV8kSw
VMKEa+7QLNjX9WjYBeVBN0lW9oqz7QTvVPY5x5ZLETvYyITofvLSaSYT2KC+ziux
y78yS5h4af4VPxm7e7BqIZuXs5mhYZ5LvwvijBeL5hW59J5hRS/4EuB5g0bV6kXO
eZnrV6nuAcwauzsjvxK+maiz+EZW1/a15x7kyMaLb6wkjhNUDxR4j6EIOtMXIsP/
J9hFqHQu0YRHx0etPiohFn2WNI8Gjat1o3tONuDQITQdNA+3oJbKG0Iyd431KoTU
NprqFrjTrqOm+xjp9ZHhkBX2HsQEst2+54wSIN5P9+AeStCfrlciy+ZeZ3X2Hi8S
LaCagLs8uFVHXu/K2hm44HS7IxHHJtv+DjzjcoYHdgPeOJ5Mdp65T2ny6qRkDeS+
0A7kF5OJcTjm6S9srtlBrXKxS2PWWmm+uIVhz23ettbGtmhR7QyW1vp7PfQV4K3d
R3NKFFAjVQ6ux4HXWjOJ3WoJ7WnFVGWBufx3i0SLJ/K4j0tDCoIy5p+evETq9WHw
7g6Ar3wTj4eLWf1EPnMJwUY593kuXr2IDJ6WIsumfWOdsUgZYwCHl58ZwHxF8FHJ
9/q8mUgI02v1yTvcHHk2BZReg5xIM3Z7kNFRxzKMJPnRTEXFzypnHffIXJhLGq47
tRT/Pp7LllcWZzZSuQxekavohcJ5YqnYnTg0XNswQzsj+18+M7N30P9PQ+x3fIEW
Kxg3AQ+/UMcUFSpPXMSYhaLt5+82Dw0DZdkkhFFbPcjIzVk96TsEzggELKzozxQK
cPUgd8/F2AnFZZ6C/NI3ndSdwkevOzp4k5phCqehACsVG+jzASPdLmvkSZACQfRD
OjUBX+0DK3VCg3Zg4Lh45Y4BJVDi8QIkz4wUoIKvYHkBnpd4C5xcciBUVS6MVJml
C0NBuLYlkcbEuLWeKF9TgSTbwhxZoEnubsEAPVK2idm/XGn6rmuiB4CfBME7CMoO
UOGPLPgx5xxZbbDHqW1mbWLfSftVTWHVgsn8aozX75LqUsF0dykGkSYYemdNzduL
K1aSQahK9k8KpVK/T8trmpy5o7HKhi3ktnC/1KKollw5K7a6oU3hmjf8NFcoC+S4
HQ3C/Fs6tYd4Y+7ogjGFDUeiFykvfzSlegbnF9mscywJug8mChH76PBcCMM2t1l/
6edS6d0RMq43QwH2N5M4UfXqHCCmBfov2GKu6JqXmM2y7CuCVwOBU4cOXhFwNd0z
Mkmbx2qiOahmqGxejps+fUvVRaK+3s4spl5Pa4ifAtZ5CrLYgpgPLvRUKiRho8jm
GQKal6lWFhxVqyCCPBmrtAeOEKh6k+xIXvJMGXIBgWwTi38jIyvhsslMLOzrd+5P
dp3aJR2d5JNszmlGvNzz9w6LMD3RK1XQovPBba5Gsnixjhl00ajyI3gj3AkuwIL5
B2W0Er6MrJV6Pmm1xYdhu7KsH1OBXFk1hLg4Wze+KAJDQIfY+wlfzEEjDlAP2/hF
vexxRxIwqOdcmuPoPAS+1U21hcbOE1DpPkhhEBTZDrK7reXiVuMGUhrYXDQmIIkm
CcC8hBScdOFhyJVh6qykYmmDsHt5/i8QXkT/6ZMCgq+fHrESUta/dUEu3QE46hmf
ZwWKqc6fszVbiOg/kCMxgTK87y244/iQyFksRNKobA4NaP7BnU8jJpYAYlb1Nru6
IL0qbB6wE/94HP3QzSKsNs0wNVCJatvNX/GD4s2R4ZDJxQv1gicmCbwjlDFPvh0o
wnYd58tpdTuxiQCrIeNtp408nm1a7l/8F3k5GoxUGJ7xn912B2/sb+v+NNTjVfx7
lLps65cE34POGcUp1QXUUANhfy6+8hSVT4qfIEmowoQ+ExLoE1plZPeX6pwG6xJ+
D+7chCbu7T3uSknfIyclONckUPulWHmwK8H8Dgf94HLZyukeiQUev3oXti+AP2gx
CpL/vqAtTDSm2FdWEeUfJbtTepvDBy/GMPWA+IRnxyzuK3jk3ow+H/FkEuziwPwO
Z5avkBpEq4XR8lBp9UeZ/QAKJYOJnKJRBY4GqKsXGc9/NsFYI11SM39qHmwcXOcf
BKE7fo2QP+1/01+y40x20+v+YI7CYOI8Nl63P8WH82aQiDz2VE5FynDe3Z01Fhgz
HLPX8tpWVdlCmxMDV3/DwYC7XHuMn7kagPCkRQLsNOxS2vdNWX+Nh28qq9nLAygc
b/27m45qb5+GewmRoMHgsONocNH9Wn7HyGW4CBeV9QbyQ1YBpd1tUTPU6wHhgKIG
SiA0xEhgTF69NaERlb/5MM2FWsX8fv8tfKd8FaeQUPnHOKBoEO4qF0P2nv6MWn69
erSRWp1kd5bF7D/2qAbjJasYkWOq1wBa3B6QTxihdTPP4YbK0o14/GABZr/8WkS7
uX+iLPYBX/whzQD8ugiQvRGtjrI3qgiCi/+Y3gZpEt7b1YCLOtl3Nccm6IE/5UvX
GrrWYlyc1mcUmNVjvDmagUiGeGWxC8QzgPUgx0emWCBMx7YSuly94li+/93M9Qx8
/E+bFhDtLmwX6dy5pp+lwha4uIaw86YXG38Wiy6vsv5++HJsCRx0JjSS43j3xa4p
iyMeK3/JhrpGSuntutsWGVfP0K4EBj3Yd1IdO/0xXczCF0HmgtTQ0bFScs/V+nOl
7f55m9p6Nt3CPMMqC7wsIznsq+vdaLzk+10bxyZoFkxJuAiOAx6x1E6Du9Z+j/ig
VBWlpH5YYsFVywjuERjnvdVwOLCpqYqI251OAseJWgXrAI9uJckog9ZbiZwnW9iI
8xu1ubbJuYRfTaoJbp2ioDkcN99YUcdUxgzIsjFzYMQAG7c5x2Phr2IdRnclKh4G
/fGDZrMEACDkMPS0MT+euX+z5MSmcGqt8gsE38l8/jyyaUtVvT03uA0KnPiYQXlx
XmQb3NDyjd37BNMCVPSLa9LgTdfUEIsZ+Q9YedCQhMuH9l776Yi8tJcn1KB+v9/Z
hsZtsNm6pAmmei7p8qVYVg4brW1BaRttTeunpwknKPlsHOLp+lFRvZt0HVfHqNhd
hF4Z6lCZQX/VsYe0ZOO88TLsMD1XpHJPKkpDFSUEoDOFmA17HcQ2sMEfUz9JIKN+
HYNql1Sq6/UCekS0TVSMKptCiCSiqhbhtzy8nUQ5Sda2LvLysydOXMuM2CGrCpJS
NVv+8/KDBo2fzQPT9RfpcrFeeAnxavoUQnU7Ev413vzhNF72XtN/9xBfFk4kuyiN
ZWP0mqvfy2nT/Hr6umVdvpD8UeDzQ18jDws80XKD3wuJ83M5Hv1dZLOQKpYSyhCK
KJkcsbtz1tH9OkZideeDIw2utrfVzXxMmj1rsj0yhGFREX8Ldspg6IcPc9XPrCqE
omP5/PFOklQUQQJ5ASSg2eYIpCGELFqu0gRQP9WLCQvhzoTY0kJD21rvBGgF1UbX
AGyBe6KdoxVqVbSzXtegYoEgmW6TwaQi3AM2xXuaNi/yClfTeIkdcpbzTVvHwG8/
+KVa0c5wq+6sYT9g/4pZFLpXXVKxODIG54U0b9gm0nsQ0ZDLGgOD9m7rX4HhDWQb
qb16JV7ulS9OUYcmxayQjakCLBESQ3OY3952cSc+5itJHwjkkmSD3788WmgBT6mE
erl2jWTU9PqDhqosCnaph9vl6P7nPh1EWzX6j2YygppeiHjVDoK0lHumulM3dj8a
42xy0V3Twp9aqNxKt4WUtNfiLsgShHSVkqI/4h1pkLrajNuDnz1+xB/Zg+gMEWNr
D85Kb9trR486x3JT2z+tedLe4pvPZo9hQvFYwKOcPtS/G7qwAGNpoIZzMP0CcRbG
cTMYbqAxQUqoV0rayDwvyUXDQ6aqUEEOUi4SupnjE3GGmeqY6keX/3M7M33cnJzt
N3GE179LIPFLo0m6ODsu9yzO0YTv6NuaYULANTNX4nIAG9ql6l2JpORAhFTccasc
bN/gJH9c+tUkQq4o8S1BSgHSI+q1ogS7Qg0zIh3HPqXWADbd5PGdCqzju06g/ao1
FAEftXEHLlzTNv+cWWelkBLl/ZRW+Ju/+SM2B3dBoSAzFUEMhWMOUcUmwYRBshXq
+UIfTKqidVKgQMqvDBJ9t0OfAiO7rVOBWf3BCegSIk7x/GtvbTrZ+x+q8+5q4axV
Bd63uYy8sUIcYqUHLQkvStsGInB/SvYc8Oo3coasH70lZykkJJ9lL3RlyaUawgLB
maax2pq95LXPr7yta9Ak5fhMroc+JuiX/7aSawOe/tU/7SlnEGN4CERnurhUgfZH
IfikigbotMzjDDredDyvl0cWnkidhB6pYajFi/Z5KXytSdNtp8wOmeRhuXbZNV9u
nL5PnG0aAk6R8eEUVWOknuBivSQ/tig/5rZ3QDxbL/6IQveCHNAPMRSe13pKZHgP
nzuboqz7TVSehd+aYh4ewEp/8spxUnAftMUT3dyFu56D306vYvZIPt1D0gCdqUxK
dlJEC7gYh16veywl+KtlG+rTHS5y6rVnifET4Wtn9FXTfQ6A2q+ZOw95MdRyDeL5
wwRYxbOzFI5OxOXdaUAk/2klgT98Ajc29MBtaO581/icgPgAyzCbOkw26L/TQecI
8+9csqai8bt7oJ7s0GCqbJmwwJvWz50gJ1HxFD3LEqkqEoHnja5vmwuBs90UFOX5
kkbFg5MoStFPnnViCA0j/1lzgqK7Ycy6DFZ4RAN6Ujn6lW20c7IoD1eDDELHeweY
p3RwyUTzdhqWOey//6hWZfpazcoPJhD4s0Lm24Vp74uSpkoQ/5x28YfBFV+RkD3h
XWJJW7w3p0863ccr+ilSMRmPqvxjINS1kg6ks8ygDOoEVUBamtQpv7ZHAyVMstU8
EQZmAwbLM9fOWatXhs0yUYdHCAZHYP3TIvajReKf32n1V+47UGWi8kA4UL4PtCAQ
i0QrH2QVVhV6sQ26tPPtBcfrGyiP9PX5AGkGod+TrcEG6b0gQgR7DwptBIcusgBJ
H5b8SHQy84i460crbZDmfzpvC0wgei5GimdzBpRV8or8kzOh8YBkkgtS0NCPwCDk
KVdzcIsCxsv3PQYG75r3qiVcCMVlGbrOU6O1iT/E1qaRwG8wQp7+AuW098dV97/M
vD4PfthEMnAg+nT98NoFEFYinU5ZHqMzrrTEUsWzqswAX0aQ/8urj82WdGpDRtVX
zEgtredoBE402+jqOTDqGettGPYclsK7iH/EAS8s1Dxzv1MSjSJJdQ7hsqc6FmM+
+KnDv+bI78I7gSJZEp0yqbDmmJwH5fteM1A2oK8wgSV5rO8vxLU3etEU6On8idYa
hrHxVpWgkrG1zY0/MewMqWICnEjPpre9BPuOaG7DJDCAMWWWeOf+1qhMwZQWNqTF
2NVJlcvRyswRTy1sRGYhaVFP/HEbTUfAQpQGh2uxxcIQf+Qr8blC9ANCYOqSOQEu
dHhCqIIGzog5lh5ej7yJPgmg4nZouQlqm6uELfmVdzSJkn1MH2gqs+5TjFsq+EKK
6kdUE02ZIO2+zBtfMfVzFP2V660OaQNhhiXUQGz94/uOOJXmuSJFUhUmlHsURGO0
iRpro2Dxqsk5DhwuvkE8mH0smqMjofkGjQU1ryXcHBZS+kfUCJ/Oz2w3VTMs35gN
FGoHiQkddr8zzaac+xkjVYAahyRIAtCqbHGH2f2SnHxt379jrnUyDk5xEOTAMCsu
HO1E/vBMv7owRthdEHYq+tITZhTPUfJIZT0W63Zo17dx9S6iFidqGsT28u8cSkWm
NVhO7F5GXqHaYUt5UhetZZMf+KkkdR0Kcgc/+z6ccwdxQ3bM7729Ixef3XGgTEbq
5nw0kj6PiAcpWEkge4km6pmvm858ucrhND/r9QZ5LJZ1O9I2Ix/s/aKInyLhRYhk
TLPAKReTK40WEHPJ1gErmI5Uam5p8Ae5QrpwgzKIdtbvh9cCfF9I5v0qhMSaLd/O
78Rj2S/xqttFLNDn4GMADUW1mBxqpjUJYQsfjSr9pU//n2JatcJA/oYgKdfcEwVM
1s6KchGSEEqRlvcOc1QzlzsZ5qHOLTOaIuH76Qz88pbVe39PzzCi3PP65R3Yaxkj
G1U6G3zaZ2Wuep4dfFJpnY758E6dIqVQxWsukSy4OuxQiGZbcmwAHQ8cxHcJm59O
TAI6ZdW9y0BgFVYBhET+XnR39g95Am3RAk9nSyIKoWkYBUdhKzXQL3TH+sR9KP+n
AHrzwCBG/yyBmOO5BTQy4aVkMuJoA2fMRpNVX4Onjn9Xou9Krgfg7dea+qi8OBS/
28ti4lX6VSFu3r0Nq32WPMJ2rn+2M8D1HJNuxUAUE/6vi9SWupv8ElcCuVJ655rs
hvHsdl9N6gwuV4QNr8IxlFpCvTPN14kPoP1mWWUA/F6GlaVYUCrP3zwQWd5KdBdv
172/TyMHRO12vyUmJ0bTUjFkbyVygB52OiZu6JnURsb4+U+Ekm+vM1q6fdBeMZxW
/VTBo8YMavDeYqvTVrWD5XunGXMf1mkVWQxcyvoyoou75y3f3ZlhwedUUxm/iYES
bD8pkRbUXnB8Wh8hqUv8RrClNOR7PyVAh524pJjWf+ahQXGWUVpvAfFI0LgqYCX6
Hm/4MdEvGeiZVfVIOrk2vLQTpGf7txWrXDB72d/sfoJyTvDumWfdWfmP9M9E5mqN
/PqrkajYZRyjS44XVtxFWeJrIA2O0hb0gIL3Oiwd85wgY7LK3VKm28x9vdx/uRxB
B2UWZM5XjkiuqQs3XLPpzXCcjQfEVaep88Tf3YuIo4JOwMGFwZ3BJQe+kKod6Lrv
myZ9Dv2uEwjYuuYGa/C2EdX4UsPuRS6xvcH3p40F3juUiBWK17GMf2nqjZFvNATV
PGIZod1AARocWwOldONt65COqt7jbEaaPq81kUD+vMW9Hy6abCkH+bqesf18ME3u
3AOVZr435IrrKyN3FZhJehCMj/PZUYkwMCnGhwLcZ6uu2y7SDzU+VahJ0Z2zri9W
hkh2GcVYA5x8ajaKRpR8Z0ZEFF7lhWCOhF+paOkIKkT1Wxt2jBsVbpGElskErf4v
UDWnsuM9WUbQif03PbNhOtdBkQB5YwA0y3bgVIB/xuXRoNIYLoxKg+A1WKPEJKtK
4s8E3PthO0Itbgjh5/vVBVDg1d7C3Tme0SqT2PSRgbeKFlwK9zE1mUwFnDpC3LvY
iJlfdHeRoUpo28q9C3sMIfy+X1ASLE6VNzNxkZg+OJJwBu2ZoAA5+old5Fj52N/1
AjFoC9cT6Upt1osvDjzzazAD2AGEgMDKYKcSEvW8lBfUBkahyXqXe4jqQbqJMx5i
G2op6STN4aEpynO2VRJdbfAUHAHRF6tdDS45/72NwJeH652kZcmRMiT5jxt8paNn
20lSTNrLEPRhS0WlOYkmH/c3dMzecvnHKX2IoCN/nM/fyWhEHeGTP1KV9lmNlc4K
njPkzf42yZRLsw5SwM98aaYuRjr3Oo40vheStxBQKVWUfXbIQq1p6OZdY5ncL+wH
+HamYxDMxFGqpt0yvP+Nfod2U8cbYnIuJ6UHKbXeGJ/g2Q2qgCtroknQhiQeHgUR
Z1lsqVgLeqWbSdrdwqIW7D+uUOlG8t1j+/l1Ubp6KbfYlLSObDBDN3LFvyUO0+mt
ot1oSdaDt0w2oRp4H2mriF86DPA4RDkjYMiUjuZH/vR9ASk8xsgzNUclq37vY3gP
NFSZqyIheYlXgDq2RAcmq99fPNElHr7E1J7fd6VuiwDVZ+kz2SVlrmZp3/hJVV0v
fv9FBaVShxU/lbXKXkau/nQolWWfcvGg2vK0J8vf3pYbH64IF8qm0O2LHYFbfFtp
KefEkbYWTznfetNhNM36neUlbE8iOzranoRvZivmn6RVafL6VtPmVvnXqr2WSnM1
AOnxpRnjVJMQ4sD6F2ZBQeISml/9mbJOIrVgnkUK0ohMnFh2MiAvQZKQe5G486wG
EsWTB842oG4HpLiCZbNxzO0we0BgL2ncY6VdJ85QiGYxlSXgnfW0CBMnJ7Ih3bPN
1uxheaUstzIets4gKdnAKeG1w12qsNQy53zsG0M+AmcrAyKbG8bin8Es1StMuuoD
rE6HV3/PJtTjmjxqt8FNgvSnS9Lfb/YvY6xiAAdN/HgfG2GcjF/6hH07MRKEkbB8
qx3KyXnF5sLMO702qz/i2aG3EBDiPZ7NPjamms0KQLy059I66KaHC1B7JDUnWpzW
vMkgeHwZPmnbS2Yl6wbPO3Tchs31wxcsm0jMb/HqenU+mthBfoiqMhxLJYPDdy+X
OKmBpXUcQAp41whPV93EWSXx8EiSh+ouMQjv5VixKOU/bZmMzLnetKoguQYc7es4
G/BCoq6DWG/6bB4B/pO2T8EFvOnFKjk6tCwqYmhcAXSuDklRWWETqcjrPeepB2ZR
jEO7Wzvs70E8vJZP9bl1mhCuPO2t1UfvZWCi9h0YuON+CfDIl4C1aKluV3lnSlB6
Sh8+XVr+4RmUymmY1MUnNdvmFj3VxbzGLkmIhlQX9RREZYpAWtS0pR8E7FziAjsA
641g/pUqCqhKE99wKTjHXU9UC3SLeWLdDXjxCG3xfc0j4KTVeryO+2qP1y96s8lk
Oa07C41YGw28uSJBnuVrrUFZpMjfseU9wBnvCk4NCJTgE7qT5gepRbdBTq2sLKM7
cA4NJaGJp9vBGrE7ksSE0Fbrv58xJViGySzGS9MI/8YHHn7XaiYhPxTVkM/UoPQQ
WYsYOS+1h1F3tbGHg56JbFISQ8hFz5nZ3gDG4L1/d3n+zVhY3Iig/WKwHdogXzjt
hoG7peWTvVLfOP47FYcTzaLbPefX63DS+f1YhDSgj62k6p5irOTPWwEMlUbX7Qpz
eFURzIvIbegCFt7qOIknaErqd7bY569Zo/7FMdB3K5R+9LLRAoCqQEDDsscSDqfb
Zp1YMRjOp/Z7Q4zdFAGbZ9yGwO5ZGTDa8sXIIOfH8vwjO2Qf1JKa1tq/TvRhAnge
MiCmAGMWJg04PRw6Qh59QCrMvcMiyQdzLvgMiHK2wKFzoisIhWInP7GOeTfbs0U1
G4c5l2Vlz2f4N/Ra22SPxLvAtnDQ537Xs7wizHUDvNakJaJOGRZaDKr9feWKBLgE
P7UepLR+cPVtopvczry8QEWe5NYFUhFKidqYKovORGnJa3nkwdKkSlLVQt+3lyHZ
abuibb1W8j+z9PU+kJ7xDRfu06wSf9lAwAx4DzYHtCfAQLDNnI0F9G2qTN+E+69l
mT2GFNOUE05xcOCEMezoPbwAbnCeS9W1WXHe2CjN7iDViCV5T/u5HJVmLeS/3JC9
IJA+6NPcMzMo6+TSLhLVg3PswAPHu3ltNSkdK3lJqdAZRceRjl0ZX3MNncOjNcpC
E6dyPnsgAAJyIhZLor2L05KJmRjo9YvfJscnnLhCmaXgiyFi6GgnhL3WKbJf6mRy
HkuenFJZezbzMSlNkmOGhHMUdyoxAZuF+cYxg7Q3QzmbKvy9ITIGObaOn/uCKzIm
XxArbJE8UpGOm1dKpUaCzXnEaIl8wo/8sT4tQTM1+LJQ5R7ZU2SaE6DwS/jeLUMl
uappGVTj5le2WAN61b9ZfXQICtOQQ7Mr3JLUw4QOerq/0Uq44RtzVHqQLtnGAuvr
uSk4+pGqUdVtBKDCdbfUEFv3JlaXUZ5ofvH2mXTq9cLvoew5mz/pHJKFc5S+K78v
ECOw69xrNxtJw09J+oGZxYalFu/8f9XBaJtL4VDHn5lXk0bdHuxUlXWXP0u8l7yp
UG+kuTUsz1R9Zi7lws8acyha/V91zmdhFiNJo2om9REN8oG++e+VaSD4XIyJdfg2
I3L8nJMz1Yr2vm8EMfofE/ZUbgbQpRSObnOGNiXkcURImbnpHB6jN0MsKn2MqiKC
ws762C8nSuoiqbNpWRgEeUlg9NxduMa3z7ORbsbifTyqcSbMyLridlacAuKtYQ46
AgQtiXX3TRUfZyCuiGFopp7vIsPQi6dxh6lCRMxEapEQETGkzopX1uttao9LLpUG
5a8PW9KBitxPDEEggS9Wc/SNT3XKzgB7yMqRlbiSHe3fu8NVgA3Q10vk0mVJ2PAC
OPg0btA+mfD1bR/VnLKhZMCWX5XT1bmAVUEOqKw7DlsoT8PikV71eZZceUgRiRgc
keM3LT0OzxJxKwggnJcPcuggp1uacWgeJ3j4Mhh+MZv4L7AaVu7X7cC6x0afxen+
R4mXZ3oMdTBv2SKx4QKVUJgjCwXovfTqclmO4L+31LJVoMOzWOIFDqdPmCjx1qYA
h+Iy3j3dVSrx4QMcXxrtIYbN9nArvQk5kVAiZl8rKBYqiFupRQzS1npkuiIVfYuO
KNwhSbAKSSSKy505UGqh6x9MH0Xkod+yov1ERoHVFVqqY4UpgnrHsFj4rDFaa3JV
7H3MjMLPVO37Vx4CVPnhqLXwzpDQZDUjhZyikYaCjYfSf3j3pVnYtD0CnC6JIjSj
BhgCN1oiGhMcYGKqf2nGKAkkOm9RZo5mrtqvOStv/efirOmDz9l5thQAd8no0IcU
VpYaVehJ1miiJ9hz38I7UwGEsxr5v0cmUZHM1DUumVCwAh9UDXCU4TgcoKWL3KSz
vjNpcp74H2VqN+qJjzTGnM3bfv7/uwY/pYAY3Vo7YhOgYgt+hZlk2j1VpiJvEzGE
9DG71Lxh+e+cAERSZAp8lyDXFGGHJvp19e7dOKLaXHJspkhAWsF4xrb17l1PIH8D
WB7Fm0qf9djCMocX98gBZpy7UA5FO+/6DKY6awD3sJTACQJDHBEg6gZBjMHyo499
s4jM7IN9zXNNGpVg2k5fP2Rzf3yf8GtI7FXZRjKWNmWLUFVAs2YlHUMLEBO3WjL5
aSlMel0469DVwjfJZghPH6hE+anKRj1hmUF9nc/TwSYgY960gvd2Zw8OGjW/k4xy
pZk9MJ9qXXNscEArc/482gQNzn//UhRMVnR1Z/WX6/6ZpnlZWvpvPyWK0mjThkKf
HM+syYVu6Yc5kcOHYBWWuU9GmkT0MrpwlvMJ+SECMMHa+hDbdP+rMyqST80my+G9
aRiIP/5pX6veoLhNxnZJbLitGX4E9BRe4VuC+O3Mpe/+MAn2G/4LsUFpxsuvNVPt
9CeturXXQoHjWg6H7OwwlkTvj5jIyvYOufPz8/Hmnsavc8U1TU86aMIRNxUYBs8N
WiHvafgJoJBA6GSq4mbrPmfTKT1fK6TkyEx5fIzFPQOzTet4JlB3nS8Er5q7a5L1
FaVNSugLXSSIKbA23co8OtDTyEaWzWd6Wy7B4Udwqs7dQjpVy7M9dN0bQIl3lV1o
1ksshlUzDjWtVOguB4eX1iseDnLMADaQsdG05+yhRIchtO0r/qQrPmumHtMVYImp
fvLNs58K2b7AoWib8GKEiqZo2CykjDPZg64WTp3waowjC/D2LhhoVHZJyfHy5rKU
LSX+spiDmGEVT0W85i03prqJIweLzLVtaKCMXQQHm+fIEuhC1p36soySDT4ZCvee
Earx61udYmAMcd/FNwkYb2DZCgCK82MCdXBNOKed26L9t5Lm9DX+2ez6Aim0ukwg
pP9ZPBxGigkXHOOrPBXCQUw1+Q6de+RrgDSoykRYshs6+UNgkWYNH15tKaTw1q/4
MbwPTjFn4wzxbWZia1O8u9vYKypeQASFRVlgnzO9bo1yyVu4wKWs2P1o6AQ1528Z
ieisi254z4qI2gYqBLt2NQWyKODZHzSuu3dlmbZ7XdUXQRKZrLiQp5A+bSzW9cuA
3Gw1krNtm3gsMQIq0w69mHjQjpqM1h+f9pp3NTxn413Dh2l6k1GIBiIJUBII2DVi
d9tNj7DXnN3/SiazC74+ruTMCMy7CUw/g/U+0U0pSoPD/485Y62j1Ek4szueRKGo
DBdRIHnv68U+XuWOelO3E7IUoMCYAYtlpR6+g7n2bKNzJQg6VqkBUc2WsG5kpAy6
tzLtpvosoACh6Y9WTfs8AzP90pTsXsROxJBFmcT29yhNkRxEK/5Sfu50HHmsaTvQ
sRePi2aDZwg1NN+sO9UjWnAUwKBAWzYnUK7K411i2DoKabY8t8AZymZieNDuEbAI
zycOkFne5tU+GmIMm1JUShF7hUE9iDXzjunFz9FZBI21wsLsgXwBXvbf+Ynwn41D
KjvTBy6Lkbag5souWAoSYUz+ALlKiS0JJ15CFuac83olr2s5F7txgP/J/RGxLwK3
SpHg/dHVP/IoZm9aeYZL4FiYZxWvOFOW3gK900LcyZr8QI7W8nilOBZZILdtfrHT
I9UyxI09ijUjsQsy4DD8/YdZduwLEwFTm3FcMydIjudno3mX73LAAKahLxup/Z4G
QN6pdeIA3Lu/DWR5T9Xm/9KujDsGMgvNvF25SdLUWFdb6rnRExXr0xHKTOtmYB9R
/Uqp/lf36AH/xgW75dLlxTp+miXRKVdK+BI/PnRRngWbMiT0BPOwAeBSQziXj1wO
kweVr0jYrsr0k669Fyqwp1Ba4WfKlnzRDb2Vgm/xtuXih8cDPH0WQobmelBl3IXe
6hEH7Ppqx4gG1SDCVN9vDChu4mLVKKrJDBH/bWueCeYPj2XrVahToXBGlLoQS5TQ
+TfDXlCrulMHWUrfdU76cjEVbmmkm27YMzY4mGABgVBKZmkr4O3Xdx258INHhLIi
EmmgK/oy750fm+Q1bRkz7rPJJ4mUCY390ZO+NLmMbUJSP9CIIcMPxLXYBmECPKyU
zTLyFXF8Gw6kGJaYbeEQURF9zxxKoo/o4RRF6djP5WNrOwbOg2d9sgQgQeMq7yl4
M6nB1//qhqSoh+Al60FZ71DyLz0gf66I3CSRDX6VDtQnT03lGFbHT/4UxX/kItgS
ty9WlHgyJTsyP/kel6yYAfDX/sYbHMao2WbKJC9alJ9FjQAC2xaAMN5kRFCg3t46
Qam/ti2y0cyaMnZJ3RZE4izqvBtnELd3+Ce/ncu8Ey8b9n176NnTd+DMKe69bfMs
NvA3N326OQjC/Zy6xX6XaflI3o3q191cRwRRHvc6KhUSo9ONLIg1iiBfSbw839bU
YzMhQB5n+cJfNherbRpmY7WAGthzpvSf0NExfAaaB9K+A6p+65ir+OBR1GzWLARH
m3hbkcRvb0psAVgybQZfVwEhH1Hycwhxrp6EORE2+/orUUiig9U9UoXJH8H8dPKE
Z0WKzsWJq85NVcY94ihf83+D3hFQ6Qa4n/KoVw8dyoTHKRQV0pV1AfWQRjDbd6ar
gnraaBQXVbYrzHTvoxTeHilbuf2lIS4ZlCBH7xzRgV4H3f5AzzYeJNU3Z4rnTwvw
I01a5cywEBmLO3ECQ2OQmRO1NPv317EFayo5s9yWuwUJVEc8tnRmJKCfmqJZM7nX
D2fN8NPNY37qwSfINVsbJi/0f92sn2HS7Bkpx5zPRqr3sPA8Ccf4nnSqi3q0R6Dt
goKdf28nnvq2ASzRgd92X5G53mywbRIHFwp7qKvIA55KWhvlbWsGEDScFdyQTetv
H/VLcsl9p/zNVufldmfTs5oqu1e5sfz73ahXvqTZqOAMcf7YJxoxd5F716/8ZDMe
NWTWfqbkIoXFTh+YbA9ECyFnWPdkMCEc0R8htPOIv51QKqLeHqTTBCsBv1ToDpcq
z3Kh+6sr1OyIk+7REeFVkkUF9CAZ2ZLStMQ31WlkgxC4sjOxou22Hl6GLPCg9yON
KpzY6elz9pSimI6IQEm/WxONbeJ8IJISCkC0/q1Rj2WltNSx5Lucag5jkWQUVncD
etwtGJu1LsPHhShGT41ES3HIQe87jcoaK2oUAi0sDap+gpQoVRHS7l3eTWgpaQVF
g+Z/6xLV54cR5GQO1fGYHhBp/8Jr1HKc3hchqW9FpF2SzmZGjqvO8/UibMK4NaTO
YJKAh/TNpLwtRHv/HsVCLe+x9IKn7EmCf444uS8KIGNdUAIxL5Aat3qnQNvEyCMw
beRpJNedbD2j5aaGoHbbPHNHcxci+ZIExEauyB6KrGyK+nNbLXphL/JimJcwQAnL
0JFslTX6Fo2Qy71XSmdYaB8FkuLpzf0b+lPX8vtJtjwk1Bb1yyaYangoV/tx0d2k
NXE04OhKthtMr4dMAcAJoAXBVxAlOH3o88StCa6e00EFrwOWFwbeVvwXe3KrOWqp
Gwn+Zk+fgX06d26WoqIqMXQsaEJ4kVxbvTVniW+qNvLpot8SrakPixLF07bchT7V
DJI6BV/3xulMryIRGyHJLSjX6qIk5Pay5ZYvGRYj0IVTyYHO373kDPIq2ftN86sK
diOfLqm4f0D16rKmGGOCwB0Evug8fZJ+erR3LxzeU0kJi0XsJSDnhqDT0UPDPwxr
yY6hMVY/BFmXNzpvYHT3yRugy3Ltxl37pIc0W5IejUxtMlKT50/5k2pXbOLwFyKk
X0MmV685eDN82CVsEGl7o/ZcaNsVIMf6yHCSKAbclpdG7WnJHWghmCEiu29JX0FA
2VeDyWE1v4FTrrQgWeoLjz9cbDbAVu5v6VDEkK+L65JurFYeBWNl1Z5XTYlUozue
69XTQpqTFpT6Jv1vXBNqOHuHZT9s4Dvzt9O/33s7qvDqM/53DnWkD6XptxgDF8wi
3kVpM+FUjzDbr8xQY/8PFXwRpcHXstnFqO7CWrVpiRd6KpGSQaxJ2uVv388yaayl
le9vcDhrLg8Dgtrmz9bxjS4OvqXP0KISgyW+PDLnd/wMMkgkIJDCbCxCQ1vN/qco
q6ApY1Qe6RX+CvFRhR+vubKecWqkNwtgK542SCR9fg2TcWTY96lCsIIhGCmnQq+y
AeM62K7v3WB68j1SJsGs+yknpFHibKVUnprcEhyntJOCvZ8Zb1Y0KodPd0wo4b4Z
puCUpWGwGGEd0TASSCwm+9iDbZ8UBtTHb+b9jCRHKH4X9cZMXYXPJ20fTFipOhZY
VcQ6O5CNEg5PRecU3V548gxP9yA61eQ+KldF/psWi+lf9AU0XupJZouJ2EXqdMuU
Cv/K3UJnCy8OvKCcbmk1h64hpkanTwn5TQIb1Id6y8Ue1eFGW5qjK3BoQu81w/Kw
/dsFPV1dliyJOLL7i+edGY/nQgcNS/bLaHkkCozTrKq2cnLTICzYnnxbQLovom3c
koY4R7ofUDI3kcBYJ4y6vatn/rGj/kij/Vmi4O1/MG1WQaV7DPr8qJpAk4Q0B81T
oQYIAAFeNcqhO5h4l6d2aICDMQ5L/wPkbVPQe/OVizlgX6ZRu3yhB/phf0Jd/vMT
leDqZWYmIcOnRLoUxTjg79dsRJhCsU47P4NQ2xeUl0gFMO8kqCvn1hCIvHTVnxSz
PPFwAkoijlCLPzn+O/Bn3HSZ0XZ9H9TH3nuDhHyjiQW4+aFKqchcFAyaN0jHOLU9
n4l9G9n+ri3OOc//beoL6Wqm7EOo4tF86tPhwhz8N+yiS83z84VjSj0YU5Q8VXwM
Epbyc/highCn4bkRw/V7InNA1bjhShTMlOnxNQxK1fOJ34IIBlPlk7IaM16m7429
Ynodj1iRpZiptKCELRViNGHb+KC8QZv+G+6X6KITAK6je1/0c9pUr6xdS22suDD0
lCAuVK8eHzcyfDIEIPcbzOYe7CNSfComNfLko6HyvvCmolioCjkQzqFQ5DvWRUIF
6lrPrpm7iVmB5ns3NHq1aGHxvAvKo/YogaIm7toggZgg/2mQjLcGPLC9PEF5A/Kd
fKQ6zVslLP7lt8keo8lX8b8dU6vZGLS5Ivsw81NWEWLJlSHpNiiQuPlSd4LOOWlf
LEAcxp+ghscFwJmwGEy6BzneQYC7WzPx6WSJlzTB6zd2GmWS7c4SO9Z6RmKShx7q
YQoa3B1BDHOiAPMnBBKfUuC1zz6DGGUGel4oaL/9jD+jwN7G/CP+IUNAQ7IaBQzE
WyAhbdMDkHg/2BJ40e9yGHRNPMwzUoKKVDNOS+VFGphy/oS1CIByFDMITAIq7033
tIed2BzbH2yCqR1p4GUpg9K/T3P1DT2qG408M4s0SjQ///V2jJp2Zs84C7F7dt8H
gRsIfHh1uxuHFtQ5Dika/wkZauzGebfUoDL/WzwPd6pfZiqykPRycLQwJQI2r9qV
DL3LglHAemIzsAn7KkCe1ll71gN8YECBFYC9gO0ig9es8YwhWVRSbloDRpelSPon
trUSvnL+Bz7J38VQVy4evQnGCJgyexIgVa0wW8gkIpPRGWL9fZLlBa9EZ1ro4Xsv
Mg+rgLtMBn+eA68WVt/bB5qEEsp3dFdR2tBPcru2SuZWoe/W1tBG1IFzIcjfoWV6
SzzsW9jpeZVJw8ckO6ECzIZBH57r/QkRev2ps2FYSQGF1nzi9gQspWjC5lTx9pyK
Mf0Uz8r0X9t3Sb6MOyIjz/mxXH7VFxhbF92T+tUyiAk16XzoH3Um8XsC6rjbw3yT
n9pbnwu89idIrIxHZ5rSoYiXIHBKu9u/z2TEQjnfvO5DkHhDWdhbOSBU+7DU8exf
ireEmfLUH1oCiZkiqtQI9zNzAIfc+iX1vwtrNv0toRCdF/YubMcpplOgOuIVkIlv
hbnbbbacHPCbuMtf1RGyrh852eK8bc9s2ZD9ccmMwyFktZc+2eLDdJONSSyJRUTj
TD4RNjVp2+lveZv+jyBFN1hxCqOEHQ+V4deXeCeNOl4h12Qsqe8q71MtHHRcEYHb
5zPDkIT0W2OyDWtL3upmH4EmH79K3S6cxKgNnZiV2d/FVKZM7n5pZZ2yUbmFkmgC
D1y4VU/u1mf49PXDJnRiUxrkGvsLL0HlUsMuZccqrjTEYkfB4/8d/jI9nelI+hdB
WmZoe+AAlY4nhnz2kvMNGYG7g2kkHU4cVHXpcni4nfC5jrWlbD35fCsr5qtCIWJF
38MX0utdH14qoxOnxzJdm/Lw9DxOu3eW2zhPAORL3CB3vTdKM+aCH4x+DLdFbqWq
1m8wI3pmIKGDAFZSZfF/HfUwSfvM1li6epXz5Q4m6hwbKX2ogaho7T7gZ5K0vrx6
5+CrXE5oKCPS6V5LVAu9DFVWHKThl86audSlr8r/6/zraO08wo6c3IUoyWqctOWg
CcxzK2eU7Y6cswdN403Aj8yhA6RneEfTdR8oektV38Nw5tI3vgZnujrFg/ayltCV
iCr+N54Q9hhRX/r0sSPx1hGScxYm/vYDYNc4C5lBHK2760/spTS0affh8kVLUlOT
YD1S3Rz18pfgfOoo/WPW4XI56rLjDQfhzvTZsIrV9W0VpejpazckG6rG+2kn6O7e
5MFAa8x9CD8CneiEq2kQs3ekeBcaKN8KAzgvAn5y3WeFAAc8fLJGEhUyjbX/+Ydg
EBx8UusLCSp10SUk0oae5xHa8vsiWiFRZhSK0AY077P2sgOxCUhGaY305JUGT7xv
bMDnR7bQChCkZvZk5zvCsS/mZcfOqSz2S8bN8n6jIuB1+wjQKMjxzBMmnsCfEI6s
ZBbeSkX8YcIogP2OZfS7zO1iJ6a/k9A6iOud9jgPWPlN30ZRCzbZSgQlDlyJgoH2
u/cXlFeg3aFHhUR9G0OMa/35AonZhTDP3uDQ/XbeHTDV4MzzEbeSXOorKdCp39Io
via938mjqUrMqkyufcWfP4UT3MdF2GzsgFq4RmZcTx3OsfntYMZkpSNsfbTFgBOD
l4nuwZaML5e/yPKjtn1ggBJ/c5OSwLysi3xhjgHBJJQLsaSIKjbtiAoBGS39ekIH
YHdG2HIAzPC424D5z/R391LZaO6W5YWw0nk6pkmCQZv1NcTSbZQw5D/NvByVJFWX
1ayV8yiS1mAug9+T8iW9pc7oCXw3bxu1+JEx2G5k0XNhqnmluYLe3gogH+2v6dn6
9U7/Swhtbtv+TcYNAnh7AqNNv+zVTqLX4zUCa5lQSSRzgryIhBPabmC36GiFWEro
Ebf/kzxmfUB4EjnIphlLbVo0UJIyK45W5wrLuXHOcT9OFx9LM02ptjqd6357652P
CMaRhMh2DATlx8biQANUO9nzZr9BKJyI4XJ7vaGfLldv1TJxB9mQVmGIivxSz6jB
G9NND2vuXzhtO/GeU4AjGv+xU+6F3kIVwvlVrqD51zgl+4gB3VPBqK7CHSUCoy9+
E47aQjmBsF5PPhwivyASIlxcFmfWrG7/XcGMUAYHES17HplAah1qR8RC1UCOzWry
TGxWJViSfrClmSBGCmOyzYlMH3FnXHdIaR1Me7n6+Fr+LN7BTSBc0EWzdHAXj5+H
sTm/QBSYLBwkQAi3ToXmJU6GdmQlQVaINRbXW/QG0L8kFM1Jq5/Nq+Wa9ZjaAJnF
ZYKpv/tjzlG/OOLmOTBMFdTwc5dqUiQZcbmWkoze9GK8ki+Obr8vmwdsZ49x1HBG
wKbKZj2fiZRJU3msIZMOmr3GrffWfmPGh2U0IdjHPS2F0jYTqqMTrnytcYXjXHFb
C8LczB03c7OU1A5dB6uK50UCu3UTfL+ZtV4Wf8nIiIU0K6H8ooZPbz+2Z0lrRhyT
deV9/0M30nnLeGcO9YPf1YqTL08Gb6FQwsfPMv1pc7D0zqH8lL/Jnr9innmmzoAi
zNlvpSfh1ogyfqF7YSzbWucUMXP94pIHHzammbavYNvG3clI8XEkMZtnUOmcKZls
F2OUnztJVr8oLxRV/5MgBcRCG8XVSBG83KQCTokrddXQ3MlqhcZj7kVRHdKwrY3s
P6qrkIzKbIuS8/+AzU/0U7WnLHHdIvFQ1kV5AN5rz0MvjKVrRQ9rVKTRaZ6pECEK
X8YlFE9MPAcXSSgSTZgNgT4yNx+2/wnlFQqCR5aEUgSwbek8jVrH/HTt3vZCxtrD
Xi2u1EX3to5IsgdE8UNKbPfPgmKg39rShIo/Qtnq4dq8T8YqT3FvNk1r9QKea0Z8
dehn6em0rdbxneU6KAln91CVatCHth7zDSuCUT9CsIFvNTjpA0M8MG/NEIMeB28y
H9f9fUIb0+tpqzQsjcW+4432oaM8Eg5Zbce/FISSMllnLxGsNuL10iijftRhHHnB
8b+C0z7Kbhu7bBMhjFdSMW3/UkFgmZR8FsHcWwf5Evq6MC9WhmwNCio25F6lS6Ht
/e/rexopq4RfQBg+cpQLXx8q2uHNoqOTh0iLBEfvZt7CwMn3M6EKJ8lWRjHqpDtr
RbayLLSEWPQeoYMCbjbOBNf4pDJHKmu7ZZqcHUXi84jN9G0122pumfNaY4VjBG6k
T5f7uR9PHRq31iizNncT9UoPA1GBk+IqgqrjuFeeBUVJN/SmiL//ewjEoj4A0MQs
R6Yh15Pl4TcAgxygy2WPNvI2pHN5NaPfPbx0iuvFdu0HLUWkCqRBQ+KpPRuN5JI1
PSSuNop8MI0icMkd17J0x9sZcj1c1FeH+/X+OHyhTnvJ5w1KH8upEb5p9yo/hfTj
4hGRZrSqIh1EPIP34clegT6Et8SOR93SQ9Bubiuf3gxAanNr0Oyd+F+xwtj5lhEx
+agCOZEHCVUDjR4lT+YoTuZA1KWZFbYdkyy6GuqMDhBw5bhKG0Dsmk3CuRHbTBmq
i2rlJNUxH5nAiCYXUkqY2OK3fBGi0JLcaMGUfzm8YPboiOhPQUmV8Ur5CUqOQbIC
ufwOQYYe3K0Ohcwh72cSBz5q42bheGYq0YlupEiOM6zyD8X2mwBFri4AWUQQrmvk
XSVk842QDM7PpbcMuqxeAJ0Q5Lcz2Nv4Ekf344wYWacAueQXOZh04+x+9GQe5HCp
9i4K9aSXMsezvdTg51GpA/J3lrOs4Rv2SHC+X8pCdh/3/AOMr0VWsHmp8wWnYtmf
AOBcLlcD9nSPwbuc63VJsfS7xQI2O+YQV5pDXy0+lqNReP4M1PqUTCAM7ihrHS2F
3C6LI1qmyEzezczTRivm5xxgKiD9z63+zsfhZRhBKte7oYwaIXggd55bu7q7FA7/
rcOwGRdcd/nlH0Qtg/EzAfYcPKtX1CXb5T54tO5WR23Pp5t0+7mCpq1TKkJ6axCF
tMk/dUagKha1WI+PnXvDGNidlwelk9y0TIsJPw4L8MI1tJaFaN1NxQQHNL395+xE
jWFlxJuaoYwJakRJAVmJ2Qd0eQYuvSoJVbAhlcEOspFviUrOpUFM7wqQO1ZDmXVX
iDi0WXQYVJyCeQNfS1smY1dpsbu6W22nKECTPcPfHt3wwJv18E2CA+oobFyNcSoL
QyBhjOpuJrnXsjtEhl1mRbJ88EqMLMOHvPbg57utdNUpBFCkuQOAhG6XF2cmWot/
gAxtIU5alJivajSnPoFGPfzdy9KbGditpzRy6mN6CEljnbaDDoJZe+xvgtbzrIDZ
FExGnk9wZVtGcZVzCYzxmjX4fs1ACs6Sgqio0P8+QBueTwTk2oayi9OOSfjekU4Q
PSckvly3rA0CbXN2lOcUGdDjftrcEzuKHriWUSm+wYDqC9g/mqQkZmCM2lqzBtER
LMgIZR9wLgwweK+OY28JZEcOPXAFexdWvR2s65PXv2cg3MRUwO18cj1vRJHQhWS3
MMbFNQnQ383dLwb0qONiH0pW9KNAtUizessCOy/yYVwAIjha/faZuDH26FfobKTH
j3qPit3TIDdqnL0VMZjhKNqppG6zPP6IEALYJJZfwPkx9E4hxqXPB03y/caOF8be
CPnFDblCmPaSrIEhi1suJgcdDw2wPKBzPteIJMrYX3OeDKnfAnlAu9mahl3Fo5kA
ukIAfc2zbhflCJO1GjXb/e+8ug02TQQ9LETjJBdShBd5BzRn0+dEEtOAUc5HUvyz
HMMPQ0Y1NC3s4zTOJEigQhFxE7yJCFJvk23jdTJ3ZPTMtO1ET+ObO2lsmS59VMB0
qWORROUgpWtBAXViDR20bgsM4/UzFEgkpVeV4bPjWPItwfQW+CnezmhpTkSI0ZyB
p20gV9xI+NmblQnUuUeoF2apnqrQNIY4PYePXdVTL4eg0RusFTt2Vn9NLiwYekrE
0M9xNmE8fVUXKX8XmXgxNY/V9oG4h+jQIutMsmCQTVfmKpfKHqvbm05C6l1xUTVf
PRqL+Bvj4nnXo39FEfZVdFNRM7roTwdYe0hJ5y+YtSFs9xRPWstaLkStgAOXRnk8
D5+woqbRaKfwkdEdEndkiX9Nt3w0xEe8mxD8CNBlYSB91q0msJgVtCfdJTwX3HEO
s5krb2XxStxCAeXSzUzuUzF1CWB8vsnAn+Muoeojlv/aY1O3oRTEaI3hGn/DPRSt
XqEKplyNCzI1BecFKgafHZhp79cI4S4BStOxCK6gfPUq3B8oOr545ZIGTIsWwa0U
OTmTNq6g2OKkNlzRZIE+UaNkfE2IOqB1e+dYpdni9mNRTWKM1lD9ini3glfeHQ45
GMM0dOCmVBN2W9EEyOx9RPK2ZCehnyAz+gtmotp0jkjOo4DHpQX6qjjnB1JUiKyz
zpqmDBQl1aDgtNeKnS6CDsYZGbZMCneR+bYLNL921T38+dRKfR4r9XwhrnAAxVI3
yqLnY9/ntu2SpkBWoxgpYi54AvNLt33xKn7iQzAK0ydZn6mbEVUVrvakuyTCwSWc
EIC4MQA9xF0YfYikQUI+OkCuTsI6wzYij4eOozA7/n6fRqt63kn59Z8xO4zlHzw1
EJgrTJfLHBfdesbXY7Gz+Foc+cjSMOin/69q1powuzFjnFlXS+LQNCGgVq1gCHKQ
vd6lAOF9ssN3bPYN46TL7siJLTdDKodqPBlI9ilKA6qpOZxin684Xffao7KkbO2r
c6zSCsfhhuoaudb+CO0wXj/1mRZre6ZFDTwfVWApMmerTo8p87Mt/5bdrKuBmanT
n/0KNiDoRFRVGzuNNAEVdBJVmJlv7ncighEyO8JP96HeTqHlD7v7FoAcykRB1yUD
cDm8gvaNQv/Vez1xOcsB4M7zJ58Bo8zRhIaXIRIsFfkNe9vSz3Mp0KEiP8Bs6Zw2
jTWYcqIkwhZvH2CDkOO8dpquBb2dwWJhLeMhd53BnbN5avkN7i+kqaRzH0R6/Gtw
dkXqtzbUw351Uli7CJDi4xA7QRr3PVENP8k37t+wfBcKmd8N2i5UBJSV1xZHjLRN
YB6xtMCH/EjETpMaHuj2PYvwOXIpLjzoMM8XFB9OaiUGIb8J2Q2wBLreYPj/L/0v
lNBCkTN4Y+/ECXODm+jSuTOJz/bRyJROdzgkWPj5g8RgRAGxWFoOgq3HN5h/HGU+
ZCu1ENsjM3cXa4A91l96kNMsYd8s5Jtj8Glk7wU7gi39D39jQCcK/mguG+zvPsJx
++6rTf+Dz6UY66PTHoBDocfNYKxJo9T1gXkb+TdC0YpfxkpCMY9cxTlMhT+gxFWI
nVA+xkLfL/RGaV6jps8+6F6IhIy5aXpNhRVNdVlcj9MuM0hUVigMowI5My1+zAna
4a2TbLD+UWJS/CtBwPnXtdwsn94px5Waz85gfUdCPH8Pgbd+KfDn/m/xsXO391g3
Q3MMuLiB/olA3JokBMvt4d27EHCAhj37ss5SYNJwfTTOEFZ4e+GuBNiIOnLFtZAo
46S6ukz+wiRe1ni0BlWyrmyLxcN4BgWK7TgXT4z+SQO+0MJf58hp31lK+0BZk9rH
GXAAbZdgjgY1R4KyvDuQ2m2wR6+TeElvwMoTBwWcdYpLTvfYIKK1RuSTrA1qLd5B
rx733DRBsCg28SsvWDHte0ZZcj9F/m2irXF6clWGuAlLHteP4yyaOOy1CvwzUI2e
tIRiIjQVQXCgTQupwGuj6TmZuHF/J4T3Noml8nYNPao/Xp353y6a5dq5Vm1c5mz0
IFok14nVb+dXrHObgPVNqbDHfvZF4OraZpsEgId3Q6SSCnV7UOogVudKWTvvxdvV
rwwgsiklvv4mpIyX6rzewQFybE1V4ypCCq0OjulNgO+G8Vtg6KijKAgzz4pkClpo
FzTcvqD4ElIh9tsPEhHOCwp8aBtmppk3/QUtTqh3m5vI5Y68JaQEbIixi+Tp5udS
Y9vsaOUpxZ3i5VGHH0rp8AcJAbDkvJC4nm9+jRlirQx9OgxlOLgvytX4othna0l3
p66PUNCS0hguQqBd7jS6Jm3/xiNdLUN3ZpYpq8SpvsbK+ncrlIABlUCydLW+vtfC
JeEVZb84KNyDHN65vroNj5daG0lpsFlAklQ40afC6HuegT93IHtxfyg1bATNKFo4
HAGsCC07hrp2vLOFabZ/NBVMRsgtp5t5pIHH7yCgubntxEziIGq8TYTxSbfLpa4I
cgjNCsCLoknyKtZ9/eZdJ67dbuMdETIMNglOpG9toorLEaMfuEQVK5WZOyX9dKkz
GbGANwSIfcC/B8iPQ/WSevYTmC7v/+P2H63tKnKFWDyKS3RgGp9GMXlT5cDPT4aG
ywdRBQvVxcBfH00xydJKpUySRurcRYqUDwi1GjZC6pB1n4RroYK4ylTRBPMWdQAZ
R4ojf6P31t0wSwR3CdxgrBSP4BccdH/YqUePIF1GlIOhRDPOU78r+rmkXhJRFGI9
euLObVmKHUTf0REyzVLEL0mZBbqwCpI6sG0Aj+GvinTNZbhsMOe7GF+0PQk9fGR2
zDT6q+FyoRORpQhy84d4/vwvzlSxjKUX/XVPjDYaOpGO9BV32iO7qHZuobRgOPqn
BRl7tc/XOTFEcLwym9PE4AXEt4JFKc4Gc4uWr8n7mx22Kq+GbRyMA/dIuo9hX/Ue
5qErMuAIS3oJTghZXrga48A73hG+MurS9UpIdeSCdh5NkmVKekIaSp6dOy+597Q4
FoBZuDo4M7mGGNIWGWHcEvC4hbk0D9mQq1SSLsw6Z4s03Tw8Tt//UmT6gN7paS7L
XUaOfqLUvMC0I+j40RpYWM1dBCjVD3bg6Tv/clhTVB46eA2V4yHg3ojhF/zlOaFV
iN763rAO0PI6WCYHeTfBrQHpKEI9aXwwhPkr9HQ5gdpi6MqIRx9TSXXjL84mItWU
uLSmBhebaI0OggTybeokjH/Sd2iRaQaT/PukLWviYAGRqIqdBxKHbBx5F65bWycI
HFeLdpAXOQeMp6AkSKta9TlRz1zJpXZdZqpgWbR0WY/+FihdAGRe4RSV7u0RJRoG
A/tgGd4K5JeOw2fSb0hsvfiHC36wTBrExPX9ZMzQVQwyPmp+xf4ExT8N9fVmi6xI
TkbdSx87IhLz4CAvuuwdCPxESeozQLAlJ/94s+E92JXsU/ggHK0rOVFiZDpfYFK/
imnRB4eNpZJbW/x4yuSUptB0CPl2LlNzc+7+xtR3ahjr6yEA2gWos7N7nXFqJJZT
vP+4noDKxzfQ++jBBhSvWwpv+QRyosbGm2heIk3+hN8lRHiPAd/sVndBDZ/7DJNB
78uFzo3yzLGVTcubjemZxGnGglTNT2YH5D6CgtTvzwk/BDUN7yoO+zcrqux7WOCf
TQqu0nAD+rsioBFeD6WbLShTvD8wbXbTxJrATcStTqZ8MDsLkB/O3u/hLQzTBv/S
tL6gTCn/YCwvy6z1pJGHv8WE875aPFg9cQUKqpt0xbKxnkMdri9d0jk/FB4Mfgc6
W0RbzyPFCgVja+W6LdAdjFBYXpkbwOfpVrWCMlkL8poSROMnNxwQWiWpd0wmlmy5
NjTAc1ETfPHQusTX3xYbQgL9xEDOi5NTHuBFrkHOC6QmZcHOIObBtkqq2XPjwmku
i4VftQRVAkAmBlSn16UVMAZHIeqhfHdn/JPUS0cFjnJzCnv6VdVMfwxofuqQZCaf
WNYTDJk5LW8T3dyyjC67lGCBCWWEGRFZbWGj13oJwJN8QT1LiCysRmI0LzrjuAiV
4ZnWPg6iell0kceyGoi49dfTDebVgP8Fxmgi5IV6HpcaYuXU1UIgTBjo5k8mueTo
GKMsO0uI4b/dgIVWXzRD5ZbGnJu9627nOoZ8kSYXizJ5fGWJrW2ozHJIAaViJHEw
X/hGhExu2WiYhIJsyYf4NcMQa3fhhCwC37a2YE96DiiVbNh++A9e+tjGYkWvYZgu
kusXQzpy7x4VEJJ0qjEWG5BbbFaiAIZRssA2o6jfMvLpRtuOf9anulyN7EwvaP/n
piKej8nzsYCeWqiM86/UaFKUwik/15m6yFgX6IH4g3Ala3Waxn+aY5jHbfSbSljE
ScdUFLiuexd6cggGtyxnERYqb+FFmKgecnHVEyeersPMRbtK0sNISTEljEX8G1Tz
tcnV4dXV6WKS5gdhg5f4gXZqlmOV7L63etAoM3LcQXKOa2DfF8SKUKXoXiuNGx5/
uKHcBeGJoHRlcwqnQ7ZwwcUlVg6RU3Ez0vjOWakgNn/B/Pb+HU/PojsT4NPMSDdb
s8hvKCDNqSReehdanxWXqvHmC9auXw4CE2zctVAhIRsTDhD9rRJdTzg6IZnS56pJ
veFsM1avxdOLmeCruCe+8+hrUUR+oz4EYwCCLhnUjBUvc/OLaNaH9sWQGwbpmflq
y2yyD3E91ICRjB+l5eq/c/iAZAJm8J1XuzUjaR9NGyo/ygSeoP/kgjRV8vrsQbaW
AUL/uKCfJwN8cSE9+5BI2yds4Rh9sdgmDa4tDEiSV03SkJ1fH71uFAyufsJLuU60
Q65hE058tiJqm2Vc0wdmdFJoWY8tSDlbXvaTvUnamfDx4GGigdWEZCCdKfA1mPqy
/3/PRkTxvtn5C1uCOkqW089eLJ9wru/LQO00p9zWL0Wzgz+ziD6uEJTA11dgF2FF
mCC6Z3fzBxloiErdT6shoTbqwf9tOwD/AuWRn7fPkt3ZAzxmkeqRjMKpWnIqoVrg
y8e3KU0mp/A8QsbkUxUIyRzYy6fm6s4xG3+/c8GW+WbYSvEGY+05CFCODK9chuMM
WNQ75hxKhBMVniEvspcbJ1RbLXE4tPpgXYO7Ls2E83NujLYixJjlYkVSDwiho31r
21kyjN0US1IOM2rZ3lStxOCgBqTAU9HCu4ryTz9Rf4yN159nQjldShrhXAGJpyEF
hrLZj3p85Z3bMphS9vLZFOfz38DxgHqiqHCg8w5WSUgb2IDJzEgSk5tuAEvbDVMf
FgHLgiiv/Mrs5IzhuR0GAFPEzYVP73FIryGlghGe0uRvxOhKEu6hDO7egujEBEX/
F+vmYVvv4lGObuDPA/CmHc57PX7znTh/M04jiXlJiq8NoWCBiWCaw7al6DbT0qL6
89qyDRVmbipv2a/lHdFwYYMpbb1phRwNWP2sInHuA7SUVpI3Et4/aUOjAfbBYiOS
g0vwY4LIi7+8h4Nrp7NzRlL7eSE90i9lwUVAnR712E5pMdbUAdmJ7CI3xo257m/t
BsrzAcroHbMrLCLFquSAM9UXU8Ko7SAJMVjn9nuF8AbHm1p+l2mCnNAUJrK9IuAH
nxvgJlix4nxJ1cl1wW/TUygT39fXYrKHeD3J9A3QL0KWvbiWRfI0wf7SWBsgHEOv
gfVJYsaHLkESKLHs2wU0pGPCMIzzS/9ogvujVDwrXlQ2vC5Q4grAdwTa+KU65TQI
aM3C8OPpcKN64lW0TRt9OiEnM+iZD12mCru/uqDPWMzltQcacSi4vrfZLFrbov1O
L32nijCGeSx81tfqhkeuIN2ezccKo+wUs4oerBWRaejTuKpOhcMWuNiIYmFR7JHS
VKYAwXM2+iOXW1/NIbncegFw+x96QGosPRIg3kx/ZFiLj3wZbJcYFHESkm3+HoKY
ywbs4TcYVC69XsWrDIzrJkL4XZtdJ/kLUwWkkxmZKUIeXM/yKJJW3tbXHj+3mt2u
Zhlv33gUd4hNRz94gii+CTOnpFor6tEa+QhiPAji8g3BbmiznF/9Xij7Ie6MX8b6
cexOGYd2OIotk2XK292PSO725oQEm0r3ijeNE1TWCRwEEs5+Z1qJy0OnJrcIqgmV
be7eKGOlqawM/BYBLvYDacXw238QydqrBn2S1tcybR4WxvaMGk6EGh2t7TBKNEB9
rKtxcyQjQPA+TovJWRkkvnIdgG2YgvNjXchiEIC1EpRzPPLg/eRNR2QlAODGTFBN
07wMQ8aqYDi8QP+lAU2d+65Ib1bk1uFJn4PwFzp7IqXq8/xz3/xt4KaWctUuuFNi
sX5HDcfP7Z+4pOg2I4k6kYAEKF9g0I+zi58vu46JPDpiHSgpnispKfdNgwjiKONZ
shSyaUao0GY83t5NFuKrfcX5AvN67ZT1TFMA7z0pAhlBPWpZOEEEiXJm9E1vEnOQ
oDtUbSI83oQjoMnAGfwXHC1rQVPSlgcWdzEClYSIqGQIDagfrPGPnAhMFw5iLp8K
b0yd7xCg2P1bjU8+xWQS0x4wyEBheRJYSc7+5mm/P3rzj2HJKl7hwUIrabHAgBCY
vCyxF5+wf/eceRJsIfIHsrakdDASryYXWr7VStA1dB/NSDng2HwkhtRgxCHHkqEu
TpuLWtNBCBlwZuQGf57vC2fdxsbv6MZK1Yewtsksma/MMnFmPZGYTizGEj6Fv4x9
EJsWOYzoRz1r0Eek9tHEdD8W502V7jpG/x4E6L6oAabNkKHOJ3D7jSPZUkq+uLif
29TfkSB3PBKzTg0nTlCqWjSKSpwKIxD9HcGtHfr/A8N0/oZUCy2nYwDLE6P93mkN
ezWJu6j0coEyBn1zODXzFPfi9J1mARqW5X1nW+7HqAs8vjsqtarMwbolZ07dzbBl
tEun0dSbGnU8KpQdag02tut74W3sYCXqiJQHRbS7L+FxiyWvSFvYopuOSivQ9q7o
7tuvJvB+ZGO8SdkY15ScbrdYayh6Xsy2N17jNntB4S02FZdrnnjWUEj8057tIoSB
ae0bObJcTnQL5TeYF0iPuMos+DSvOrJTxyaUhzKBBEDlICItphwDNA/UuPJ44fH8
8jIJf4Ut1NX5pp3OunS7fCS5rX373o3W5Koxpd0txjsS8ZtBfxBk32pox2/mDgQN
o/o5/kfPO2PROqw2nejjq8JtQUE3zBsN5b1pZ5PEPv4R76H7cyXcobv9hZDRL8Bz
2jo/bPRXyi0z/rkCK3L9FizCdjGFMIhbvieuk5Pp4oIr74WMUhNwnZ5R+fazus2A
rhHuXPDfuiUguATkHMFbmuNqCGDtN/9+I3xfDBJSUS6KOv6Opzh/dCZKw22jA/2T
ONLhUR2S9GtBJAB7L4y2g2D79lw1AulRteOYedwKTSvUvUsCaVclHK99uww9Qfgr
S6dn7Y9KJlGOb5+R23bZlwJdLow670tHsBgyavES6vsl4y4Aqmww+y3gTBOf5t18
qapffhiLbAw2RtORqPFYwkLWWXjF4445KywrY6YqNewOH1LB4KMZPQAVjroDuuj2
y4pkjlCbvBKQ4NOmvQaXtYWoy86+vrMwrwOd7T/HKSTK6r6JYXrLvcdil7szhIRu
26LtzT0cmhoqeSZkyWg4mxa6QmUTQeg/2SUJlSvDUqqUHUGAshlEwcyXHl03SKS/
66hqrNiCAQ3xPgmL95yysruiROuX5wOes3kBaRg2P/E+rG+xDXVNmF0ZEfcJhzdz
mt90YJzMtxzTFdqm3tcDv4MqSxVBndVpoQvHSNykJKfjTa1IEko85mLM8T9My2OH
/4fDwBPWBajvX/vMvyBj+kipH8uiI+39/s0PLSimqiM0rvNYkRoUd4KeYXzLV3jc
vNBP0tK9YtYnWjFVaGEtElT/R7Rq82SABVzk5afrgGYJa+PrMNdNTyx4TUxeq07y
7xBryv50WDvPKH6uzkWRffBifxhm/Os8SfOx/qrpazESGJiHlUM6ThegTcLO60u6
f8/nwYGxmy/xAx5THUiz67Xq2mniJZ0Un2NG91j32kJJUDYZRDYzjBnQvm5wxmYK
QasIoN3XZyR3HIkij8Z1K0rmZc4DCQ501al6oaVs8pQn+tHA728Sv0qM5RRgS9ru
HV5FcM5CklTJfQRVhc25gRV+vHRmL7qEYkBTpbsZamIls4L6o1A8FttLIyJd5QdB
uwEJZsBUxKhwS1i0IuNTQ9eWm0HoS8WoUcrR76jAOZS7rg81gl6oCbefMygA5VjR
a2w1l6iBOytIQ4m+70BAnqm9btD/rpRwHbPGE/6A6n+qWidoXF87xIU9NNIYS43G
nWY4UUmgdPoKYsju7ZxUnS3V9Ie6DLmOUFY0VDkIvMsyBvFeP2D+b48GA+r7AlOg
f4lBdbEYRXDod5nxwJ6WxhBf6Ge5YBGR+HX8MfGE6wryprwPtputXszDD7nh0gak
6C50cU6fKudB110G4i54qweFQ5j60qKeEU1L5trPJPv9Bxv8TBwqe1F0K0nboeeD
JUWvaL0/yZGfguBoWmDVKQZIB0BkeI0sBsjrbnQVeekiP1lUmcVs7XNYVp2i7Vs/
9Rek8Pi9TUiiz3FNgTcQNnZi4IokjoZ7VP6/1rfS5PA+6/i02nOXztfLW8iDOQzt
6wWgxCht6el0ZC6T2gPaL4ROzxuohxkvoZT/bpuRO2wR36zl2P8qZSzRE+jyBCWc
fN2g0SovfQzk4S0Y7+vm8GsJpsHjgotQ+MnH7JamYtWYk23aDBgkuZJpYs6AUz0B
YjThVN74xhxgcNeiBEdRFea6jReCEAVmNk7oqtdxjpk1v6uoH6RGjul+jg2+hbdH
zMNwd9rIMK3sjkm8YbDiVwOBJ3i4Ze9lAV/Pevf87Zyx/7eUAXlxTCRz0fMPHIN1
YW79wuETvmHWBvxX1RvZveeYRvjWYJ/OBf6hRW27ek/pbTh2XW/Yh0CfeobZfqiX
RSekgcjDGzSnM4Jh17F7gnFxUbBf5IORs2ENNphyAPKqVVBseWU1yN+Lh/M9AB3Q
aKFRU2kk+B8j/VR6LeQqudo6WBEPfDv4UgEPa/Qx66yzFHUymr0Yfw808YOIxUfK
TOVqwXHLvQakjzW/hebkvyXS/t9oOc0iHtIGjh//fTukLb/KPH7wCpk62nCGLfoj
C1Y4JY55ASobrEB08JbV0vVqN/ztHVGlKmvLpgX48nqjyuk2QDFP+drSjyyGyAlJ
sHFTTeYbZHz8jKHJxo99yT9q8bh/oRGABzQ67bL9sYV1ME0DeKrudJ2bFg4Dz4dd
s6AvKB2Pqj1S87uRItsHSpo/V6lbpeJMFlEanRMd+HGC3BetxVAHDajEhsBwzf9P
21RpGUXrE3GpchuOfOWdcFsHv3QL+MP/3Yd/YxVw8qhrubnWd0GnEgQDZqwVebwm
8sIR74M6cPRFNviRhT7TwTtLLPhf3/2ujQ2yWGNtrV1A5sJUrqCV1wx9cJwPUz4U
/sm6gLACQlzDopHffkJN0lPGYXsIS5bL1fvqfcC06odSQxae8T6z7k5SbszC5gL1
EO1W4WnSyGrxokNhmy1P7cOWuhH7uuhg0fNUQn1iureoCvOqkLL9pK9VlNYYZQCu
BLfTW9aU2//2ETWq4z3GEJzgrPh8jtMpYRl03WYnTZTolkqdY6UaxUs5nDuvYV1M
+urEoh9iSQuCs0NEXKVQZXhCRcrk5OFKhjJJhjqzHxgwiNU2wXgxxTGcbMMc282/
FJN2SHr8X/1uU/EZpumEtKbNvNqKDB2iq2uRPfAPk6A0hpO7QuKYo/zW0M64RIor
ArHn74OzKkoZw+UBA+lUM/sdr0E4M5gBtekLZXfw6rh2aSEDzlESYeW7ErTOuQ2V
dxeIP6Jycs+SRqrWBgMT9jrjsTSfcZ74lriTuE5uWhVVFnNNjUmaZ/QgKt/sFlyf
SNoqVfn4enYApXteh7fHP8Nfni3O/WFr7gOL1HnzsdizoHvjC3etj4HsiKry9huD
lhZy/XSiad3pAkR8RnZhdrXfpb4jrnDZMIUvY0BQ6F4Vd+YJ0SyJ0F70FluM7rQ+
vDuyiSE1Rgpsm7uD1x8yk7MGgrPS/ONQDt1snBNNF3hWFl3ownP8tmIxOtxxRJde
bwzXcEJ8iIAHRR7JOuPgZfDCQps8Izr9XEj2Ug5qjk/JHmFtw8BHC094W/VkgZGQ
aZzBZ4wb+kQ5YqTkKZehdqpYa/kp75r4zAk7jzOnGil9K4aamqCAkxgN8Bd2zk2w
cNGdY4fRq7pxop0s6viNSLUY6q+9xO6iXjMJxIk/Ag66q5j79ZoMF/XLfrfZkDi7
DQB0ZGJBb7LRQEp2K5dPuSvbzC/H1c9esoG6XEMODBym1VAi1+V8Q0XVQ0Ebin4S
AzkKoqZ4UJ/D6Sxy2foNid5RoZmK6m4FtT0qWVQAyZzpu+LJyUoCLCw9uy/3vzcl
HKLMNQof0HXePfjwj5jkdoVZI6+9xIe/RJOY8Mz0GvpL1aa0pHeMQX0DFXp7rdeb
l+YogwjX6pouJOnxxawqtoIUP+O0ztpxpK553n+hDachDoY03jRYXJdvPrYstCc+
R/KKgHt1QP8dRwBRgK78TlqgqDCT1i6BEatn+bVb9PKGbCxketIe2nlbul3+N+Zj
Fem7GuJ9lwK68tpn3XSBICMKjKhydgSiXFehNU43HnBltMxftcdiW9USemLEQ4z9
g0qNQtbZv8qKmPkwm4Hxg8FIj4U/r7KaWep2GDb4769blDChONmKtwgzEYofsiXx
srGg0O9eZXg2l1LOki8m4zH6MaruGAn6TsSejmyJTbKnCRSoFcD7AV+NRV/1Ta6I
ZIHgU8HZFK8/W1d5SrW5jCrVFTuFsM1NdBEKrou1C0UKESZHSsUKOCOrSBIERZeb
NBxQRT2t241OcusWO1AvKEP3BYsiQXFYYm61UzoMDft22tFT2jPPrfdYv7YYDBkQ
cZwjtSQrZgnJJ3VoNqLYAYu9dLmhFZwtyEsIZtkcBJT2M7dWg/w3qkMfOYXaBOIv
1iYmAZh9QWcZvvexC030UsK3BUdr8GCt2dY0k7cBugyN6kAmFH1gBJ/HJw+AdWm8
e4m9B2paioCn4VPpj1ecNh0/zIiJvdZzFADVMXSg16K1XAzbBKcfpQGONwDmC4GH
A4EmbUgb5YKchNlDGU/ra6vzAEqgMZ1MhVYhMANq7Y73Q3ZsbO2Rk452m6wCAnyh
PMrXdNgTWfZwSd1I/mgxZrNU6auEIRgFaMSZdkkJW95L3UridGUXweGywguJ6vCb
ORrGWvzpRb+KOFgNsDUWrsmPvWjlkd5Plb/ewLujkTx2la1NSDqDUPfzfSW7b02f
Miq/zmQzhUYuoA0uZB8eKspWNtd32ZjpfKIknoXoQ0VjTYDgEMs8XKZILAOhvy5I
jtupovF7H6bqLb8OyQoD7+c5Qalt7G2bOIZUT/STBq9ADITmsaM8Do9gP1jFpNig
uYV04sgzNsJf2hZF15dP7wDCshlxNL3LLzDTwR2L2/ANCh14MbrxnwLeSvejZJl2
EkIcDrVRrlUA3gydZyG9DS+4KziJCN/LCKqXJs1mXfkHcfnQGaoSvunXHeMDCrm1
kPEGS9sGwlOpQg5J27O+mD2pkRbq3kNkPrz6y42FzEB+r6Z0w/vfOGso6BIQ4OtF
Y1ZN3ya4d/uHV0EhYIeiV+wkTP1/SyUvNCXizkywiXLMDAdAnc0kEpta3Fw4qUL6
KDdvPPDVjUvlaQfh33TmjaL7y35rckzD+gWlEhaNSQAX0j8TrviuMfUws9+5A+ix
T9BzRIduQWrJATRmohCGyucqretDEoVRmPYEF5RVrRWGVR3s1Fqr4YGWWilk5mim
z4nYctKhFwVNKvwVArsaXRgG5TmUwqcc9iw0Np+nWU5KG94Q/soOELzArBjbmpLx
rkVSVVBroVltZN9uSi+JNi2HzpChuJbsDFAnzC8a58ZZnK5OKfSW/W73ULX2031/
bn6Gd/2ohwksPF8db0F259vkca6gWaeMiQktosOFK8OBxdcY3bwP5OLTplcigafy
sLkhxZcJRx/d9JZUFR42VeHlIDirH1Mvimhg3NR/RK9TebV+LvRgAh1v90wY95Jf
7qZsfvCZLUQbKv8DplIpd7JS2/2SY594qzpJ/MWVPMjC3qbzV+fbdOz+DDrb2Isu
PNxezdwDXI+GtnYsIkBZJQ78Qqy8akxNOdbIg10xUq/4Ppi9KmwMw3OAD/1Pm+mb
Z0gy8T2ValVs2VLuQF/za62lp1L2M7IHqZT8us93ftj4a+PQKfLvi7xrpicLa5n9
uP8qCS8QtzHXA9De/K75fgKDwBitg7rA8WrfRrjPH4LWaZZm+5GzNMRFU+CIToRP
NP6jeP4WrCCMDc4d84SyevIHXWURugTQC2UgiYmSnmkdIAG/kMLKwql5djc6iJ7n
P4xrqkJ5uPmYQcQCMlKMjsT7NqFayru0Iz9vonkKqd32Z/i9vCRUPGznXDn0hefN
KBNA5Vuzt01VPI9Hwy1kH1KFaBhmCyyNS1EgOik8uAjqqVTBL/1hDFAajhCAuE+j
wfbp+zyegjqlp9j9YyYMr8vkQHdrMcrOcOFFhGDcVGWLWkHZVOUtO++nrsmETpxy
AkKbqrOK+4c/gNkRgJPTP9T26qcfJdlv2aoC6GPlcAE6+u+4L4sI20yEfb/nOG9Z
E2FVH9fGAZK/Xmcu8foOcK0uEfJcXZIOs7R2vmWTnD0sNumHab0+oYNl/nIXRgdm
bUJrbHyxyCKISsWTdIzfbkQXpPvah3Eai5SbXbG83c0UXW6mVFwYRU77jGvdblb/
qb2Ix1vzJ+YE9rQsPOM5m4S8n1gxAYGaCovEUjof1ZeCSbGhNmmGlo3W3ICJXnyy
hhIMeR6Emj4wtuwuwl8t0cRji1iOwR6pq5r0v38RFI1pMsVBVWkNi6GKapBTfeB1
TwN3+SUsdOFfTYoGqvX3LcBhN85a/swJEtsZpoeHnFz45RXclq8Kb0mDoqLUImkj
gNRjOgQTh7g42IdlOnIGeT/2mgY21BSYakUR8duOP5DXv1OljrQs0EXNC0suLrzR
rM1gkN1pMacAR57PAFew8KNs13vR0Z2VIY2Zu28lch7DCAnBskkq8GHaLj9SnFfr
8A9I+ksfVpp69nTZt2xeF3xm1WsJbRLv++d4ANti/y7V4rQ8wOcAVNsQ+a9DukpW
pf8B15YTj83zZv3xRnXoDt3j0aVRCz+ibXxrA69siVKiPIojhv2j7igrMhfmnQOY
i762txzWuDg82V3ShahS7iR8dviCebX4cG0UnFoc6Mre4wMr5RY8AuhgM93ivLEg
JLvWEej2hXylN9jAiojYess6b2xHslczT4H6mgLH+sbk18QR/1BK0zSdCSxQnI5E
53lPFGQPah9Q/VCeQNd3c51e4PKAbsGjqKmBrohMbSE6XAKPuVKrjOLRZqX5A2Gc
esv3q0fqt9pNdy4k4CGKk4RQJTa1x9U1WAroMmrKv02FlfNuhrDnnYVFZu3GWCmQ
7Nf6iY9JpZZ6gFDcJg3909LA4oeVWPOQk9INWGJa29fm0gQLp6OWjTjYVLJ/926T
1P+oS4dGYr3sQnLA/LZFZ7Mgc7LRRAFYMDRX6HiEpJlRWNicwSHOn8/JI96SOQuK
8ceJx9S8rcomSHN63ah38L2ZEA5C2w6dtMs8R+KSELBXY1Yy76epmY7EjUgcx819
lKf4/mwvODA38R4B0L7hdgac2vi7ECldN6Zd2OpyZL3kQVLJ38eY86gNe1ANVvCY
kOO9Y/bJhvc84YdtgxASbioRs/mY1cT/DQzUef2W8gNdqLWkXJfrhSW8ugcJPiSx
Dd6Wz9GX5UisrIccNFRk2UZEL9WGB808knLyjXUm/rbOy+JBLbYuJiHi/qCYqqKw
0T5y03tZba2JIN6IWG3J68bume0/C8pxDnyrQWjQeK5ec/ZLFbpPh2nBFEEolm5U
bZ/uf6+2ut4v3y8yD9Uu0snnc68MajxKIMztcIAt5XuRrHImSuLLs4NCLqZDpgVR
ZvHX0Ru+oqWwOXDm+WsyCpYHUyKdvsB++t4CIKgmH7Nm/AgcjuPq5pDUIhtUBZ81
1itbRp7X4UaObmntWOBXkXBLsTH/ibOm3Gb50mhRYw5hDRJliHXTla5EdDk9CGoy
cbjRWAwj0zW3izkMYuFMWa96yUAg+dNpBzvtxZBOyjPki0mpQosYSCq62oaC/0do
z/qvK92mDUYIeG6WesftjJDLj5xi4TdVaoZRb73sJRKPLJONpMU7YLG3qsCamUQw
eNJgJ04UZsqYcM+dfY1Dvo8d+fMfjsuz8cu9WG5OIutvJes1JMAqw26p5yLLVVn+
ClrokN6u/tPXLyCSDXrjnaQfcZID1h60KbNcEgPnLotuK4ng0UeH8LjO+URxj7j7
gJ+MNiG6priDR8J+vsqy1Lnt+Wh+///Mg+h5UUOK9DmVMwqGwUCwzrFrpnDIu6MR
rl6mMdUNov+aTBbImGWVhxuJ8W58sSr/Gz4LehgB/teuS1oMQQTh8nA/yVqgRg+E
P3jszZqQZcxXJoR5ngmwhG+mNrcCpI8ArKkYImN/AxlX6XmLkoMDhN4tuafK7N9p
Epoes8/EfWV40ZXTQQOjQ1vWRzCib4inxKM6iBeHc8spV+TOKHhodjyn8/2R1dFR
GtsW9Tu0F7ks8re6ChTT/nT0KtsOwUn50OF7dzey5AZ6qxA4S+/W1cwSXJdp+UeX
KSpTV0LqZWAsV2SwreFe12j+qgR1o2YWlXLoSJJYagW4YKqrbePQtUHNgjSjWEoP
pNm36wpzOLH8QQ4w8u8PzltzIQtdpfZ6oGJ0jZ8ex5iAu17f8nD+7ug04kY8rBs/
Owv92RRylC3MkaagWnLqGhZSNgK1P5AM0uNih8gBRLkZux20unWIszW5FDCsNmLP
d2U97ZCI3F8YEncrEWH/yuIu6DqT7FahEm5z7DRE4G8Nk2HR4XiBES9xns+dyqbs
c7xGR6OXnKNgFYYezzVjlLQivW0BGJgVFT5bMoO7TWoyzKtl24Fo+srzx9BlLcxe
9UFosnCDvwpCUZgVQi19afpTjnWvks3JXBVjz7WIO63YZru+ZbBO59OhbwrAvK3w
Maj8Iq157jflrrTFRvAEypsl4TQ8mIGURp3+FIdJqlDA9TnjaDPkfLLCWrDhMv0h
tgEQLBxgjr5U4hH8FLJEtqShm9WToHVa/9NIXzas6yromY76TJ9jy9R5fvSbJU6U
CMzC4zGp7FTtqDC6Kh8LS3l6dA0/CbuaqqKJOQrTne8ut5S/TQ4/Gv9SoFT1EM1z
GAFWHgAYmiLYf8MzTKY0mG1zsUccWDwEM2S8f+Aa6vfBucYYMB63ZEWvI3DbERrG
ACc7dyW1td2nmWFkdVbgJbdQjVCbqy2zmv9HgpY2lHjCcn+3Iy3G2pWzwUEau311
+scNYQkcXU68/YLyT8rugTkPSiVBYCKuB3vOmt4WZUOomRIEMyFvFwRBcC3PUVua
LpiuTo64GyjEHhg3TKrG/G4396gAPkCJYnGTKE9mIfzU8Pe8PEgB6CyWKD8VbH/4
7rtz7/FGtj9AJz6Qm9g86rAYl4afnaqndp6vXriyDsyKIyXFkpFd2iqykM0sYrR3
2t3CXAfKsLyIgB9QzhggDDIdbPzKQf437KTeUUU2iSRODtBaC7KR3sFUWczwF1hK
991WX7abDv3t83PmY7GmbPhp+6eAc8FV2CR7Hz56uGGe4n9sCAAPeE7zlhMooAjE
oyrL4J2skz82VZzQZwRLFtDirFD5q/jfBh8UzqzgsbUW2UnlPSANyWzHYEl+Cwy3
6UsyaxugwuCnxdc0mfWqmV5Moie3HEbjNyCl66bhmvidQoTOEKuodki6kvFLol6Q
5b+e2qvC4JND3zrgYrf7/1DfGzzBj+EiV1TGPx1kLUzQ7P8xd+vKm3t/W4dqowGh
NkzCKMB8ldpHtOZ6TBGmmB8VXG5TsN9DtlfCAnyeS+FoRVAvJA5hLMictomVQn6k
luzgtE8M0pptKTr86QcDZKrEIqPMWOBZVttUXAAbdSNWKttsNu0kJ7Vt9By0lVFB
tvkXb/pP2IeO9dXf42/fRRBkPtaIT6Cam6rIOi/rSO+fM9qJDHQIFDEhkdFcfGaE
c1XWNr61Q88k4iy1ByRe0u3ZhByetE+SE3D+M7uwti+d9IjugJ9JZB6Tnd4e9eaL
863WVCINd/VrKWz5vXGcbifgFwdluFuFGGjePfrOFDni8V+QfoHZF6XG+rcxwqtl
S7mIgwZ3oRWlMJs7NkVMtitHGp8K+Vgt/1krURDGHCL/iMEEYh92/40cjYxoH3V3
kaSNf58aEfQ6JqVZeePCGX3ZhEK2iV2J0SVikAFjzBt8jOOiYuCRLF7qwPa/kWT1
Oe1PKNLYPGPJnmJftrk4tMEnqcMa75dR6NJepa34AZyA4DC5CKx+N0PaTsg0go5V
OdioBpWbHucmM+YZl2KSrQQHSDECEmeBrx5SSCl7q00VAWdNN9WNt/R/Fv5ZVhMm
bcP/uH+C4+HfaXLjRp4g/kCRrwIEkTMcK9chAItJtWvfKrZcS9G1fiDHmrcLSrSw
YZKlB5g6a+S8RWst0Bi4YO+gtqVl/a8d7ZSN5Cp6SDYOzLEvKe9OWSpJNW5MVaFO
uI2xmnkVu+JXogn5K8VmMQfMpWHory1fuzhK6sN1vEKmrDLEBZr1OxrRS12E7Wh3
YIOLgjstaFAN7ab6e4dmdyy8SG+VeEBwtTxWbW4NHd76wOrVcBSvFPB4NcykzpW0
f+ELj2E9/P1B5ULu21Mwf2vifqybbLfGcLfx1bAMlfiOS+whE3hcLkRPbBZMZEqx
56SUbWZqIH4xaUuwAflNs2KLevQlN80A7oFjz6kngTqc+ok183BZjtK/vgSB6xmG
CzEKoys0OoN3SeSSSBCU/veHkqh7a9hwFSFOEPlchhk6bkYHcS0VY1bO+FUSga/V
kIDTdhZxEzNa72UbQm3EJEA8+SfGXcMqmNDZZ2DTPN9Rhq5n7RcfFzgBL8SjYhgh
MvB5qYGlZyGRWujZ8o3id08QoBIXH4p0LHoiWjHxzhpskeYbt+fwQQ3ERkOjogxb
ZKxutUp1B7faxg1OYRd5v0tQJ1Tq7edPKaW1cU9/874voho+/K+Frou63ZjE81y2
nI1R8slYQJOrlbEmwU/SUZcuEo6N3+bO58uUfs8rHnJ3D0Z+InhU0CxzuA7vUq/x
DcfyhyE33pn0azAD3NQDGGVsF9J9yapN/5kXpuh404NxCq2dgqm8yF4TGpNkzqYS
P9MuxDBUsPxgv48+VzyANl5x69hn9ZsC/+dXbffQW3TuPRyOF0ZeI14IAgp7M/Mi
DgiN/TBU6qQdU4rDIosGFXl/q0PjJcl2TU8rohuCRoJriXBXQhRdJWLPHX59nD1E
m5favBvX19Uje8FxhHNqhJIYKb977LLKc45l0dzVM17VkPs68o7yTHzrCkIsvpkt
KB1izX87P8VHrTgsGh4buUkcYZGSMUifYJDbqLVzEVGPy4dy0WxSWv1K/PQKU5fi
Yac8GMrAGZUr3zNPhBxIpfY9jIM2HbUp4vv+BlEjpiOgPHicZ+F0ZyfVAgAO1FOE
lrpDO+Sph83cteh/DoPYLKZdrL+Mr/KdC1AatrA1O+c=
`protect END_PROTECTED
