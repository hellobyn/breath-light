`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BX0y3D8W/faTPJfCw3zrMOo3Nhn9a33W31dKb8YuAGyYWk8vikWTU67w13LoxIl
TO5izCBpDzSFkU/Vwjb22vfl/DOSAmp6V6okV6RHKTTSuuqZfd+Y9FvSB/lDfBTJ
D8eBRUyVUX5PQBd3EtGu9sBOphrljntAD9QktebJtyKQ8dUuo/hm2QlsgiRGcOVy
guS7mxGKACUtF8SdIq4Oi2pTCkHqsmC0as1ewfHNG+OgQ5kWo2rsWjDCHDBQYMYL
V4oMrsyagIG/CSjaXb5bMdx44QgLS44rSSkiUxU2TOBYxkoPtSLUeuXIs0k2Fh37
BXSrA/t7kN1QaYQ50Le+pAUXND6rzeGdgK/L060Zp2TV3dlD+rsZpL4bw3QaMsJ3
1uDEsusPooIqVMD4+vX1CbW9UOG3IUwbEhGtkMpC5sbuJiQpKyC2bEpE5gtN09Zb
6joP7nZQcB79bzIubd2PsCg/Ys89vceDVLd1gBVsPGPxLXnf4lePR9HUPJXbYCuU
rVToAQShFE2JJUPArSjxpyWn/MFMg7cdV689PmMwuz4nNfHgTxdcdled7Mywkncd
7V1p6dFFro3MhGkuUZPjZMtpwMd8M39YfDU7HJW6WdbktGQkRYaYyA+lTGSafoAF
YFiMfoue0LJPf34giYIGmNY9sZJ0Erkg7GP/0CLNoNc=
`protect END_PROTECTED
