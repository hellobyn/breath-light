`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMUpgfnxzY6RRj/nPSkTnH8PmhQMVmjV7mM5uwT1554Fm2S3Gtre5x55ajTYZliP
AdG/5vT/MJQxrys1v0FiJdjvDztCx9HdJfc3wjCdnjfLDZei82+QvSEKRAH0zrOk
HfMVa4557RImI5Dy5r3WIEbHU4rJMB1qYjp9eoYtZuK1axrBXtxJGSVHc9pvLgGe
Klq48hGhlq79PCPZQ9Hv0TXtJPkpPMZL1T9ia/wx95v9BHZZdVmdsRuvODZCvDtH
hlcyTvaAXlM17xDSgHzmZKtnTubcD3ggfDXJi+KtZo2uuW23LARGtd52QIF8X/uX
gtQfW2s+lCmxSmt2UDkz5wtKlfzuM2143CHG/HeonuBQvbvnKF6hUiAF9AvuYRVb
2zH/+tjYP80T58hO+I353yUTphfdi83cRy0/pI/IaSpjampey/TTKLGKfn68TDhB
+o5VwLkC7j9KyxjEUoivPMwn7xB04Y0qs76CLZXGqylXB5uefLKI7uA1xRTxiWS5
TwDJYEpQZZCI9g8Byf6nq4wvGH8YYkfpqq8jTbJUBFHjMzc+uqXQrY007Ecbisxj
oQWEoJIZ/H4e1LLrAnrFWZNljkZEOdPbrdk9NunUWL1UDNL8ZykNMsmvdKczPEQq
kyZRriRcJJJLVBccW7DBwXyv9xDlWrie8YrwKn5el1BlCcJdM1s3mOgdttI9Zoyi
6y1Xh+9LujUHRrgOwxckqswXCo+hXx0ESOe2sTFfxVLJDOqivLtLQLwbMidkS3JJ
viF3RPABUdJt1BoPEvj6e7J54K4a/THmKkiDVRYRVkg8R+cmWCg8Y3nhlcHuPX1V
2Hxrxei7SeMZOznfPFyt39sn43/WkD0mC8vfV0EQRSUBetWLE0TdGnitL4NUZohV
HJcphZzjBTfw2/E2JeUeTAwxeeybqYHu6LPJ9DAgUS7v08btbFOV5LfM7KZS6w9y
YuGIQ08VhOun5Ljq9KH7vxnOTHYf0exLUstX4PFtPJHRxdc0BqiJpnfYg2v12Mye
5uH1hiq3umq0JLeYmrU61SH/J0lhTiGN+FiTToEBRtcM+9ngUHrACKESJCu3i1je
xD5zFqg9JvaoLVQ5X7fyuoNsbUgejXXxPPViQisfvCxUgrN5YrMIZ+8vAd6d10Iu
7Cts4MlJKvyIyM+iyIsSk9zzkFJep1eLC1cWBkeqZIsbQkFY595e243Zw5D6SFFG
`protect END_PROTECTED
