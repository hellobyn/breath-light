`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4rGPaZvZhorBdqIUgMaxe0XyImu4RJtm5kRrjlUWpeWJoavXcF/aQG6v4UweEnM
YeyG/TNha1h25DbeVkU0DE9MMRI+YKNldsHHZrlXEEKXvu5RggqGaKklL6Xv1JiZ
QYc5AckmlxqqpDkMneoWNzzq5ThBfcSpRp/pTFmun7Y9unraU+u7FqauLgHsBG1A
Rb/h2ttZzXbtNWfhm0aqmNp//NTSzkgzCNRl+89MBtPT5BePLraPi2RGcZr+WEfA
LxDjhtmXeJX7jnCVz51grzof2obn3OoUdRnbtQ9g1V//dCzKcqZyTzJieanSP2C1
bCOBEQby49Iv2aXMyhRC0vTcto64i/GxyU4lmckhOLAV02bScz9mV2XRvuo9Ddce
8dFKufqCZ+2AM6lLHfsr5wek4pNYrjgUDsI5VxS2zptoMt2M7peof8smqgREuWEj
BbbweDwc3SYg7slOOYOMe3kgnx83u/p5Q0MUF7M9uXcNMbaXlRB8Gt+tJDBdTbeD
Tq9nlmmDyOwhkp076GBeQkcdGKGo7jCb672svMQifzHPUnpMtvf+TsTFnUjk51J+
uphvcOT19Esi8XSM3xUhYnrgyerVjBROh9fnzAAV7vAa2PdbEKg//hkGQxr5eLC3
3cXCqdqeajTSF3LGSeVFSAMsH6wTMG+gpaU4D5gi/Thwd1MIZJ6+987vWOPIZ6px
vttUjJlcrFUOpothwlnqcN4JRzlo8SKXi/6CZ5nSB3bTysNOaZubGzJSDsRskLMB
cmnqhwGSsSE9SzTp+PKSUsXNB7EpV6JmGUI0ofSE1R+utT0jlimHHEjqsaH7ncPG
L6aNqdSlDtCt7nIn4lTWQ0PK13iQUCY3f/7ftt1uItl/cphuE1zdt7u7GPunMZN8
sR1DpK9v+FlwlJWsziBXCBdetSYxz+vqNAXYK/sEy4O9WuaTbTdHQukjtlUT/WZQ
xDMnBAKyA+q82CSQwMD48FnwkLYBJBpI/MkeYX4ah4DWqCsmADVeTAZpaMoefQi1
bwtevpibm+MXDXjlsBo/cEtiJKiZwJWuxtZmei2mr73uVcgK5rlmTcXxkUqHY5e9
2uAtjM+2OwCi/oKhKCztl1IX3oVRact4aRuJTx90+kVHLJME+QHAkrV/GBuL09hr
fspH0S6eMEME8+2gsJiVn0tQIR3f87gqpLilNkkPqgBUokmr5fT2cCRv6w3LhbIq
v+2VqtTdHPbIscej9ya42TFopJmnPrvtl1perFHChReB664+UleXZGPnkHEuyRtv
ilK4vAweCv0LtAkcpEblMr7y8rv1G5U2VWH3ryoPRmI=
`protect END_PROTECTED
