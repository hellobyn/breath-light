`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKFrCzCBBGHjmC+owuHdE9EWu8YSGOH0nip0UQ6SXHf3oOZ0rzUMRsfh6KXtnJAT
+OlzJiIj3/I+dtb+KGYCmPRtWFTBeCwv6DhzmlRTEWL0dW845KMFt4aBhbpUczzS
NIvq/lqtgqbwSg3geBIO1CkGYRYeO5XHoym3i1uw73dJvkqrgvIpwVGAHCNU4v2Q
IlPMpP7TMM87b8mq6WjQHDGLAGpYIdg9CFaivjqkdPlqvtLqDup7lzGP8TMOPUzJ
6SV4tH+2TQBGEgyeY6vWqisQ7eDaMF6PEqnFYwHs/1F97v9UanEB1fHnCU/DtYZZ
IOdj6/GYbcE4SowV+hel51RQwob9nNbSkHdcf8yJuyR/ptKZEy7z/XEjmTBJBEy8
MZDPtozyqcdtdfAjYLnYrunYJDyLpUwApPipbXZtGWKRMeFwIsvIKnKMqnViIAaR
pco9i2Zvc53Yf3SFAkMzVr5EtEovG8fnhaUGFEPrXssVqo8nxJBwPqReD/F9o7ec
uQl2Fyeg1YJ0n0lZ+Ttul1uBYte4Xu5YRZa5J8vp1XUGMBRODEXbo2eJobdc812i
Isoi41CJfX37loXyG0g5JnyM780OCye7ldxf+9Mbe6iJVIMTSNcPKdwxmXC3XHZr
sBcpecAOBx1Bvzm/UCbNVk4rtXoJteT9t17iRbMihA9VnDgxibb2K7KMZN4rBbME
9yC9Mg6F/w0Q5Cz/C1E9hikB5nfrr62KqGff8BgM3bVpFWiToht3OGhUVLj32V1K
nBvxjL1cjKB3d2hUEh04vhBUkjsjVLolBSuTrChILp5DK0T0UiN0KAN1vUvhLLeR
ZzXN7SUtXxoBAMPfUafO0AfodGLaYRs9m1yob1xY8oYaVd6xJp1CEDHsJQRphG7O
rEDQxROoZ+P2lKWvPRIbXP2VXGxxrG51Cspx5BJAH1TCBy4wWRQkYwbiAf5eG5my
aTXQGq4pKtKxpi1Fa2DUiIh2wo/NrM2VPe7Swj3mZJsTk8nQr6Lig79mrLwMMtQb
PmpLzI3nxkXUEcp8gO/8eyhzPRCr6fKFkIaR/dPF2YRfQcI8CWROEjrYoaMZdbX+
x4u5LvmYpxjoRWsMJWwCfqc1niUjVLt6SqDg4POLV76sc2MNgXF7eJWy/Y8F5iRK
Y+GGEMROxWfjaVOpGiK0RwLxZVJYLCCuhmtKl6ZVIr4GTvYlx7I+7+x/DINjk4St
MK5zffj+byG/pb9fjlEMZij6kOadG5puaXQng04e3afWOaLtWTizKiacqieXv2HV
ntcoistBYUxiDEf5ohGVmIygqCPKJOlnCsNSi9aUSq0a+cC8PmGupvNcWMRFiWQj
gXneAxwsbYBfHoyWu2DC9Fs6N3h935brPQuWZiG/TVTExNf6cdLPmbpjQqO3gFzI
1YwysfHfdyWJx/IRoNFzMQ==
`protect END_PROTECTED
