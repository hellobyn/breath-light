`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4X1JqfDkVbRJPSwd22r2XUcJads+H03F9Hi0OsejU+9sbX7MSgPodOD5UjgRaJaM
P3b2umXpPEbyo9vKBqw0G13Sismex5MZQ0wuMsvozg6KCdyvsKpOFGye/N2gdECU
bflXsOKAcT67dXjfmQs83DkwuCs96TYfzuz9a/t86bFaySjt6FNoIhhKNpRCBcNb
tctsLq87k2UHSH6pTvYy/4cfGpZa+8E0INFtAJwhttb6BMcUuxcIUzkdoy2A61+u
w9Wot/Ni8cPUt9lsWANyB96xLMZk5gwSMukQ9zYz+kWEW3WhJda+1RpUE/H2Pzcb
Ep8WJJ0lJoxA4MGkkNBiqDqByrKVAq3WBWGGgO+hrSUOav5S41FThjMetB/VWdzm
BPpl5RTV16GCpRB4B3gGcK6wo8wdm/5i11fwy/DULd4MUY7qdD7htGCpgRhvMXFF
m7AS8t+Nuna69p8hW1I+FC5OWcQkox5IewPrzWxVK/02TTa4qXh090YcMgGgTwZd
l1mCNjEAF6XDcyUyhU9oVGbq15gyJ+3eD9rIoFv6NriLLZZYe5Z5CWNjGuG73dKU
YdAhQN25w/IADXT6aIOtmurHJqZeWp7JpNE3QTcPyd3cpnY6yyUzGSsMBywzcPg3
jf6JjBMlAiKAD8mOQnI94+Ng1mS6LsZPduLiwMv5hB2rR6l1leSYxUZY3/ihr3jr
SrQrfsEvP0MxPE6TBg++CAOKtCVprAFmbNMcdnR2qOgZXNO676jIEQY8B9WYLnTk
yRFWTl7bUfm2QZp06M+hH3pzs1p/LElEc4J0NYhYE4hMT3NrKJpaitws7MKr95QA
CxhYuZp9dznYtjjV1AfupA==
`protect END_PROTECTED
