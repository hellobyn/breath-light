`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8V7QW5EMGt+UTD2NvvpaQKgoaZMtSfoQMFnxeUeOtvY/h60w72T4a94rSEv/apG
n9B1ulRqx3MBa0QSkUidIoMSyuXskDn75UKlZ32UGncc0VfPKN/9I8LYCJuivsNz
0Wq8DsfwYXXEA6H1VK+UY2CiSm7NMfTqwsrwJa7ixEb1Oj1fSwH76t+6wqWRFImV
whYOMKwQCojV709GjMYIkKlc1s9fEHzk3jxsH25wW2kFfEZbcSXJnjVipifUev3c
BcxaBbm4necDe3hsrc3o3R+MZV6j8P1VRlkttw60Bu8DDxnUGAFx+yDz79TtNitg
zxKvhDdlzKhc2h0h+7AWB4cnQg9R9YdLx8E+cz9XKV8b7taj7Y+300AK54uO2oi8
ELxU6znmW7NcZJZXN/2oNgQXr4L388m6rz/ixgGWnHoHuCAu7WvtSImKgEFFGFgT
gKaJOWYYccrGrA3cpKwND26GLMsOOFOt4Z8I+0k/GdEeoeoL28X8HgIPoOFVCLYP
fbirk2KLsHH1F+lIRFDaexpxCzASieS2HKFBKb2RWvMmzg6RQ8vBeje05flav3Ko
CpkVayrHcTGmJAZwORML6U1vSxZPsQrFuJNBVVP9Co3yVt4tTJXlHCceXUVMYY9n
dX90m2upMf/asDTheEuDP0Y3UwjOrf3iwLgSc4t7P4jvK7TyxNrt0Su9auT3y2tT
NtYUkAclZYPFKelKgbPImB5yFyXYbfZ0RI2RSqQKws5g86cHecav5zJWN1fzkUBn
oWgj7Z/KR8pMQiWLuqlkbIje0fYGfLDMwB4D1z6MKVTb//YF+HoUNF2jHItHBSZk
VWnw1HkVevQYYPAuZuBKkEDVxy1aOkVM43w5LcB1lH2+IWmMWFh4izx8AHkCCrqm
f0g1f6wjgBRUJOPaiVEKG8awfPz+Nn+u4YbQ4ElFWfBesmWUqIRGOs3VMVVJGF0u
4dffQkQhhyyppLtsfCGj8MvnSpsHNjeg/wqY49OsULunO9AyArImQctTzaSyPgUW
ZNT2WqKSOn7V2Jc9Wr3TzShr/WtV2bFII08NiAAUAtLIWiLgwn0VUNQjU5ujVlMJ
nzPrK6nEGKsH2kPzkz9bVwVGpfFEHeagOvEeioxPik6fXQ04F/8P+G5GQvzU/vLj
ZmNyHGR1xr1EVjOS2X4fO1HD50NvQ0JlKEQVj8Q44f3HL3bbCXU3ZwW+Grj53A9/
dJDFFGhiiaqNk7+giF4p3Zzg6028AyEIQTSzmC+if7IH1GCGkkk/0Mts9KUJYUvb
eBo6ubQs8ICjWCQOCtqIFD4d0xEhnwU9oaSGnD1NWciW0FU5aqmOF4Y8p6qQUhBr
63U8WRqTMN3rF4MAfdVIoHQwRrOAsSgZesypC9gh++DTyIZwbEJQIrMlcTLNFVxV
fbVs9VdFKCDkpriUXsyDxau3m8S4omcsuAhp4AG2SAsAN9kuAiplyvbXSoJoHYGV
siiKRg+BmmSgI73fIBQ1Sjbn+nSWbRVEQPdlLhKyu3Apy2st9lhkXoCHMxa6JWGI
wAJ0BfXvxhiFptyRTDVjGuWEzUjMiWs+W8D+J16diM/ORmN3Rigz8tKmpfgASXG6
2il5zGv07AOyM+h/GOWSnv7v2oASHJTT+ONEdVradKE3HzQKGfpFHCcikX2dbzBf
AUaok9fbffqtBYKIgjAGiQNQO62DaINOl5HZifruAVbT8RvFFAVer0zc5WhHoJE7
Qvn6ml0dOK/YsKtZW6cJlaPI9aE/6xJF//NtNnb9xsYmwE83r6l4w/CnQv7uFA/x
jtJPGLdNRP4BfDuWA+i7KcuvgceZmugr5ndnmPqXz3im7RJEMBtPplyuyTXxRpyD
Q4gB33tMDqXsb2Za3xv4CV1OfTur6Dm8RaACoA3ytAJS6Q8jk58l9txXBWpn/4mb
HwFXtAIAVJ5vHRhvC3AidRRbR6P2OdlXxjWr91cZAGH0KMQjV/i6DhyzJy4v7UUg
JqpWAhH/voHwJDzklBCz2EVUaCQqesk543avkaW7kA0j4e3yz9BQNusISqNcEWwD
NCpcJoBjMmgpnBfNW2zLrryncoqYT32XoMcD0gUMl3odpIlTuKJyM6La/OcoM2zK
73ruYdITMVmEaX88ob1s60S+flr2Cw8jEjEHCTrds/BIZPjsT7IH8VG0h86+stky
mlmkNOdbvrLHkbvgxteb5EqrwZ8/1Snv2YH7hp1M7yj8xG5r7ygES45X968rEFEx
z+FVWcVXebqPKiiQthegCwk38xOssMvM4g1NcgFAY1a96Lt/SnYiLj906AmSsl1B
nVIIAnjLOBnZ/D9Dm32sxtx8hBvyyYAYUWEOgdwuqq4Ne1sakcOouYk8vwlsW3J+
VRLJTlFAccPfKuqLCysLy0oXAAkRxt1WhcJt342ae4kvdaCqBVvvdyHlH1oKoKu/
LC8NmGNnkKSPZnA4XyyDM+l+qY8iNaG+T6EeoLCVQxlVmlUSSzFP0MTaqr0KdV0M
gUi9mZAx2IQIRzaeTK6ATwMlbSsG6TUjZ4aaivlKPCiqW8OIxSirTPCdaFbEnhT3
zUup0i0xivdjI7vWbMlCUwMd+HuA2htwFgm0l1uQ/0bkpffUsB+JKazKKHadQKtf
aAvaooTNF7dWBO27gabR8A==
`protect END_PROTECTED
