`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W4wDvtiMhL1dJsleKRA/ph/TlXD6b1Gid/NWPPsd6MpAwzM1el3y/rvwoCBb3pmA
QFZgFAphROP7a9np3tS182ft2mB4PV4XAncSgznbWR4j2rox5xeU34xhNplWIzPT
fdAOpHsIC0nPXBVodpfyIjMKeX/i6BppCTWKPOmAanw4J4rL++vBZLHKGmaC0vd+
2bpnI0PwVfPxfcrtE4JhmPkY8h/p8gpcmJFe/ePysVG8t4un7OBZq8jzxWhSq+Di
hwpeN100u6xNNjGzGGrCuzwvSN+XlGoeKZymIngN/fkyDFjmHIEit8AkLrfeWO81
B9LOx+DO7skBJjDR8VeZHgt6q/qKCErk9HTPTBC+AYuel8LNgSxMOH8DTxbf4YlT
ZUnaOY+HaqYgmjbT8/OM8yyhNbZkpDd3vc8Z2SZvjal6x2A2NhoLJT0cIXvbQw1D
Uvt4knyRgU8Yh17omzhCM4lSnOKK+HdEaGlWHr3aFj7dCmErOiIninMQWh+nC6q2
Dh2tQFviO4ZTGVqmxZLgeoUNjTh9InDCtzBtoXj0oUCoesY5lwc2a92n4xM3FPXn
K9Qo/DMbhCyuz3NoD4mBC2xQEL64iP6cvYAAvfEkALiv0pTMGkBjN1rmS4iiuNfx
3JV9lQk/IgZgtp68fWGemSmOD5SVG6USvq/jSrQiAWZFOIEGHRyqJlqoUCcT+G4Q
icQ2gr3fDebVgHfHIVlSPG/vURFWxRyyCUFVJ2TsMFIHqiFhqO1CKQ5cQfWlx5Q9
xgO4JMf0V2oUS4XWmEnaaSKQwsFBbCldlki7lkr/EO6akFMcYuBJ1AyxNY9taTOs
HaDo7+cxv+adLVNFbuXjYNTmA1YHVY4t4MVXMTqZJHsW3brpevr74+lBZhdsi3gw
Ue3kUYwQDN5UJscHbUIiwQsR/XimS9VAxHQtzonour1YPlJ6XYrJaRofzsZaaXYp
Ae2LovXkN8b2b8hzo73vr4ns2YRfwRUvjKzLFMEGLvusotWcnIuI4b2QCBb65HDs
YoyssqVEIr0lBp5hHvAl33berT1PCdtla3cpj5xDzTUHihzzRxMF21NIGprQ6eE/
m95q+X3EheamlqgUhB8tNtGgYMFWupoZzt9tUKM/pFB3lgqPUKZ4AKJpZDANLGez
yaRzRDhCcO466EdZmzxCEbmahaFglqrScYubogt/HnzFOXJrqQYmbS/u7VfR+ABN
mr7FNZchmWCFvXxNwqXORjjndYxk+tPmXkvFyRI82EVaM6dPRabiblyxWn2ZYnCt
WpKFealO3zmcaQKMux2oNN8dP2n1iHMsAKWOjjzyA1WO4abA72aaUTrYW2Y5BHrK
nzKehLZw+RfJjbv/Pi4TUm78IL/DqnQjODhTi40Jo8t7ArwDPYnWDt++zfUfg8vR
kwtzklPqf8QFPyWo228oOc22zdeu4gQWeVV4ZIpGXQYPzX0cMnkqw6DkDEyLHNls
fZIB6qwsGlo0oQ6/MoYbnd1H/+rBL+l23sodF/0ILAXk0B09Y1OvUpgagcDgDBrT
jydi5b1sBvb3Ms+Yu222M6qfO97NZb5bIr1mbjBszNHvnNPEXZeSK6gSYE3kB9NF
3ohOiiBK3Ek57GUEzxmrns6muEXtO3+NZOFvKfYRx9/6Zv8+yL2hhsE8UMfC3+vB
t22MkdEf8P5icAmUv9CpJ6emSrfQ8PBzCQ+JST7qpp8lsuucUSQZJr5ty+6Ww8UY
Z7HJW7AGfT1vr+LA4oBFlqA4eDcK19SSk70ey8J9XtxeKyElyYnWVNF5I0LbmQOe
iFdwDyaNz/82UtVlswFlTyy1i9zkBnR10uJXOP57cUscEjq0+QaNtthKLVhnnugR
/bneG+yYW4lqXfQuGHIwAKc9qv+UXUBKhEuDhiRShPMxxwVwu72HM711UlWhyXFc
h/ZAVnB+CoKZh6PIi1FEsm4ZHdO3dD/L7sKOUDUxcopjZpYmNd6HrqMv+0EmMBL4
8T0BeE+Yqnl2rHM/DR5+2hIOKRX1L+JUCc0I8coNe3uYrNaY4nrzZqQMmfxJ4h7f
WxEPlixzrK0ORWs6yIdh6aZoQxhbrkFBH+MLlRAtNMqEc501byyfiBw81fSPL1Ou
s6lRQuD/ZWP1HSrDtX6XFxs6OZM3ialiAY7heebeuEgfEWW+xf91g938GoNXZtjv
7fznysklsLOrPwBmhTmQvX++j/peks3mEpc9zIEulCeNOZ6AS+UnEl7yonumFFXf
kkQykVb56Ju+Vada5/Odey+zJY+Kt7oypE7SpykFZXJB0tzuioG8soQHVQ2YIYGM
N3x+V2W9aIlnFUI/Izj+55ub1i/bhasgzlhQyztLhWz+VhWfi4nKHPQwHvBE3syK
sho5fIWZOtVPBONjpe3Of2il0ECxSMjqis2wmUhS0ITUft1KIFV+RLJisv5zfDdX
wX6j/tbtjPwAe0NtekWOBu8fVUfZEaKKgC663zru07n5RFnUEBFHng7g6yghKYya
Eied6RTQaCDVA9hqZFlXQFHkZwJ99DCiQGoVIDrs1UQGDUicc770nAT/d7HX0hYt
om9f0YftSx4EmMHO3U4u3MwDmGs/A24Ve83lVt9yODPJDHrj3YYJThWIYeO24PNk
yxXIp8nsyc8TQTWnV7qn3lkaHOcnDvlKrVDEixQzbsFmOVU3s2OkNANSy/Q5kRN9
PdSjZeREunjKozLXBZ1EUORPl9btcfPKfDj71Jl3MxNIgZ5nQfGQYwb7WOkpAD7I
HP+6UZJEXsLP/IqG8pSAyMTreNWFKjnGOSrG0azx3GwEsfzCFU9rYNpBj6kNB1uG
+2UUFuiNHovKlpEjtfrEjcf2ifIhxxelJEdUHBoiEpGUS8gXn4xKx66vBCmP8Wp/
3HqbZ4X37iLXQ0+530MaTH+AMIxPVou7/9/Lqr3ql7S4m0199rPtwwK3ZwiQV0M6
a2Cn86El+kyAarpTN6Th2r9rVLk9SfJlYn3kyCA9xGEs3aj0piYVOeQ8t7Q7Yp/M
HCIpQzzFU5l3Uu6kQFagvsQuBGruQI3m5/bop6SmXtHBUYnuBLU1XTwOqsYqiCuJ
XhmuEMVeq+RdJ9K9ZmCN4t+nFrTPjgy70geNknQe8qPqre8uDL/kjrVNgqCD+suE
kqi7vW6SaKvU34Z2E7JOoDqJB8+zSppXH4QKTiLTeiagnLAF9aVT/tjIygdEhnlY
vwlHJs1gaV899PxPnIxqhy5SpiQZmzRVxYOplJgq5Ou4uHZvGzAZz4M33rbiuKCj
1ANMiMuLydHeHRENXjKsxv03EMkNdgqeQ7fVQWKztOAGsU5aYqwTHKC4uehVK64e
mUz68Tc3k8nr16EAQ81PfEHrpdw3g3sXxvx9H/zUGcYOPPKKFDku/gl18MiaWV7e
1iv4QX9VtIdNDVntVDjT1Frs+iNqh8mktCp/PY/FJa8UrGH6hk0zui+JAZ/iIN+N
pzuim/Nq2N4g1m5+9/vGNh9ff6expff0IcdMqoLPPzMzz1vu9gjHNK4lQ0OhkmsT
I0sDVRoVR/bj0iLwCPnTggQwWA9YSgGuN+1ms2OHNQ5xrHPHYQX//mdSd3mJ9y/v
t8/In/I4UD8ou5UvdauZi6nfvTyImQHIKhoRMF4GgMl8PYeH4vRNkd80dm8bvP+K
sh+y+M1BS1QLaeaFo3jyHH+zK8jiMPE6n4itIPr52q0MNWsots40MV0367P076F5
eOir4dIgR7f5v5ffkiOLWSgIwpsl+7+7gVzVlbvCZDMpdV2nCa/5vNIxDCxdG98Y
zlweBf+GJrCErIlLMYIULxIxSvMf/oFpTwF9pDy3XToQdhVbYOWEQCWDq5Pdqv98
PgG39CgkTnqbLwlnWPJGQgtQ7sIqnrTuGNC9YqUrshQuyiRjKPpXn2OAXz4uD5YN
WETnZq7o8Emi/J2SfG0ErnkZHN47q6xSTjRQIy68xvFleEZX+02rRAnbBtj7ZiBI
zF7xsq4NkKUFduvxTHyrLQuEgP0tvYY5PUWwRidt+BGEtbLSJrbP8ndy0YxUkWDI
yBz0H+Je1CC/SKDWdkMIGUuBQ3E4XAx1W4e4K8/E4b1Cn2EGJOr88x1ToYP7cOL3
RYpe7Ozhy3We4yr5jGeW/k+2ekdKf43YF+BFyQJg635yV0pEg9rEqbk15bHuGE0F
4pnNqEfSULoNPydSRwsbIW0qYgp+8OOrVCiHBHXJ+LwaKzNrihS1dAtL0kv6xh8t
Ic78MAwiLRUbSG2Z3MRMWKGRxsaAAw5xVUbV/7ShqZkQsvplnVsYLoSTX5mMjQgO
06U41W4mowlz77DioJcMnd/dmvtVfTnre8dqfNpSUyF+EF8Xk+2S0FHnqjWPcJqM
+ckv9yBmUJGz3xQ7QKKbq5yzLbhQiJAR9xC6kz2/wStAfc1PvbKYYPDAPi9OzCYP
4iT2wwzA6CTPzyJVcEH6u30EA0fIxm/pzyrv/plYo22qid/bp4W/k85cQAs+ruiZ
ijiNBJ7by6nRUorMh5wOJksWPkYHIegYdk37Tf+6nqeMeK7zT9uY+SKoYiWy9WVN
eHqP7az8XLXcTeWQXx8kUsFPUvfSo8+u2ME2QqCNeWGyIwUzcyzO+LE3Cn9DkdQI
SBDV4D5fs5ioq/kfOls/inyGfuhYm/b31eHcZRhTwj+D9MVFx9Nqke1UDrYt+32s
UAkeqEG9EHncL7qpEerfq3pHFJol5y2X/QrJGnuGqk5qR2JD4+EE6QAeslLwcdLU
X2PVMeLSroLmplH8FJml74XfEDwMbor4eLpGpFNB6ff+WOnnAEaECxh2Mjvvf4NO
a/0pbk72mq+08ycmrZl1vOdRZdo2YVVJdBe0mZ6Dh8FvXwvF5yX0ej2iJUq8DMeN
Ng6B6XVGSy8kpa5vR3gvcFpeVKFyw4vkLJviA+mzoocanLLE2dvapa9FMxheFs7e
W0SH1UtgnE12GeEjkRKEWBSZkLiDRU4A/bBrUV4XykQ5cX8dFbl02C+rt0+90+9e
TZNaOebGKYsAFucCF76RSseRall90s9wMpzjYjKIVVjbCRbVlwyRTAMAPN93KmhY
BUdoIPTzAbwUIzvLIOBAwkyvOc1+WxLNfOuBjExPrqedfupzlPsgFNGnk3Pu6dU0
PrkQNjeP5L0PYZXZ0t2ZwdoiZnq4EO+6GXOOkcAFz8Edsl+p9U/r4Yo6LoE/69zA
EPEUS7/N/Dy4Nh+ykgdEIJy1p8rKks9pZmRNY/rZIu8WiRwa83O7zNE2cc1jXQ2o
ND1bp7FVQ2lW3mjvHRrRbOInK0qzxgOfafNu+TqDVn+4dzluhyzObb34KFfrxVmQ
te9eERzLfaMfSABaG56E9AfONAg4f5nLp8pVe4/M5PniZ+176d9zpyR94RDeVYdq
8NKBFG53vH/7ynfNTtM9GEgc5jVDPXhJX4exoGZPYJJufb1CNBYzTSvOWvTwe+eS
MNuwT0TFnIFuf9HEsIewNIneurys85DgXETnvMVEF2VSE4ByMLtMBKJOKmUb3mw/
B15OQa8ZIHIoFpW9eFtSLzzfr8Y6A5gktCWD5N+anS+MlLEsQM67HMXggDKmfD3u
183O26DawGTovMybXmmTKqGjXw3A2xxeLhMLDLoPNthfhaXbW/r8qfw9/3QQavOa
auHfP6CvSkvRjFTDJl6W3JJd9gDOovLOVBkt0E1/bd0RmvR3/sA32HMyNf7Sw5X6
Ks0vErNbOvbjAP6BZZDY2FG7xk7jB3KE3iFIaWvgZ3vpeIUJxfotuY8sFQ9k5Gg+
C25FDFJr9EMPb0SN1yQtDtvARS94bNfT+JKrbAg+SK+V0y2y2YYTUxkpZxSA1klE
CxpjBIOOG4w8ZjTjy0wk5aWkvkVyxyzsZbHshqOLT//FRHmSIMfGX7NqWiqvfk6Q
f2v4LMyybqobUeWuVB7k7TyTxdqddi1+P2eL76h2+hnLDBAYp0viuY2GuY7fJgvj
tmdTTjWXr/+lTic/oaymBvxq3HuBdHphFX3KnMDmWb2GsqVgI92XzCYFeLfOJe3p
ta5Q/coTF1semJRTdD9WyenE2qnd6Cas+/g+aeaEIoMpEW0bJgaHhDg4HJMj/uHG
Nm50blDPi4kr9C33m3Rxra+iInNpUOwxN+qfX0nbAhVJl+SdpUR9um4G0X83YHyt
db6dP7MhnY/92Lg0g/vMJQXhNeFbVCK1ETqhzC4RSJXXmMMyd43Zd0LumM6kN8Il
b1+GmJ1IQ8ExINDrux+pXblwqkOSAcSf/OYgCuMmvhMeBtck8G6EibqzRH3VJBpk
7Ap333299NURIqjl80AieqiFVcovGk0OPGcQKkpTQM/QTSyGU+EO66MF+31ZROoD
da3RkYhlUY8G0DoNmPwQn+ZV1XTh8KSVS/CuXLriQWU2w5W+RMMD65lrB0iflP6h
RxQeL5sbzEwjJ/WQGl3jMbPXTjwK32CAfwFpkqVvcILeXZQyzcl3UnJZK//lM6oV
xXRZfF0ep3TAKtA7sPqP1UXRMZfCR45WEe0h5IrpBN9YKa7bEH/aZQYCTaS+6qwT
VI2e1qv5u6cqbsYO2BbqlLg8GWanfkW2v/m5BgN+tm0aYwRP8mhbv/Pjsv1pIWml
jnuf73zN3QYKQoFmE90kuVA0i7i9KeLtaDTHG5cbgEnguNsKa6c+nc6ONM4gXCF3
CGVIEMuNI9q1T7tjLtEXztitv+GNSRBDzmt3zAYNYQevITGDq8cWxtbuFRqi2vVQ
9X4Rk0mqSoIgv/lWj/4TgT69GaZ1+NCFUrGUxdWZn9QxsSHIbWcgFDdbl/zwKURu
bMfnOM+ZIDk2Z/X0DGzqXMUSxjWJeP5gj2zBerqA/ehNmNeJzI9x11TN236NlST7
jhn9hpdyRyC+4QHFdXvkL7ACzw1N2t+pK5kXmhMLphK0V+cvKic8klrPzNVFABSy
KMcoK8CUN3x5RiHX0RueI6vw/QhfXYOLq2xiPzxVEjELmmZgQAJ9XcA3UYpatl9O
w2ZdFqawVl+R3lhurieHhiD3uz5sNDvYwTVCcTLeHRPGLDpQ8jIKuGPBZs/I/kJu
vSccwgPN0Q9ku7gZ4C7zJZ64XWf24bS//dOSqV3NIjvkntO2P9HSuHJMnYHgczKK
ACn0jb9CYByIABoiQlMmmStq4D47HitJevlq/wkUx+hDwF5dsQ2fWsZXo5cLLDtW
T2DsEWUebywctjaag+SFKFGlSxSwxSOxa/mR2jFnv7u4KuMJEPVsWp0XaB/Imxoe
DurfooSJYWUF6gnVElxt/zNPqB2f8mEQyThdx51upkjjmBXKtkBSC97XD9obKTEP
jaXWJ83Go2DMGWcN3zo2vYkYUoB2vjjQCfFZevBNsM3dbWocJx6B9OBMn4G+wFv+
GfgoEjlGyBi74iVnzKymdLMi4oJhcaT5vUP7nX8txXCxE3hPs6X76KylvPk5bsAm
jL8HQqXzLUJ3Xt5fh0jjLyCqmqMN3iYO2VTWs8FWKMXec+A6oyIZkjTM9JBgZlsr
DT643RA+imFi7kPak/H0scCNLmWsmJeQd3iHIrU44m7qbnnuQuu4xj8yXYtwWlu6
NGlBUoHIL4SGkTOtHYOcPzw/MJsbLwKuexF2bC6e8sHfp2Oe8zlgk0x10X8z7QzL
1f2uGujrpY+dlC4sPLBiVDbBGIeCbNK1fx+wHp9n7tN71j+bLKewaLbW6IcDkWcr
4oZ1lMPHvzrO7eeRxq1Cfo6USbRpfguZTs26/YvWpDx//yZ7ojfhrHITy1Ytm7Rz
MD1jzBDCgCuBvlB18MysB7G2Hh7R+UvXLOQyJVm2Dg/5tPHTi8baxf5dMP9tUqcQ
t+SesWKtlOpTfDRWT5qXoVdLgRxvXu4DJA+8tJ3M1VMD2Ge3p9GSTMysnwROOI8y
Gm3uLaTKmxYLSS63JCDnqr7gzhlsPdBbBWt6gGYuJPixrRQOz4siniPIwSiEWpRN
w5E7r9DessYgriSEhYxI2w==
`protect END_PROTECTED
