`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVdLk/wtnvCqhWDls74qdTa+dL0EUrTJUnXXzxvBRB1s/aET8X95r7IwxotXE/En
jqWlLL4SRn79e7W81G/YuMRNssj68LmydYYZRto4fvR9EmYJhg+pawcP0u0dFIAh
LQ0fYkSDBCPd5aHt89opfJWql9vZQ24OpTXobDTZ6nsmD96JVTPCm/5jN30af0TS
edxE0jQpx9Ujl2V9nEzLHsImSUBcfAAqz7lIuYyZ18M0UjgjKEcwWJQvX/Hytf45
Y7n7binwePnE4hGruBs2TC2/aRax24Yl/WmG5cTN3WkEO6YEpJhw4G79wOPiJKnI
bN96pSWarW1te63j4JJOzebvI7i0yRBfzCawkZv/b4/kaD0gT7OhWJXvFmAf5Zrl
argCc8F+d6hz87Xd2nmBrZJOti2Fs/Yzh4Y/KuT2Q/Vq7XswR+HLogQSUt5A2fSU
HVvno+n4TOt5lVYlupIudO5j1x23/yZzzZtqENyQ3n7DHnLo/WUt+SVGvbydHLZ8
4MOg5kMlBB3iHh72wJPGY6RiVZk7Vw6h6vzzYGIYIXaAi7iQk4XIBNK2aSje0CVz
/1foiIdhw68KgYuUBCHymJgCF3g2q7SriCZAe4QP5b16fbVGw0hnzra2ehPVL17S
1bOO+b3u5rW5MFWNsjZC+aodcQ31cO17kmqYW87u5na/APKGHyF+Qjag98V6JcCe
KMi9UK+gKW5oNtPw8ZxnAo6T+cePI0Tymmg9x/Sm1QRee6OvZja7R5XpInmkFLUR
uHffXClYi0qsWVPerQ0TeHLij2OeoKPNLXqRmqq3w9E=
`protect END_PROTECTED
