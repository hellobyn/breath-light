`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8T4RRGFiKemtIEWb66T6mNu4JRAx4Ce13MTYAzzhxKqj1SuvKvtAxCXIJSzfxzSG
gqE9OYKMbMimUlAyr6YikhiTRcFAJYZerMPbF7GAQn7s2a3qDbN0BTeywF68UxXx
UPmdI2vMHR1Web8hzFIJx1BLR7vJL6Xl94iZypeKoobkStUNXHjpek4132CEsEpG
ZtfeSbmGuGlQPHwIOnzkR2T7Nczd+qEVv9shPJWstE6wSgerwh0PmVo/yC5UDhtn
OTuXPeRWoemRKxfQE2ablB83U7r7ZTiqeyFp2a+yhvkbIxXfe9FUn30fODTiJ5rN
4fGPOMgg1xNTvfcKbf3Kt+E1tJo3b5jnUFwMATYMDB7JvjuitFTlpVXKZImDkzDj
QhsAGWJ15KKdwGBGojLAVArayicWKCUe3NtvI09QRvYhRNlySIpzINjaElViABVI
1g2ZNmxNrqNajn1Bo+1/o3aCMbLE0uPPw/L02F6FIZbmnvu0zjxMogzqMdGvm7/7
Mjg9qHNuToy5R84UD+N0RSHssPEPr2ZmR74n2+T08yPFdWcfjiAvVf8kU9KA+eeQ
pQoGC4dSkz6qKYQjVr/RVEhuPu3ehXtv52bn2D8mfH4=
`protect END_PROTECTED
