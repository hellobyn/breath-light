`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRvStYqu7wT0bpGbe64Cc3k5rtmsMgilfrYF+S8UbzAVNkmoLeQkbi4goM1zFiwO
z4hc+e9bInb0DvUEL+kWC2qn6xDWLmpGTPE5u7DoH3x72/Lzdv2NgrMLjnftNIWP
ivTTQVX1VmnU8RuS8KQuO6JEGjz5NORu5+3CvyvXqP4B50wEkJ1tUhIXbyLnP0PS
h65Bn9uomsTjQz6Iglv24yw7U+QKAXuASMIJ/BUpnUEbW5sOxoFlcLcPuVHuyXas
57y4ibAg5Fn0zZ4tSnP1sP8jTb88UKYSzodwQPvDy5gY4Ozy7Dnw4PcbqKygmKA+
j4ih+JL6Mt4YUS5XVQAvFbgAdI/xBufffdvCZTA2Dn/IMXfpcTk81wxmyRPjIVBu
sj3yTDi1UAp3O/bOFXGAFQfpgsb75xnuXorxqi0IK3xv3pmhopB03oQ63yL3/8pg
2RVmMNnxvXIzfp+87erLGBJ6bWOpPuMXc0WEyY+upPWnagf3jCJFJIECCsX1kuDb
F30zNGfvIV+RkoOjQSYm6mKCllmHrgdi0MuTovig+Lo2BWFnP/Z33oXxDWRWeqVz
5kuBfQ3PcmUEo50s/7NLu3Gn2vkYHPgkEKPGlQSUNZNOadMNRAzu6br0DgOVa/Hq
5g1KBB8UG5NDy9FqUM//xBLJ/qOnOiLgzJz3CprNmrhMoENcCmenO6nhItI2BA2b
g+rLDI+RCwttzEtacirvBFbbszE0ZPKvnxT1dxYaU7RiIyFg+Ss4RpakQjyR0xG4
WclOs9dj+5uV7JA8vTyEbE/8eHDSvePIVcAr3hnU86vbgYjL8uk0RzSrDvalTEmn
eyVp0ccAWJcUml3gvmzMH7kdpsJDJkioZAD5sHX7IYrO7AFocoMMLqnHzbw3WNkG
iCD6rnkka/DIFHhXXe65gvaSx8jgDSlaRv1C79GPtZn3X26/9gyo5gzr3NZNAwge
rAincZ0FB2LOS4kh99sJglB5dKJ/GrWZsjUdJh+w65tZmzrjgjt96gLQkmcJgXAH
DuBwg1n6z4cmBPZYuPsQvDHcBhdq1cJql2JNRy2qEWLwaxCQOwNeKDCKTdXCmB0s
Vb5hJLQYvkl7iUOXHfNHl2LcgwQOXEsD+xSZc+UxAs/otjd3IQHjBKq+fd22W+iN
DEK2hvPmXivQ0Z/NTugegj8WzM1Vgn3L/4vSbdycw061fxAycjzQ1bq7ajtV57Dx
7S8QiXakTz5q3l7VssH9Z7YAwwwHVLEf6OwqRYUcLCAn6L/MXtLewK8N+fWFCmT4
7fXKMT5R2MJnD0RB47eD4iyd7HayQ1b4uYBt65uEdQP9JlVEsZqaTUuGH9/kxUpg
ODkWXxAHWwjWHu0k6Q93IZ8E+4jSYGhyTi3lU50LfjklOWG2otaEK4hGLNcaDopS
JOIHD+5+jdG63A7LLBW5yToFPOPik6QfN4QOEgoErpkRUO4ror5QPU8nvqYDqtZH
r5QCvfd1RZxO3Nq2dtPMM3EL8vMar3w3wYRuyI65g4VTlYFIR56d/sjmwVhJxZ6z
Jki575kLnYsJ3QhULJNky0PkDI//ppMoAz6tujCrSn477azYisJ06yw3UMNWc4ao
chCrhVvgE4+AdR0DtZeKSenjK7hm57lgdKQiQD3J+GoQsKBIQz+oJop3YBGf6C/y
fIZJw1ZNxlqni3Sb5PYJdqqKveeV0tP0nZKgj6YE4txrwYJ1dFW9wR8g/h1RBOoT
bR6h09qmQnspyDz1OtLZCD9I/oERmx1QCsSIkkGf7YP0mR3k0Ri2vrajwOidoZNu
4KgYh66gyBkch4NWhZ+DWpVyPqo8okwembY3P912cajCMV8CiGG9gMMGwPumahhT
6MDO07wwnLEwlGUd7UaoxLz/LU1H6EBAFfb6eOHO9cFCU34yB75h6I8N0h73rSSo
lm3AVzSQSK8FY/qV0SwF6VbCBWfIaolmTIuVulDiY635W5mSqLaU1EA1FN216cTk
b/7bUmAAfd8ZUG/s9tlrxUBSTL03BGKTdFHLbWjd0Bx2++Q+cEbvHmmf3TsRD5XY
5VtkiuX6q9J2MhV4lG/DkeiPGU6Nn2Dv6hJTWpTiKP3fyYl89yQ9qTY+OogoS6t8
JZiefht7cQHb83tyT4aoxfYSj3ZlzMlJZuSt+17LluFacoGxKJ99SQqSoKQp8j3u
NqgR1fBTeiTEd6yU6KRA/kd1diRoP0+pytTo6/4umVR/QqiDtSjQ4jNi9rEambIO
fgCt7EXPoCpWCISuh1wRmHBWWWLWIW4IjIBonku4iiKpHDJgJPvQKLFux/T3iEaD
c3m/5CAikj8e7GlIUxsUwzLfFEXbAeYCLjnco8NU6HxeH+xVY+zOejnoXYZ8qyTj
ZnVDPtB+5zGQCBzgB/XvszTHnP5Qs7QOI/GRCg3NnH72XBDhS3MFJgd10WuduY8V
aiSu3fpN+HWM9KkqR0K6Yfuca66sF9/mI6Ml2P/F2TMzYUjIqCVKIl0Eqo+2pQ8d
uj6Mmx4v3Aj+0aPt3LHF4OslGCJdf9U3xCztFk9kYXK5v1xyQ8ZH8XP67jBHBy62
Gicl/hq79qPq9g04ZYgc+jj6Xl3OwWbJ0iQtEBcMBk6voYwc8iSuYx2HCRJ2jOBn
IoNLYYk67QdAIIMEoPjFjHfKpTqyOKZE4aRdOGkwMpF9tzcqaXefR0wftj5bzQnj
MSXoSjPcm7rxParNKcmO+J65h/jmeZVOQwd/SD7aa/cqOWgaA7TM8hXOq+mAdCVp
582vcr48yAs1M9gV7ZhTlNSFDPspgBXDRRzM7oCm6zYEMI5jSzoe4L1Id37VyLAh
wPyn1YV3nt6aAbTcF84+JKUfFWvbMHZgnX5LQeC+qRZA6oKBjCku4S28620mzgr3
XUTBmFnLYHYqb27GnICwQkkMYFDBOVoGj5uPEtZ8GLQf46w2JEYGOyj0afhl+sZM
UEvoiLgkt1Z/byUYeX+1UxpfuAVC0060Xe2FMyP4DD/1BmAO+o8KlbLp22qgQKOP
dm/HZjZYxaIBJT4A6JQCvJ/TQv2uA9Z72OdJd/zpEyLJVARAcqS31TOd7Ihs1RhK
CmH9nScvBGNocjtshNxeQ5suN/oyCS/WlF8RwPqdOU21I9P3YqyYb74J11ITNM8a
66GumU/AKsGvvut5GOGQAhhtUoOc5L/YmKqDtOMBSEPoYa8PZ3OaUYL95AFqlctA
zBZCJr+RBIG/g7QHdGDSGwHDYkTIEZPpKtKa9TI1U0chRzmcgvis6TAbvzvr9N1x
wkjt5tDTkyO410fdsaaFyg==
`protect END_PROTECTED
