`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0agHB8yQL3vggw25RXnl/Wu5N46BMGLGe2VfQ245uEqjIgWLu6YVCPrWg8a07yz5
0cOMOMHIKEbDZRBePeuEKQCGIzClORUx9NzM5TwQJ9mIwVlmAfBTV2jG/mt23bAA
AVWyGfBfuk0DOVzHCGzI8PK/NrbSF4xai10vel6bAi9DDl9Tr8Z1XTQCJfLQUFbW
HXWlhFtE3p2i3eCL3dyI1MiOVzgrq2jfb7VJKq653cxTbfUXBHt4IxfjnCrL0Ykr
HTnEzb+6RZenCCRTnOSgEkLFVJHjjrnDQ8pgz4yr6dBmpGHoIKomZi48pRZWn/u6
fMdXkBurJa0Wr/bcqoFNiftQkAb8lHG/ziRtmSxcRW0rFtYVr0cWRYuvlR/RBTfJ
6iDfAAnTurqhAUwfnfKwtY0lKYMxSQDQv15A+u9cRVakstugKnRj9UGMkYqvFOaD
+178IZ7KbS7Jjfuo50GH/l9yVZwmRR4u46BGj6ZbcROZuf76V/jFHsw4bzZ+4XMN
vhP4YBeHhr7mfpMenXqjRbI7wbhHxqAHcjJfXLKSJfGg4J3L7JgnTC5xEVEmgW3J
JdOrmGsa6cYXMRPueKMCkNC35EfT0V60ei3A5oYhS2xHN52DIpKChGPrslI1YL/L
NdBR4hY4XHdxDNrMRT/bEluDD2/sO0bZ/Ee6O1EdyFHQQ7VELqPIx+iyvfEdjX40
`protect END_PROTECTED
