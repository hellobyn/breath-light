`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eV7Zz4YEP16e5qQElE+vFdCoPYIWStpIOagqIi6erDSuSQGmvnTDWuaji5Oy7yAs
QomDmSvj+xUV55AuXV/n8+r8dW9jdeIQQ4XGyVEMc8U8hpmYwfJcuae0PafWYpSm
fzj3jreyxVRc9A5WrO1+aGH6ujnZOiFiiTXRw108inbJ/Yj9oZKReAvtXP/rnNv0
7g6hmHcjudJWni+uoVl0viDV2NhknpHzG5ktNXK75jIIGeN1QZkfOGYPtTjV8xDh
0XLwMVINGgGx70NBtrZn3r0e2DY573G3PPUd6UaJbW7MQyB/aObamwemzyDS73Ad
JBF1vcxH4VsZGdPTZi+WN6GLC7XN5hXTE7GrB9IH+z397T1oBpJY/H/oaDFbIsY4
i3exAVHQCpJ14AIUItxEymz1pcabbxO16EbbFGLHFZId0ywgAkg7WE+eYr7rSLjG
h1xmgPmtb91QBcrkCyiKj9FQJxZ+uznUl/fmxvh7SIhr557fi7qWLdJOoUnwxaGs
mCI7sCyJgFymIfZ1bdCDTICeS3W5BgXQURqxmI+ZlAlWAYO9FhwwFIzfiLFvHUat
TSyVS83eyn/Bm7m0zqYOLhrFwhRWE5OpLp9tLCzCN1yHTB8hmt7FCPMFIFSAV7Iu
QY72OD4f6aRNV15PrW0tvGPCo+KAm77zkl++Rdh8DOkUocB31MT/bWjO6U1EMWqS
uutq0qdo5Zha2HDzM0Nlv2uGJSGUDJLXalmBTm9M2r0il7tKc6wzRcN4IUgUGqmB
1DUJIOYcU0SXPOOPB26J4p2+43sdE+8hbRAglY0bN1iluQqoqOdGrKBQ2epE2y9r
XoT0obpArsPkT2zALkRjqB8PQCvq6OHAixt1v574XVswvvDwe5b+983cGHK1nGJ/
wKSn7IISsE9A5gyu+m+vrdGLIEo+ha68w9oHp/qGMjCRwGnLQ9/zcSsd+2H/dQPf
yXJZIIKZ1g/7RmUrRWZD0awXwyi10wT2jz9XMzT9CqRJxl7qCWHT/Ii7SbVXcO4M
`protect END_PROTECTED
