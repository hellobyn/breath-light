`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gedl2p1KBgyKecQPxp1KfasK4lQ3b6dd2NFiL8vsoILlWs7C1rSkWBBOCZ2JWOOJ
0A10/oCZGCreOjdWGslVUwmUvjWWVGqGspo67V0J1NiGUfY4dqeJRqEvpG7sMBYV
X3JLzStwpHvle08HI1LkpJJOMoGk4EK6IHi2QXO2fBQbGbqeSVcqKq/d6ilS5CUH
dyc2jWyX3J9bixGu5EIqnekilSzZFGCbGR5kMBz12kRW2MUC9zj7EO6eF8UhKImN
PuAHFhKTWnNYQ7RalZgw6PR/vvnYY7XdSwr6emnqAWcQ6FVs3rzfLK7l928/5Dui
IFw5hE0Pkw9tLOoUqEwTxJMkcR35H4T+g23KkDAbHjdxdKt1YC07kJp0myOhVErA
ElHYza8Qk8gVoFQDiHAaoK4I4yXmZ+5oo0N7mVcE2ungCcCISQfeEorPCXkOTzht
Ra2w7dGxXSSCtgkz7ES9vYAUZxP8Tttb0zR9DDFgYmoHc7Rk4mDJcckNrHSSW9+c
SH4nLgpEVx/KkC5jQR8OWZzUnJM7jYDuTSXiB2akfIFsUH6dGTAZyuhgDvDeBqZD
EEg+xCd33h1ZpnOzPyrlFq8HJHJ0zCkdPIWhFEMeQ6mDGJYoJ3CMbW7pbwVjiLUm
E1WpOgaJniE86fQqoWK3DQ5BMBzIHTK+kAhsq0IMN69ilREhZ2RKTzh4EgN+uqJz
lRm79x5rXDoSYw/+S8MBOxAtSdmLj/fo047YfP6etzmOF3reb8LzYT5ZAd0mrfLB
VssZpozDz3heWJsmjG6IkroxqrcDU0CWWZ+2ZuV2qwzOy4TYfkH1bGm+azZQaMXL
krEyH103utNKmKl0vrjZGtvIuwxk5T6SCkKn74H5dbA86k021k5/vEbEFwb4m+ir
+UrjLjgPbXU6RH1Qr+3Lcf2TDN97dS2nwcFDJ4Ck8hD3P8vuWXs8gTGlhNqBxgFr
rx+sxsZXGuHfzODd7hggxeo9xhG2BbwhrQqnGTTW+5zQnygq+RYagmi8j/DmV7el
9w4gYx+EbAqwz6jW/DfSWysfMjT6o242Ze369evPQ1vdj8MQJLXO/y2H5cuKAjjX
v2ZtghdX2HTliQRedoUuh7U7Hvprvm2cT6jg/+rZrci3VDP9fsOOo5bqat3qABeF
9glhMCn9q9MI1DPvzNEYgQLbmY2jdAxb4BaQcePqGlU1XNPWuFzBVS+do9gjZasa
Bu9Q/Kjy/Ipte6wczb3ySm9OFzQWaN5JPCRjJJR6Ma60VfPV4CGDcS08V119zr5X
35ibW9pNfV+WsPQQA+tYSAW+lQ41iYM22SPGV3+8/fUPDGG1Dk5iptNNDFdkZVxA
YPWfPU5LqGIq+xcZ4jMzmWKP9trCZEwso1my2/FIBj0n8iPVgRwfy+Fk+ffBc1bs
8RqHJ6+sH39logiCbHuxbmIg8YBVoIgNHIjxz+/8ylhfVbxb+xbEZYPnnRB6MFnk
UqG/egoONEYA0c7bdio3LdUBoaWpq0GmmWbEtgMIJ+pictU+VH4NneAUHKilcG1R
6Y9BiUF3X6ytF1e3xyr5OGMUHS/t6RntLBPEWAMPN4CGYLEEoF4ZQzygp76/xhui
7Q2/XqBHoMHpm++p+Zlr9hLG0MtuT3s6FRhJxeCHv10yANVbOzQdcFjg5+uBRcC8
RtMy3igs+MIbmZ/1V7KbDDUi803hxsh4AVf4m1wyKMj5mBjdWQdDibYICzJg7CJh
BctM4NGZWwqo2YKJmUwGnFrKDRAyjPKiGB/bhYWGdPcFwi1AaOPUssnuDR6EFbYL
NI5TEdYPWl1xZbziPK+uxW3hijkvEVJ6vRRBFn8PTEnYVNF33qcFf1Bx8y6OqkwB
REmQoLzpLMZ+59mCO79J7DoaAp2hgS5wTXEa9bMfLnRltsdKACsBTve5FpeyZTCc
YuA8x61g4d0nkafAbPgW5K2C/YN/gVgZOVoHOXZ8FKh6+U/29jMutH1/tfXdMVY2
UvKA6nF3vNPxKsp0G1cnW/Z5Co8ZN6BmTXs9FenXYiqamTKtzmxefjCbBNK/7wQu
iM4cBllVhNZoizR89x2LcltQJyWsDdlszo7DIBz5iU3XL/D1DzuIEiVYjhVIeznG
ygC7Zsl2zeQ8pItmA+80Q0L08oAay/bPM6XP5fit8hBfo06uRBlTK6MypdmMz9UO
d78U8mXHYiRJ1QDfNEnjlecEQvZjmEISwsc/QgjhCg0++32i8R07XvpyZg3bZVUV
6Mu1K7qWBvKWrKTBiB1F0y2zOZJylnh71K7Tubz8tuLi5pAJfppe3UnsW/e9i9bU
UAzdF4KJfuuTnRjIzB/7VQCGOepKZtNyjKMdU54N1rb+JGDMmC/5iU5ONFep1rrg
AMgIM8DO3E+xCchcseewc8DHFgL5QGmYjwH9pxbHDLc=
`protect END_PROTECTED
