`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxKYJigPBvxkT96BoICjDibh9BJLNaWE2NVsDhV1GTZVwZ7Si2tv0dAr+FZWA8Cb
6jB8o5EKbPt1mqWkcgwHwimZCNn8NK9agLG1zrof2pq4SHUscYU2gNOKX71UMV5U
0ZL+UIip+p5WXDjpSkAnfGKgLVBtgPr0Ujt0EHHBqUy8Eu8Anms0OORqYK9OWTJO
dY12dapsrogjyte/5krFXmOQpmEGBA0GderEk5f43Fl/48BQtM5wyovsH2HmdCIb
vQmxo1NeFhw3PvQlsTyfIz5+Bl5LkAIqacN7C458OXvQlwbS91AeSl70qhly3+E8
aaZXGqhYXO609OiFeLwOfGX1OIvJSD6bVSYW8AtXK71rrRIPwHaDP9CjDTN3VWE5
7ccPv3q6SgreRZ2KFJEjoa6iI+wNKmREo0M/XRJxkTE7nOdQ4DK8VXzty5DHuMqM
JbqJvg+d2NRE41y9tNxUmkKpUBdT0y+CkqOgy9bDu6z5FI2sGLuGNi4AQlT52N/Y
KX2YGR4ueJEUoqR7/JCM1rCMU4ihZZO+fYoGxUk5zdKLEvwStogvJvixtTl+C14Q
3guTgw2FtlcnmMYMJMl0Y8yh3jkmloMUNud4m/aQN5gX7kqQOtYq4oXIhBwXe9lL
RIFPombBqLScYA3gphj5dnYJp5lfCGxNWwNktUqQuk/al+0TOT9HaUeW5VNdmE45
IfhUnHSl25LgfsAiluf3jWdMg4DBTGykhlECLt6cMCys/e2X58aE5zjXz4DEAasm
s4/iZGBeTUfA3Lir8FjZdxEpYtpoGY1Zk9174mOduiO3BZVqVsnDDbUfrwh1Md1q
LgxxbONUzbQmtrWTeO1/0Vs7vEVZMwd0PyeKi8Khn2izpOSCPDPZrmqcyY5dDEdD
gHJVrkd2HSRdpMeGZe2vtN4xXZ5Bp6ltha9BPf+bIMxilYJsNetI5jFKbgedMhro
c2pV6UDW76mL4lXswu6IHMOMbTCvBopcyqE9q0zNo9ZTMIsrWhjYbZJi/sreTEIP
y4PUDy+C3U3o9STWPf97GwALGaZ7y99Lhw90Wa06nvkV9iy0GFK9MfaBEZjt2ac8
tUEh0oATmUy7YuetXwKHhdw6t0rYacp5qygo1Tz9FmbIauhgjOOdePgoXisirT6/
xINCt/g3syZa0gyPbcWTWLow89df3XM2I4ZKx+WAKThM3TNJ0dWWo07Fa6yJiP/t
4/A/M/XwIdEcNfSskRrzld3GuQ5qXIwgMjo+jolcd0wj1m+LArZuoCHoqTR6yG2k
+wg34k8q8EkE/Jcjs6ZoREybUKIeTPyw9pxwS8SZN3/6L60qr204wLHi4Czo9WiP
dpLZG82mH0EJJnQe7hs4vnNjrh+dq0VitPNGiugBllY498xvsQsUSqgLYX+7vVc5
f2o+c6R9P4xHJ7kZ/jtSP1TAzvnjMNIPFXyFHD7jdFOOgv85BzHITXfi72CkLTFz
nqubcaaRF+p+IctxlHkNdnSrIH+hmPxOr/VDdRIgTbIVG7neHA2H3INxPkXKBwJn
Ynmph3rn1lswU3QZS0Bmyfj28T0zbFzaSMkos6L0i+/wbuTzoZ0fsizm+zn+s+uk
kqAo7YVYzE6KDEoPqAwqnkJlaD7PbI7WBoKtO3MuUIT9KxLoUjnXDcDWnGtzj0j4
YiZpSY3S1xoXJ5yKbeXNvdq3k8Pu8thOPDBgnI+xnexcbCNErxmyku8MlJKl9ZKa
oGpyd4YIjSkSC387PnAVauncbHUCEiUKGH/bpPkFkMcFy3jMwYRZS3zwcfaIV5/9
xOqaQ7L4K68nhg0kPVEkjrHd2ULvqsEthvN8IQDhyW+3bNWBxQIdS5tbjzIzLaFk
spURnVIWrgQlHtzfBPilG1Kvk8MYYO3KaaypAKKbbe0iCrgu2LYhvjpxSzRSxrvy
ZwjitPAq3UlwXGh+Iec3Wvm2MODyHUwNRASL+9qblAAKTL8ByziiH/Ke5J9xQRli
R1JTzhJuQn1vDs+PE1lew6coa9jJjmPQzygOQXdcCmjk9K/gvwXjtrmNqImGlNvk
Nuu8szWV0Eh+Jw7iMJ9pqP7/WLX3OJBH2sQ8Nyx0pggiQxW9wKvCZY0tWYrIeBjx
VfuCLkMsxhDVoElcxZtQ5I7B1s7HMjq9BZ3ro0HmEGtdKYaqYTftRR5SyhLiIRqr
SU7CpFr9bxaPpNSG/XXOj8r6r3u/6n3gbgLwWDR4ONARxBe6SGfytsRPRXKphmrJ
oM8wL7Qn+9oF5pSh+3YXhDZY9LMttJPAHQrpj7CZ3LS6+SM4GLK8ZnOXBIvM79MZ
3yXwycrDZFpUCpoq1KqGf/XUYkz6SUaJ2V2tRMgh82Kvq5JVvW4fxYDeqGgVYgNZ
/Yd6lM8iwhrHqNsP2XHQySVs5OKdH8rhNfYhcdX+W3MgAZKlO9SQH3lDFNNozwne
`protect END_PROTECTED
