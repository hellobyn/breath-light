`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiWlmaaM4ehYkxcIHSH3llyU9/wqXbsZq7xtxh8P8dkMn2hb0hNy77srSoP4viKy
qtp9Hrij/OGMMDJk5hF3ZHWKFIODfS2AI+uR2Qd9bHaWgmcPMTEivI9lCFJzDQJZ
GwjNqZfUk0JgAw1Ee+9aiQeAPuGba2S+VvRWaSQ+RdAUGrXGIHDGwFk0vEgov037
I/GPy0H3RIUE1QrVzG1hHuQ7d1XUHRLyPP8nvnJE7ZUtntFAlitf+4w3qMyCQHJm
lmCg+70vd23Ihz2kxXHjVbqKFE2JOqojFuT+S0Qh5ThgO6NA1hpnIAJVhbcmVN4T
0dkQvTg6yK0cexqsEjwMVa8KSLmggaICVVtNSPxF2uab/50zz73KNRn8JZRiMJGx
d/Uv/qRoq8j5aXfX/0t6PN8nIur3R+0Dwiy3O2ej72pBQheOGRwpuqJLRkMVwJnx
YuAjpg2vryCsAi9sTVMPIDPZWkJfjvzqW+R94ZtmYv1JWIhi63nwfGYvcRm29roC
1yh84SYnyy1q3Wd1jSfggOxF21JnO1R+CeAK7q9oKbdZ+SKNwP3KGpLT2XBbsmmI
7V0vjRPe8431ouuSy4IDoJjLcmcW/vHzfzLljxTQv/VDgpjPq+5P4hLci/prn/UT
6sCiE4Ym+mTQDrBimNutwVsc/HwQCim2hJ4FrLiSDNDn9A0zBssZU6mmywfc0106
nx3bvnS/5smDmfuVgcEbVJZG81WJeZW8dv2QakRu26BWa2ywLLi/yugmm9taPptE
PErsIsb8O3gxAEA4nhIlAJOphWGa/VItGJcFVimuGxQ+B8yB2m5MPHJktJo85XSD
KGk1fRQhHJomCIF4jf88olAaMv17LIgLjqNYjOGmdgqJN3vjMc2XhPd9VwpYmez2
bVcMtUNkUunY/wBvXe27VESESI2SYC9ghPMFlDEDw0RkEhzMo5xW8WVyfp3+hlmF
m21+/0gyrO5q3NLrtt2GTuhtO1ejluhexVux6g/kHRIlG8a/axRyxQ0pAWblljVX
SilgDa5+znpoFQYr3abThMaO9Wgj8hp52+IqC3VefCVSRRhWW/RT7OMA2dCal4lX
MEEISJs3X5xNV5cNpYxlJqIEz00nfP79zhxLSmbn1coA5ySMGlayeND5Tmj0/rJ7
+yHduvYan/sdGKoFiDcVVVhuSW+9/wVhx6UxJqCvcvQY8Z0GjEu0GsrBrAG3v/Cu
4CsNoRXnt56/ZGAhjwp85lLRQLQ6RafWHwMqXZqv/rmZaaHk+IKxbvJZygp3ksaz
DvJMJn8Tt/8WlvC/kNs97+ZcWd0SOP1/D+OlvXld/aZvaGZbRBHQyu6ZN0YgzVlC
gTK3WKAOXZGLoWfk0P0JCoFXg989GsDMbzVbOr4s6L9pawD7b7jtZm3Z4qvM9/h/
AWoJ3aiZggK9lFlpw7x/I3L5TvrVodVDnJWtdCiuqRP8nCIuHFWO7UH9+a8qYex6
pECJmbE0WYPAst3TuQ4Uvygwkryp3naS3N3EwB/OIwg7CESsUsdKM8GGXvAbkgOV
kNV2jub6YFXcmyGNCDZUH/mtBxqJp5EkHGpdI2H5ARmlWwBX/i5zLrzOK3NbuXwe
gxIpmMeHcvPJFxPtgq4arXf6ZvQhQB+EljBHkT7fnLWobpb+othKYeJCkc8O8peT
3oHQHPwT5MNxsUoa/b3VMti6PT60z3j0yfTTFnHscZ089vfHu2Jmz9I9GPfnxuX8
`protect END_PROTECTED
