`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bY8CwtHdFDufHudWaJhs4Ec3AGVQRxo5YdGV7hwCmXe4DNyQMMyFxl25GhYZxBUG
fTG2WXMCnIPfQfCt7fmhZjsuQg6qdGjH92MiAp6186YKlIT211gbg25YwmTbUcNB
XTGVzqU3r8WSJNZjahEi2MOPxxtDBQ5a65Kzg5JjCmLBk4BkLUlJ4weHIIJJrBIv
xb5yYhu1LJ+mXNuQQ1IiAEMNvdPxQexDjORe5U1bon717JdR+yraHYuQxHP5MRZQ
EF6HNl2EuvMfxjs8cTR2avcH0YJ4244cwm7KeEZi9DVB87s02ZcssZREaNARe8HV
1CHnFUy6MkGBz9CTAL3T2oz5qpUjJHjpeeVY/sglCzl5ZshgSkPSC/n2OOYyL0sD
xYxDTCTutr99jzMJC3aj534rix7sq3/DWBvL55sqZT6c1qsqmSxNPPouXu0UfKlq
pQTEvEF24AE2x5Foa69o0CDV/2Qx2yWQFtAFXlOdAeWYzFuz/VU5hfyA8PDJM7Mk
u1lJ38aQFK6/nOCxIgUV84qiLsQImnpjwr4fbAfa/tTemwT1kQ2gslQREmF9pVwh
vCrvJ//xEi6jInAnLmqijJENbQF+XpqKjY+exI3QpfuRBRgEyrIC9uAp7eklRjFj
EQPL4xVqG1kR4oKGph2POuArKxYkRpF79g/if7XmMbLfvmzdk/E7vMW5NG6+ux+D
RcBz9hLcGvzQTqPE1N9edhJj4XozxCxsTEfb57zB50oAJK8LmmE3DzWmbAb8YAcU
yyxcmI+xT1x+52TRZXofeZ7Bl8ak0gDeZnKfDWMP3M8FmlDGzG30GmSNihYErrXQ
dIpy3FdjYbJxEi/eSwyybf+QQ4gpNQwnbsRx79pJqYcZNPnIno6HEn8WOoXTo5ha
FhCVfOp6cRqS9MQWVSHbmh5zWLusBnp2x8VCRtBmL5JisU9H4g/9lnVo/GHCh6kU
h+yMOWfpuTe4v9F4eZTCKd2i2p/ylkFoK4IkiTvU1ZqGw8ep1t/UvAbvLIVOotvn
zt/ruHbJElMS5UCLi7FDuUndAXnZZs0BgbSb5CYfbXjB7gQElrWbZ/D0ztzZnubM
HhISVAYEbTHDD8mRoaH7IAgO6hZE1q9cMf9kYaMsHDsX3LYZlGZNarrDQRoUWj03
Fr9Tgp9dsW+v3PsBHpMFpW8SWbWXFtetDyyjqBnvdvxZqGSC3BzIqnpMHO3bkPky
V2MqSGRWuLIUl5RlbGfVYg==
`protect END_PROTECTED
