`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sy4VDW+csJTvhcaQntKRW8r0349aIXzAzsKOQlnxvxDvDD4Q8WQDCc+o7wDNr7vR
KmzPLPONSm9SzVRZFfGHLiynMAIwt4BmybdDXBa1JXUeBS3zSk3bhd8GL8Go7yn1
lmQ+8MiQk8eZQDEJK68c6H2r4fQPFvGFCADqQRpFpbYvcwRNvJ9RzfPo7DhQkz8W
9IfMyzC+g1AF4qix26LKh9QuFGusjt2syY9ltYm6TT3eshIfr8hca228OzDDiBUs
QetNwZvM7DTOw1MpngIyj0AjeKy4wkNE5WgRh+Vx4KOmtrH5uJlJV0w4EBJbFQU1
0dSQ57Sz9/zofh4GwXyqAdQ+VCsUzIEgJk8Yjo5MhhWgIfICwR3yam4xRWIt214a
eATcIM2JO+Gfipc/Fnt1mFYqTkwQulFc4cnQGJ6/LKcGTyHRPFzRyqdg9IMn+nOp
qaRMqnnvCGkFSf0P+BW+kI22aWsSTzYMj8AQG51B48aXTgOcE71AtXbs+WD3M1L/
xS9vARF2thes41U2unlEaxxwNGP26BxLrTAfP3ZBP1JBexpdboOFbWVe6Mm9Emwj
5dmjF8H5ZVtfW4dTKQcG/zU5VHHbsOpL4OG82MHR66W9yJRnpQBo1d9b000+OEYE
IFQXmrqm/hMxZVEnQ1QIGwYbQYSNIZfzuMgoQ8v4UocAJsy0D6ajTzK5pPHhF/Vt
+8IPS0huOw8Y/7MWf79POOuWsh1KFDrtumXrSPYK+l4+2XU44uxYCwHq9X3+OxxY
ffC3bB5auiZcP1okxdYJAL1n5UyE+OIuaBg3RyA1t9mHqckbqjVZVk9RSBz/Yu2/
0cnvh8LswEOLi1aQVJeGCTLlwiurxG0rGjDpL4UEoRv6UAXBC6/fLYiv6BpUGmFb
hRuOCABnsHynwwt7+jAzATz/IZaRNTQ0l090UKeyCteFPyaKy4SBlA1rjsS9bULJ
OasSLM0yrdvxYW+c/tpB8jq7q50PkNjJrmeBzq6gTrh6RBnFPyjNRddns6jZZIyn
wSRzvPV2x6CxbVGJoIdNmk2HHHkrzfaAuc7V3xoVstjvBRP8/ukH82kiFJIoSuKB
LPBWV/1ezQMtvYtn+bkvmGDtkYo+n1Kros0UjSeimIvB6CvQpFPLIMiYEqyZnVez
aKUbiMhHk8Ck4VcV1FUqUKUpdKvl7+W5OmXuNlL9VIKPPaoYsK/AdRKMsgUIwJiM
WV190wAZI49XnLd3UZoWYgBfAOW7qXeDqkC7eIAXLF6b8pkMSo1v2NCyPwi/P2ST
D8IMLRHKQ+T3ijraCTgSgZKd3a3aAuiBHTJogttXg7BpLLknNRtKHHyMXVOSWrjt
LCJkiWeHXiqjKDGvRVPIxV1vszswEVJaOCKU7U2TbVQBHc0UkMcQ5HSijLx9BgY+
60QLWiLKvRlmgCPKbtC8YKpqlprLqxHmuNHFTCCS2hyDyDh+3ZmMjI2YvFj6B16x
tuIxM+qbkQ153eLiACAe5eX2dQf/ijyNMTWyr6XbIQcns2bOP3vz/d9DP+KmBh2m
HkwSu0343uQdrIBKDEZ+4EffcdxgBc1TQz5DTvzkPn54EQfHDJPx3SOUixiGT0KC
h74RBxnL08pHKSDoEBH/t2Jwo8AA8EK0YcJJjeHrVWi/ZYsuY1r/CmuD4JnlSGWB
oFxyDBHkV5pKnwnrWWRyW2XG7mNr+9UvG3yRvcRTuBv8Nmdz5K5Q6ONPSdgibMYF
ANEoX7cDkNsR+cxio4hYUVIOqUCoX7amtCO0ZUjE/AZ3kbiZM7aGzjLWSwl98dLY
PZzRHvqsadcJQLp/o66lR8qhQa/KayMF0taBC+IGMn/mnTqcYZzvPXIteOUHwiFf
3rG22YMSZmW8/6WLx8POtm2gayHkjUJrmDolMdqK6+MjNlbwR+sVsZ21CPDsb89g
8pz1X2CW4IyraxazgJ+LkjBPyYyIhbHNa8W0DCIjqLb9rAThYMjUXot4mNPbP1Sm
8dJOv6GcUbouMwRTc9KVC7l+JF55H601gPQX87p83MKAJuKSzF3jOmzwXN0/hhGU
g4lUo6pflcuGZTPZpP0T+XBcYYmpTn3F7X9f7mhRO++qqqpMfTcCwnNpp8DjXSlr
s8SuLtzVTFUNzbye0u+orSchux/Ye/LxZ/X+zoGkGf9+9Jo4rSfipLBO2ggiEwnv
+ep1+WUph5YZFpm67VCJXI16ApefrUugaw7v6jRdHdZ6XzwblGIlJzkR5tvJ6F/X
lh0lEUjt2PxxRWfo84N9YiuJSpDDJBgORPZSvJdPKdnCx3fRD9ch1j1Vxf0X4oV2
ak+KNk5mpBnhPzyAc5HzXd8o8PBDIA4RGMuDxI89d89cLhz11vvwARz1c3jo1CQX
nwQ9PBzme6VZsIW32m+aJpoHcgDTTggxzzYx4lT4wQJW4/jX2pnPKXVQFRYm3rZp
5LiBev1sbqiwkjvGTd1aIzCHx97HlPK6bgMdKEr8+/k1MAwjJ3KP5zgmObxhgZe7
Rp49PAC1rpG4X0BKeZcp6wgz+mgpK/g5FM0ZIamWqMW3h9TEZKPk7hXKIKUnGb60
jMu0r5vawcpacOoc7mLs7QW8RFN2lHq1GkCB2ujp/wpeitRjIu/civOsfvQZWE+E
eF74xjt1tLyMHaVe2lMavsXkH4QGTHO3UV3iX6bk1vTC8812g0x2lmSfFqoYREEp
fnx4QAtxHkklEpwBoFLdscXpKGU1wifiUncDtZMv8eaiqsGZJ85pHE1+PjJ7kAf3
AlLCG4Wfcsvk5dPtdfQ5P87jreGlxJVE2MOrvfaDPpmaoTq5r4nseOoVVMwp0zJh
ZiG3wKMvM5OfniCBl0V6Ytk9HaduiQNyOytQ8lczjgjTNjsiCh2+00H9HEoPOZbg
ClSJ273kjGJPI1Wkg44lYGT18oBthIqHiaKkXyRZm6HFIQsA8FkA0WC3OMgnX/tU
7XKQWn1anKpghY3txoBzydT+H29zKjTqzgbweU39SgbYh4kc6LxQLiCZ1DIt78tg
Y/kZk+kiGYFZa2yYzhBHodPX5/lHBPJgD2peqSz1fDO/43gg0vsrah3CkbzBF7xy
h0aQjXRash2QQDnR2GX0cdTepI1At6COFufmkwWmJqIMPMsqg7BSpgCH0/tMuf1F
42m6GzYYqyg9lM34ipTpQQK6KneV6FztF2J2FDv0KY0Cye/fDrU5s2Q+wTQNx3wI
XRBS4FI3kxzP2KRjfpiq7eldFbn/GXPJb94SqrKLOHfdnkdalZ5ipy9sAMLIuUKr
O2Yx2dff8bpWOYcXPeJWsMz2CbZaVtw2zlENhcGxjB5T08R3TABVMh67LpUyNBoH
m0mIdCri29X0+6+JDvXF+SH3YGLGlIT3eIqHryBAUXVZ+vY0uyCRlQbMIo8XwgyL
YZIdbizF8P9KevGRO34jZVGZ+gbk5Zt+K8k7iQEO3YaOUNsMRF25OiWTxB0eFRxO
UDAKjcFmJLy/Cw3H7j21mBwyGStECqW6+6m6vIwpHz0=
`protect END_PROTECTED
