`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kzcI+JmLADUfWceQxlN9YjHWF6HvHdBFWZGUmBz2MCYRyCncSKgUvs9R1n0PlqI7
Yj5S0BD2h/l+HK9lBqzdndzNabu7iHfqLrRBOso0wDR1vGynk1i6X3iKI67E5HnZ
E/jlUnPxqvGH1/iPvSjBtu9DOE0ZZtbto3W6dj0iHTp4g1vTnIkOycJ2rD8Ecvxy
FkGKL2DbMK7uqaE8/N06aBg78FNEiZMZZ/6nxBGwiEGVA/mI6IYgDmw29tYUfQBq
nyt8H4cDYIKmtzMadYN53/3q75icSkQpk58KyJtqxjCRTqp+A06+9E4bMSuI4k99
jUVkidCBhYHpe0WC7/R02GWpJJ6E72GbmtzGdLYrbMadqtgvK0Ms1AfUwSNjWg5F
O+tV8JlHXBQD11EGQ578Ie6EwdJIMWKn+0fjfclxB11UNsjfO1U6lUZ8EboRHnlZ
Katw9WgtcJNUrXH6OBf7Mi9VMDTc4vuSkjfuCKwUWHzZsmNHWUTRrbaZRau9CKEa
MpHn7lPmmvLDsAvtnf9WXheI3XQakKro0NANw74ZawOVO+6nAw8Iv/n1x7pAg3k5
guEvv1/1JHPSACTk2DB/2AtUNNoA8fCWHpwMfOcVvx6ET1b8CkAmM5pz/dG+YOOy
QzhL8duBzzahIxhFE7mwW1OlLfCBhZpRtwIxQkKvNSH/QQMY9eahFvS74e8ioPsq
uAMcnpl/GzKkLUvT/0LZ/R8QmMU3SqbqB6BFdgsMngvNmSJp6rxoiNR5N3VGRURN
4Zqzjc4ZSO6KgTeNgykXJHMELP88ESwYLTRleavH2vc9NHMAYnDKs6k0Nwjzmply
fO/A4qkWF75TVsSA/gKcuiT37SgfWY/vmH5wbrT8oqfdbhtpirs1d9J+ftbx2Aj5
jaTLDTLeEa2uHJlZki9QDVjEPN7Qr4YH0rQshw6TiWncGjQzp7MYGjxcMLLY3T3w
9K7ogJfc3EsBt9ejYOjVuFBp/n3/Wi4o1spEbgDQGXeAQfBCLGkmP8gU2xXTm2Qk
eOVZ5l8t4z7XY+CW3UQJ058uLujAbE6qhKoxa+6NbK7NVIqvix+LgE32Q6NprzH1
x28tasbkao9fbPuT9IryNpZ0yLwJarArJWYyWfN2FvBWsYfzoUnbt0fnubMd92it
ImsDAWCUu9Qya5F5EuxwhNf3Ap355PgwUxvGzMleVeVpZhwEcQRtdPgetjvFAGV8
qEd3wdtoFzvzdq8K5gAYteZa6s/txXVv3w4brMdjPDYfuloDgCuTMNDtSFZNEGLY
+y8xpaXWy+noZpKr5TrTIoYkDYc32+2a2Lkr/jcPbkBW+64p+nWqfylvnmNHG5jO
SCKhdlwWc4WMK8jGGmkvkZab6Q0U3cYlMW9lLrQOyVZOLmwThtoFeCLxbAv35oqB
I0l9Nw0890sEjafq7JJiMHPjPq/kgFrF4OA/0BqO58lIV1y+zgZq+3di8VPBblQj
pg8jgGVcabOYjggMyfuG47KspXPEOSCJxiqu2N0OMChuWKa5wIqfiDYqsHp35DUP
IWsyeZylBc5gqu/Yal85JVfC5M+dmv3hHhsu9IRB8C7ZC0FDorlxPfpbw0/zKv6Z
vDltUdpGgXldp7Tq3UIgweypH+oLHHrqmL2pECu+x+On4/C29+tbdTd7h73MugF1
Sb7lNZ12NRu9JducTEGDl6pO5KD71ARh/Dbk1n4DJmApznMf1jjBuWYG93qLGKIT
JtUvXcHfk77IcDthKe614iurFIcbdscJX6hFUIy+RSca8COO74BVyoR+q/45GQ+X
R5FaqYVozZHuQetYqrq9Ww2QBCGLLeL2kA60VLnRR9TmKyc3kiwaSSutgOUsob0+
Vu9aoK3xako3b1fFjSxAN4Pr2iRkh5r9J1+sqPS8GxZcsES20wPQ/6uNuLmnA868
b8kfqX5I/cwLG8oPLUnnPkQL9q72bDQ8Qju9ya7M0b+nGNxb2988RLn/I7rC6QeQ
i12aLJ2x8DO3HFC12dyUdCfGR7rZ03o8K5yPgXkeZZKzqy1FWfEJiNkg6hMvMhLa
mIa/L6l6zuVI81qyqtpJ4lilIvpJFUDoFnZSnO801bPaMHJ4SSLsFg/WchxqMDG3
fyh4jcNHOEhNkm3BRr200iQkVtWurOMvRqZIqUoTFwneYidNdxa7Y6wykOQrPYPJ
Zkoyqc1kDuv0Z97VNixiT2CWsMioUiynthXwo/7YEPEmijnlETM4Bd5k5VaU/+6v
Y6w8H6wY9h8192B/V2Hmv2PiIlI1LPOkZNkVFr7+TinjKX6JYZE7qrygWKnSj2vt
c9z8nSKjgFeNO14dCNsOzHrPM5TKJVt3JNfBSZVks12zKMFlfZIfx/ijuAL4MJlS
mnuzEINclHE6WMI60750leZO7iFHFMCDuY1WeUP1fyZ9PbaFK9DYfPortoeO0gpn
7NxSGV1WBzoae+3D2poKnau/u8CdOfKbwbCej8gTLoMIlWEuKVkWMhuct20TkdoG
5Ed0Z9p+ncC7YGDy3LyGzs5uRTI0qqR+xafqfJFHgMEDcedBYnLwlK7SYIBMcE0T
uido6yKzd27KXOou8sw0GDYm1TxLLwtpFrn3o3i9lmpjKoNiz+KA6qVgt+rXpV5W
GcDwiTbFspTe8JRo4b8/qsyLNNKe2G4NzZKjPCxil9RIpWLi1dr4yvV+dPDLgyuN
q9X2RBXdGCszeDZyclYjvHYSrqo0zfsGPd9oUNUSIgnrxscRs51pZO13xnyhXUPc
7/VngUOwKbJk2Q6BklgFT3hsp2uymcHSGY7GzsN8wAz//7iLkxQbYwpm/f9FCkNw
V/VyWXjujvnhpjF6rbyvEeB0WLNI6FBDZDLI5P/iMcH3HRC9VkxXXtWFdEiTBzcp
9QfmOz5EdreGepnUQCwsOaqDiNrClt5YqhTDHsex9qOwZmCzhMySYp507wMC839j
Twi7ynnR2dCBdzl8fKLQG0ZTkj+XwVnhraig6QgVo4Ov6yZPtP1UlZalJIJkryzi
w1/gg3dRMsV62B1BpMqCVYCU08vdi6UEMp6+DXBmIq8BwL5/oEVXvLyZ4laT5yjE
r702/nmvZveUoyA97kqJ//CdpNav/gIYmKKupsT87brjdteRocHbvRXvnX2uzUHE
TcFQZtlHRgfuBBG9U9g3x+VX0xmACaOMa6V/Yy3dj8GS1OFG6Hf81UcBe4WK9Zof
qIy+DM68Tl2XQnbWH0YeRsnwI5PU+7dxrIq8yF0VsCv3k2JoW45eWELOv5S9JzBq
VWpTkJVnuRvfnR24OmY2u3POSl68EZdhHkjyfcXlX/xjy8BBtlPw/xiss8+iHfUu
My2iYF5eP9pbewE7miwtDzd3UIgv580yh+9jZk/bH13hGNnZb1qkP5YpQfj7KLLu
zKZGn6zrDwdTwxfrPzTZLzojwVJMNCxz4C1/h3jeFoVx1oDJfs9LzSkqEqqf3Pg6
erOwmRxeh1zKc4xgooFyBgYBTYcgzzvRkqauomzDpRb5/JBO8VE64G3gC9j19N+G
uAgcZhKkKLJSk7jys1ovRnAI8V5Mt6fESSnXGZgqtuidJDMwICk6LCQXpurURu/9
2uyMxvf8IIENwfa84afGbfV/5b+zyh93vFyWTJXnuFC/vkQjz6tgDjrdAwMvYljr
iLcRQ5y4QChsVTu6PXsd+NbkfD/Fwt5/6lTACHsZ+64t4KdcmkVzXE8/T3mt86xj
EQVJG0gpb4ObkDM3TkEJuM7nH17/Dmi3NRbz80MksWKQ79Z9JFFW+fpd2XWuc596
4oCLnzFZxsuPrHuCXLayxyAqsMrcy4qauK4eZl1cfqdbAz1rEMVxV9JCV4wkwk5l
773wvYFYONsOoG19A8k+j2oG/sfppFPjUtnPutab9yOFcbR6bvIOYxMmLo3rIWgc
n2eUAOVwfG+yA7L8oHPK4OULmeHFA+WwG2EeVfYiUoiatmGb84F5CH6CkITEJ3Wd
YGq03b7CYzKZD2D+ma0tB+Vwq5n9nQrvcrcrqnYPqDn26rIkS4qNUc0dAqtodap5
4KB9wsydEYCY87x+vpkFrrZLDZkY+frPyJvg2yp9gp3+JkzzjIZGezQArc+yfZXl
umdf8LBKrshPvMmEKh90lBhyt2YoGRAftSA9s2s8OQIAPyFcNkT746Okoibq2Mst
bGsIkjqK0/gKAApM4SYVL7UIyYmV+YwXPH4hQcogg5Mcegys1bZBe7nrxtfwKa9w
1wxj4T/Mn03g3amOvj4FLoJVr1V9QBXNJqt72P55eVkH2eY2PDHvlJ+bZpfMi1l1
LWLkCZAGcIEewyaAsAXXc8f5jeSu35llwJGOEmcpAILALCJNJA7UK7NLF2hgL1Tf
eUjcwU/PaoNEh9h+KHApJO1fN3Ys5A+YHhry++q35Blv4xpE/9IgrqsTxEgqn2pR
anIp5M62Z+RpYGvMV7jnYfgFp8H6VLrFQJkjnh7RvLuTzHBY5tQO6kIqRmVEbRNp
yxztQKQ2G06GRHpq6CnLHv1bLogJjGn0Hxl0GHzx2RBFJOVb9TSfeBOhRgdhAVaQ
ooWlqYbkjgWj7cQPR0BaBX3LbOQOk5rvr6RpVfmY5flXIwloC0k1TAKPGTOEfZSR
84kStnoTcyMZNSbmO0zpeIuGi79o4NNix/a0Cp9nXIhNuzhlCw7/jyQreY9cfY5i
444lK/uu9iNlen/trO4JxnCepohpqT1V32uHOz1e+eBQ329XhbEPQRdc4uqc2vZC
2hUsmsKuwxkNRwWIhwyHS6J9HHabR2o3gMANuSDiPqCwEi8axJm/f3VMAMalWozb
UKWB+VEBvLCO/8IgbbZgLYISfVosyHAayFuNYfY8J2Gx6ajkECgEg8rmfKBQTNjG
l+9VJFQb1X9a2BrBnnjze8qrDAASrmtp9RNBvSPycdk9hMJ9vNQLWLba1NZtz8kj
Zt/hDlkYQZIrb4DrQ2TUDFdOoDZkSdVyKLQew5a74l7yG8TutoN3tq9M9h8UGhOc
pZCy37F/gBKsUvX70gBlDb2CXwavgph4eudWYOKcU1njMurWxu2hoih5VJGt19O6
2PPBIJvGXECNqn3cdifhMbnkBMSXv1jAhOj+CNsWLgfd475jHlqqAQ2tv1fmKgP8
+CD7MEA4/UkJW/RgI3/MCIKUGduJm5OpqOtVXXBLsSO+mU2bFdLGiyzOW4YrtuUd
PoIaclKF7l4lOihSVLECv0xCRO73fcFLEidiEQSlqa0ZrSMnRr4v3FE3oMdLS/KW
oDbIU+UOZKgsVVWB57CgWlqXpGcre/cL0iIgk2+1K5LKZCxQVmtLJ+drlsEP1jj8
v5MnwMR7hpVLAHO5WcB9J875UgMv7ytr2+ArTGFcc3xKnLSgYOr1zfvcT6XhWR/2
tHdWwHtEQummHiHO2nPezzgeysuctMdvaV3a6Hqbublgz6P3YyyAzSCJRRFdrsxe
NnqOxVEEUUFu0u4hStqnPqL6dzZktoaI/h82KH/P7bLCP11w8SE+J9QEXfCo9+0O
JXbb4ZvHVv+G1DbHpO+DDePOkdZWAvpVzl635fUQEbwCh5clB8gJFzkkZpDN5S2m
nJIw2JgBitfLBcfBkJ4W0fnj6oeLIdtsf2mqIqSNm4rGGQedsvtZT0ToqJ9GTCQn
w5DUsTorI2A8+Z+LGeAbr4iGF0CTTDUHuSFTUJDWA3ESk7J9B0Uy/QGIkTemxLcj
ifecfGSvOKs8T1irNUOql+wDKXrfulydaQcN+DbJjSqng+iGK4Ja3pKgiJ1QkMQT
v7L6hoVqQ6v3DGXfxmXj1R+BEIeSghVMm4KTdOjzxP6zQZ9I1qMIxZ19N9wUbNba
2ml7Bc5hNtSxT9lzzz8SpYvRA6Tms3JtGHz398HlsSSFV5jPUSBVn5Vs2qtlu1rb
Lo8m7umHZm4s4AG/86a2OVBy7s5JmlFM37v7pKR/57kTMJeE8aYdi2/AOnUGSivl
rSTjw44UL5NVC05EOHvrglASvgA39HWF/1gVmQnEn0l0aiWwJnu4J4tllDiG8WcV
c5akEs53fVc9Lh0qlwWTXUf1+oMNCb9sQIwCrBxfdQjUU0Mrh5CsRN1CtkR8c0ht
W9bAwQ7fCB5x4AwQOdskIYXxURlj0iT89jPzYLJFNLaq3mBvovoIVQt6w/UoHV3p
Ufpr0Uaz8v4uMkikTXpdpRtD+nJhA+wVIObLeHF400cVfLcVvQ4LaP5BtooT/fyP
tPiFZE7Ah4MKrw1cYZyUSSUzzWqinvdZVkdOGhvwuDhnz79pwUJfg/poHQK6KsSE
AOGPuUrSijDMAhXEufCVDUCHB2vZ4ob7wf1gwZnvoadl0L0Wu7FNWl5fFjSsCAdI
wuHCEQOZ0wK0tZDZB0FTRR0uSoPjUFza+MQ4sQvmgmbj+T72fHWUrnVedCq0GxYu
mChgbEqHcF5OkO/acZr01lzCpNDnEuSJlM8NO5XULcw4/nFbp4A04N2stNDi/rnK
HWdGr5c/hPYSg6Xu64oJLWUBdFXYdKSwJQoWnZwnHZTAzipAaSLxwmwhGmrNQwqz
2r3oCcY60xDLRsyHUp54NxecwQ5MMIoFg4EZs34uhe6THyvCfkciWNDoqeNNGlil
BY1lqSdA6prEYp3eFklK6pi8MNUJG7+XTrs5bMWZdeZtH6qX8zg85acZkcGI18NR
9IddS9np0X4XbgpAnAtvLP7/zQ3l94sMuF5lTNGnSL7frKZcERAh+/lSVm3dpFN5
Dp3vTC1J8etWzC3blzqVDiNg5boIg9u7bqnGcVuAH5iiji0SLuhjOgNlM5oUkbUu
zsw7/+W2FTGZU1B5LkTbTgZOo7IYBpoU9oPom2gSCAcbfw9Fit1ikaPciME5DjGz
ckMoihZf6+MUJXhAlxm0orpnA2F19xpMmhJnKTr4Uw1gJ1G+nTxDxt+pbJ6Yobqc
0yV/SBEWtExQ8FA4Hs+wpCRPgGyPUN7xKfPsyYkOPYiyjGEwjsqNxeeSCXCO/iFn
5k6QyeGH3IUx9ZjNUVr3gMsdffQEMFiIMqfW7WzenBdygsgNGkK4CxAGX9a7dLWX
kaOqbv/iPu6Ac3cxBt7xyFPWy6eTIuccmaxEV5lfUnJ66SX0CbmYuUNq3l7lr11P
JUOwGVMHfGPSrTiggC7kg/P7BqpiKAb709giqTunvjoatrILO81MfniF0Ap1d+XA
IYMCnO3XULoHAmHud4Wq++b/6bhL/RKuk4PmkQ/ElMLxUjtJTB7hJoU3KbSclsmV
ztKLrrNCzFL4OQ4RVjHtFmxyf/HkKL+59qO+qC4z8SYzVtS+CHq9+rdBsfjclcMC
vzghYw/WUaX47ID9jmx6kguUl2yGrkd+2obAwxLQ2VMwuART+lVFfeP5L+N4XDBx
WXNNmFsISP4GHYNcJAslkJpMi+wA8D7X/FA5I6bTDKf09nDsiRLIXFLOY4F0dluM
AWv/Ex5RaVOskxs7cDbxk68lMkPpDIUn6iLjfZzvSX58w1Qwh7WKW+EXIUKBNCRx
t6UxE3oxeL6V4TKIvO41D82r99hVKSxYTxmvovyQmixLbi0ule1HzTcJveXR6e0N
QMiTmwHBmNbciWAzXfFTYS7XrRhlACNMjlrRQr96Y7jxbpcv8Ob2X9xnUPAmHI3+
YGC2y8W9jh3w/CirbYv7U1A0a8tmdjtsE4Wezgl5k0G729WvSF+pUVu3aFjvOX8W
qUm36sCQmQnX0yYB86FDjrtX2wa/INjf4MXyweJSEOMD3cG/tHFwBoV428gKSnu/
57mM0+nHX7pCUC+ymjxxsh6gM5CkI75Cy/yL9yVs8Hxbt9iGYXxti3K+zaxkaIM7
ssuNJXGAAcsvA8j3UWZIN7VHNjxTEqdBgUhKcrZ9tME4WRCvL1PnUMEYGKoCi70d
RoPYL9444rFqYwmlMACm0O/jpoRW3dky/4N/U7dI2GEfrVvIhbde4ww34pmwYdns
V5pWQwm2hTsUHh8+x97s9RHLPXTkT0+d/WtbWPf2T7TvF6+CAT19+lNPcd4edZi9
S3MXmpS7dylUpYE8Gwj3ry3buDuVuHQbAqrqo83BubPOAmRSj90KJ6KhhfCTJOKI
f/kWeV55FqqmMrTdhA3GTrdi3yzGfyuu/SPmpU8j3FRbisoxvlZY4QStsLLRkHDm
IDCa5kulvKGXQP3qY+ppPANZ+iLGmQySUbU7SZUdbRMQDVV1NJZqsPki5meSiGjy
CqMk8O6UhWyCqT3Gl7qo2m1HcSMmRWXQ0shlvJqc+ZMkP76/ccRqkrsSlB81AVmA
7X7MQ3ZyQ1aosEfbtT8um4RTnWOBUhaI40N5bFuFBOG6dz3/PA80MxHAwft9sFoN
rO0HbakH4aKfBjf79244AvShYe63VFAym68lzHAAB0FApbYL5H9H6jMum8XkFnv2
NkFE7IZ+HR7f7WKPk/67tWM+fparZhESjbkN09Rqt5LS3t2mI/F8DhG70Azv3FA7
F0IFjB/+0oiziiUPPM7gxQSSOK4fptWl76kqW2rxF463hHweJnlyUxNI1y+JDIK8
CrlP8tNGnXqyTz6d0Od/GKA4WZ1hGQpRoG5/DoKjog4=
`protect END_PROTECTED
