`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5l1crpXu5O52KBgAlx2SXCG48e60klMdPI0WtsrKwTAL78lDCGOoCUeFw9Nduqcf
Io6lLYX8ysp+bniFTgQ0GtTXEKRDlWYqnvo2no1vJijxJoqOsWIXkWgfZeb0BC87
2gJ3EK+BKdMd72sVJ070u1INbm9u0w5URfFZBvE6blmfcRBgt9/4G0qEdHBtPQaE
8GFGQxDgKpnVyju6/EGDTcQkcV/yKIck1ovho27fjVU7fMnnWXSWIcaHALiOeynu
AbfLwUKEtLrDFF4Hks4YtDyS3iJQyiX8OO14/T0uhmb1ci0ilda3rBhaDWSeLiWy
vOKCp0a9/ubui25tECV8g40f8PP1ri+nzNtLnKO+sunJ1VKSPhK7R8fbX/eWU4UC
daAZmb26Uy7Iw3Xl+fx3E87dwizP6TIUZly6JmnU0OK323yXbUBWCiOdTPnlWwMf
RzR+VGK1UtpXgpOey3HjMA8RPSaYFkVc3MXXJO8twOwXav+IeXW3dMK01tfudIjZ
uL4M/qGE4RtFW0lXU/CKNI4oWUGP7XWR5GqTwUmMKcmAuJ8XFofUj5ZMBf4EZXsR
zBnEuBosqrFgEE+kcWVY78dUk3M+HynXFMfd5zuGxUkSbuM4U1FGFo3EyESq9XGZ
/C/Eu9Lbrm9oRVLSNyht78X0PsupqiAbSxVX13pWVJsW54lQJ3/4Dp0bvHbnaNXh
Xkg/WYBLcJ1gV52FTG1hvOm4gctJi9mCfHIgG0jOYdpThyBAXd7bZqC+sXwSS/Gj
5tPZ6oIzPJhzVICfr0bxruXps9fJ2f0BYalf+neq1TTSiaCJ78p+VIfe2ULZyxf1
zmfvvooAQa2k4TYYgQ+fpg6V63y9z0PZ1+EjjLvVES9J8SdkMN4llJZGyj3fEvMi
E+1957bjgjCN27cYFcOM7GnyxR9wiP2zUE8gNXaCVWFbIMyIFZzcrk2MO+dWLJ90
7gH5nz2uFxEWB+Hh3JCmRi4TAsaWVfE6HF9u64tF0BJfxm+fH/miQWlAvlitwJ3G
QlE45iUY6pAmWTcU+SexcR4+lqt2vEjURkAxydLP3YWszcscNSRSEIBagK03gjhv
qqaKaCO0xP0mHS6WHMcxE/2sMJjEenCyJz9MLNCk49S8Ko6Lh64tFOyP4nt5sGCG
vPrsKcwPfuD6bIoaaZB2bzbmrMp8Tz0XQMvg8b7+Lvi1tvvANACcSygE0LogYw2B
BgdeAyCYWmDBeiWy+uLNUChKcUYoyBdpA/ZJBnzywThLpSfAhm+HzyJemz5NkiaW
STMI7OCMtYBRn6sQgHkNveBGB/bS7TT6N49ZCNjVydVl0ojtzjpfJx2st7rXkFvu
Y/Byi3pp/Dbf4q2I1bzT25IlyoSTlG5L2dEqKg7rj+6M/cfM8A46BM/6EzrWLJSS
tvOh17c/O7SqzodQUJrcwaKcXR5mQLP+5sElLqueOlxakVOccgaAMYmGdbH5Mo7M
FJOrpRRsSpuLbUz6Bo6Uqg1inHOFAcn90d6fvDfrP3Ubnzo2ZWDgsvhWpfFDxKgc
ChCStVNNDVqpTllN+t+OB3asiQCOEwMNMxaLGN3odAmY/Jy9rLa/lG9eaqytJLJ0
sDQQq2iJ1pSTGDY+EAfFeexA+kJqXLEEDAx4wEdWZldk0rO2sr/Oj9S7fsFGPZSM
9n0ARMHRYQLkBwDS5q6H+NK944muFY6ULWGs16KCur/+lrAfT1ZotNixu8Xi5kyH
QIMOnlQ+7k/4NgM/ODEZN9458GPVGyQRWiWyiUq7bivOvxyksAm6oNJRQCgF8H3o
TfeuZQxMnmDtiJ5sODFDtfZIyDMJwi/xMCF90KnFFAy6IzGGflzFH3o/WuxMR2We
gX9ad4PUBZEDhUadR2mcs47qXhoVQO6OOO4m/0hYmPQR6nxLLCHos+/GdwHJWGBK
ajLMdul0Q0PiBSfUtRFaofXZ8gbZ+gXhEBhhOgr3UjQdf3j8UFtI37edpb8u+XV3
eSklup0Z7kOGkVTxv+wtAx+JJ7P29YHGjEg4rvi8zI7a1AzD7J9SyeNMzcIp1OHr
D8xAGt+qHE+K81HyM6w+3EgQl2MvgDBGSdTwhKHvzhWulUwc4+a08QSODdzj1U8s
ZkZVzbFBSap7kosCuKcx+MYEdLdCtkQ9c66KkQ/nf0gUqVg7C9yz6dqVbGDGipvj
Ksx2kjfMcaGaxYX6cZp7EjBDieQ23CItOZ8CDE7kGZ0e9jvNc3UGfwLbyn4hK9XX
twUf0fVw1/If9ym6wFbL5AyWnOFb9FvIhTfQFFtRkj+MIAFXyTSs0qfW6mIKtUkE
CNbDIPL+csI2wbib5JVMiHqtNhOJLhIsPXtWHHEcUiAwXvWRBLv3Uwfedroq3cQW
+6WXOLYxIsr9t/nVcQEToszHsD3iFDrIhRJswrJlBOWN2Wltvii+Gf4/vIC2oRAk
+c7JMDgdjkMe+9RhfA36y/F1fIqRB1n6qADpRShJRw78qSe2/dP+Fjel9fjoDLlv
hepxjrvJU5Ue/DiZU11A2hi3tuIhr4ZAk2cfPUqGYCwsmnDh1ZOeoCXOUDtJias6
BrDsURJBa3rt6jssCZUbiUujRKd2f3d/9QKQ7jsxYQWhUtl2f/EY8sO5t74eBx5u
4E6BKkpgt4orcyDrnxolc8CFpXK21gyrFQ0LyLQp7m0=
`protect END_PROTECTED
