`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxNS5uFo36NulTdAhjZVuGDLbXUjtjtr6uu4Ke/coe5DpMSyvATdL0/neQ/xnImp
6ATN/3e7BV0Sjj40oJMX9MKJemH3lbE9l2cxzQ5M6pvtcWPxGe5zmsvmB2xBgcW6
wg70zs3//g9GV7FFh6k1baf73YNThiIcvBZW7vlIO+GI4RBkZrDLY0SeIVfw9ela
MewPvDOIgfe9Y5lqtW6aBMaoA+h5j2FZNyQ5Y7o4r6kyEyaayBnslzCEkquhfT+M
i4RkdWCrHiVn4x4SIFoVBHUit6/zwvJjOKmQHxfm5QbEY2PhxQozdDEkEa5k3efu
U39AIrHCOjOG4gy/GJ2DJOxi1U2N+k5yt81WcuYYlQZ/ws2QRPdVQmGEjsaRI+4q
Ktn8vmDU9dRzFxAhbdsMtNBQ9/vGQsBIVE8gIrj+fYC1EzA2ggAG4f1r+X3x1Uw4
a0GtV5s4Qod8ocCayplbDjB9tc5m0MIIXj5cailRnRY7R83uoj+hl4UStDqeiUiS
o1JMZztJFJU22oCX73glshT/JXkvjnrqqii2Bc828N05B/BB8XZb83bdQAm3Uk5F
w4hd6VxBW0x+MSNW7DVsC0cWDPfj4rTrrsbIavpSDHkqqKB6BYbFr6nf5khMbBCk
k+Q3SARx7in6yF12fow5KghdQJjO8xUo3zoWeQEmk7pvOm05ym1ofWVI0/A9cdac
pS7GQ0LVt2OQGsJX1jj3iFy25GS3rRYx9MDmhJE5nbkQaeuMJH10q+7UfpM0EBG7
35+6tUE1re+bby2VRZZM+lL2VwFKa729KVJIGOl0/N6HyKz4PkKE1Ol9kO8q3Wcb
SNayFoI6/xOiIoxaTmowH23c7/PLW3jaLILNV+Y5KM6AZk7V568CWksehQQ/y6MK
4hSnX/RovzKA/ag2C9qP+G0pObJEGMORkx+Gzv3dHUF+BGHlaHwWpA8gqb6FBxzB
0tjhS7JlZkwADd34UgoksqsVV1hiOsHvfyUaDTz9/xQCWqLnD3QZj2rpHZY/QAmk
8t357vuym3FkjD+nBISlyvsp8og2UQ6Hsz4uAJGup5AR+ITtxsqNFqHkSDX1yVfn
0285M3pelY5HnpK9donR3CN+koFvCIcDp2TJGukPWB4SSKTghGkCQD5UmAG4eEfE
o3IVL5hLndAZLecGg+NvsRhnRxnjUgbpkibKwqH9fJCxeudXKRA/bFCtnU8uZPvl
rhjbIqDtm8qeI3UmKs/eJRO0JUBkDsyQfOiObujr+1CvRbKiU7FVDjgjoOGSG/B9
5Y8IRx5DhnOB6oDvAxHhk5+TQ82lcHjS644zFCWuGZ1gX2VHv591d9NarBkHv7cT
j8af6OjgtI/m5vr1WIPpXcq5/694c41sH7h9u/Q0YuRNUUG1gL/f/+iHlyu5VfOk
Qe064t/76s4cF0lr0Caz8iQ4m9CrxDkAmajkmvMmVQLF4UhjueuQkaYMv6aeRlxe
tDImoe324ctWj1dk8pgBoOxJW/+i1fIV7L8DSTiK6YbJv5xiUah1VKy773zIXVd8
KThN3RQIPMdxQW+6R5PhkMBwQ507CuHufoPvV74QlYM28BQ54ySt8bvtrjNJhhJT
hCNudfeXIj5sL1bskoixhnR77eIRdNcg1fR8LTOcu+eWG1TF5l1G5xzBIU7qJavD
Moeem75vORIlJiPOY+sD9yLZ/4sB/8z5UQ5tDGz9eo7OsQ5nD65f2lUPYaeC/FuV
EP6D0czIOy6WMQF2QdgUPsB2XLDK2Le6pBccaBBwzET9pizwFwbCupBkn5FO9RQ9
i3DME6pGHJ0H95CuO5U2LuL/ij6HlAXKuiDOugIQ9nqBOc6EciSBYedwgrNATXpp
BW/aMBAI9MnKIwzdr/dJ/nWXEGkPwMNWHIidq7oHj40sb0oB4q9lGI2PMCmykXBl
Xqu4flxN9wPGgg4MMicuCUfP6Sh9JZZqqfYcNFXeWIvanBVcWOmP800fdLBtWl5q
V6bzYRIlcADBKqGYAd+21IwdV2AO6uSUoKIMxecSmJk/Er4b/j6H77RkhKb/HZzN
YDgA/x/jdWxRNlRZSlEw+zxk58xSsRJ2w/RuvrVMm3npabOecdY/o/pJj1yulKHy
ks21Q2ajRGXE9Mt+Wvcykj7lngQsJkEdK2WX5Uov6Aq1b+GBigR9NKfCnvckVwWu
GdyDM/L7oVQwx7Ublf/4eIuhiRnkJCfJ9rApbA209YfwXNkd7azsOd/dRV/49sal
mkHa9eKtY3JdIDqTzBMCQI0zlQsUFiOEKtAk1KMZ2b3PXxGu+LrzJ3M7Sx1wAAyK
Oka/UxLwJHWOxrjeLELsV2e81p6v1GFq/7nonhehLqJBNRZPLWicGmAFl4PozRva
JjdagrEnG/0Cp0tEQcZ4bfAAGRnpb6OnHtrSt8x0i0dl1fFq/nxPFD2p+t1qiGcN
zo3vr56uIauAyJAurfOP3HPbXoWGVFFdjewFtD20LlU9i0UiKyiQVr5dlf4IMZaM
72mwR0aTWkFJeRaDrbb/3wCRdbZHXmsgu5sS20+4ZR1dnAUuN65HICdlxX+Gy8PU
pxaMoiGBmn6DNnIt7MybAlAtdrGgWh70qVJ/njlO7lk0ACX0tt+AlaHobb9iMjHx
vY+kD2MlpWCNxYZSoQT8Ef3iXrcIuoT+cyOkt6+gZ1pwF/sHm0s+pz6NlvyIq34q
TOWgdQCUuLqHimz1yAuNIBbgqSCgEhfCdMnZibeARaukWNLnuvlun07aDFJaMiRd
HMCbUmVEK6qv8gN9QuTAakocHFQqvtjyVQrsvjvYV94WWAKl83qOF/XvVtI3X89R
JLrB5NT3sHPRvLz2zGv7yTT9pMde98Ogm4YXA1DQFTR/9sNLJ/DTCAr9TN2FrdO+
0GRYEpMrJG0vm+2UEJH48DxJPnpr6ZqBonD6wLzjPJf7cJn5Qj4Jbcf4v87aYazl
nqGCLH0YRr/ebLNVjk6dN2rAodCbfLUW0cIGmn8fmXnmFZab3SYdaamaOMWu5WPV
SS4jo2VJ+G8DJrxB6nxFkNZ3gUmyKHXSoMFt9FVJoFLyWW0E9YCgY70MRTVZGjsq
sgt4BVRJzKjDeVW7ZEBdjpsNYoy5tZVSP7QfECOQLVBdgIzvbzDqMoqlXNcV6Odg
WMJwEdLj47cPuaUWM3b8tQcVtjOb7hAoVU+viZcycGodb7Igq3Bt9NNx5V/l0mbV
acKgOS1gHXbLSH491nboJLzemcizfrxQW6TeajVEqBmNjUO1RN2MJ34Otd1xrvNM
UEr+9zAeeMgY8SvHFw1hgYZJnZK3VYmaQ3WGy2g4O28yjKSh4h++zZ89eZjoQ60a
julIg61/vs697w4tAofQdPhOzEALBYIMugJ+ugpuDKT8dhVSV02lXZljX+53rj9+
Zv8g92jFqMPy2kLkqFZqhwxGLbrhpOVK8tbEZaZrmbhURCefhiH/VueT3KpdWuqs
qwNf+z36Ut1iWEwKGUdA+6Nf8ozwW+2uqI0LbC8VTqkDrxRRLxDpT+4xcdtJWDic
3cbAs8AkRWUelwWGCezFkT6t3tmhT+yEKWO4D6v6e9R++QbmKO8qThhfHXMHBuk9
xLt2gtK2mf4WRadANPafVn/Bxo+30LD1FEortq5c4LIl3ae3FQsmX4mLjdu2MRM/
kw7cijXteIshuKvCjQ8k0MFa6IOFzk0YJDMnfFQLHzI1zqDICO6sS3eJxi4Tm0m1
lXunhfWhv1OCq+wOk2pmyWFnBjBDn9qPioVcJNRsXsDfT2NpVuKJIaLNEvHSC1l1
RdYsKALvc+APq13fC2qn+mp5uAjwj7qI4cUEr825nhZHeksl5FYuGwaKo6C14ySh
e8DXQY+1SYRY6pzqzg6iGF09IyGszuQgApxy2Q1bkI1V/1YyRWGYRcovpbsk+BwW
UWp3zSV18MyFu53w14eiTHjvFHjjansYnL15BeVWAQMjZTv9p0aJ3tqjAD1q+M5y
spCI3Fr2NShM1g+XsdFHP6/w0K92B04MlOdYEFgaZw9Z7AkyF873Hp4oZ83mctcW
mar8Aa9ECv+tzRvtMemEtFScXVOcjmuEKTBoJ1+WIV9sU9nkjSwreaV38vljUD1c
K6wPBdBGraMitt1wfGcpsSLfN1xIspIPIH/bQKHlQ0P+MsFKZPzZsuKCTlvESx9F
B/JiokNWY9BgI5br0ABEkKedX7Tr2VX4Lka0KbWDvik9nqNxOuBZB3wuYy+VdjRD
62/ixPj8uWWmoGfl5wig57+/Dxsv1EwcCpBo/SotH8oKvZUAN9BkNfVUnpYUykAw
/vLOxnxMvTPGMR9wkHchJOB+8Hv9TFuo0TdFxEVLnmOgDeONTY9RcX4bnoZAG45K
HUs8zB750FoShgE/zNioHfoiMr9rKWlNipGAO6hcX97c3e4JShUUIt7dOBxulamd
/zeUk/5i4zYmxtzqwjWEBWhe4YGLuhT8QOmagLZfWofsXsEnR0VJblRMXBOhvbuP
cMK6Bo9xwHebQFAhdDnqb3rNcc6Vik1F+A4f/IpZD5l3QHji+NFf5rAD1HEDpglQ
oDetAalq9zqAWnUxoOlMa1SYlZ3ZWPfiyNYusNSfuIOlgJ7a1EbNUefo9WbD5kY/
8oWIdHUCnOrg0t0iP/fLHJAxwifRqkKAHFa5seeGzSxw1YkJum/VxjtDJQ/o5mKw
lnG9q64EEeZOK5BS/E+J8EZPn7FuKswUSxP9Ck7uhmKiXcBOxgSTHdHFuwq0479f
drha89RjIsH2B7JD7hg26KqOPk+bMT/Ttp30uOkvQEtMhBMLc+DwvJLlfaIIz8IG
SPjCSCobgcU5QPAHH7izijUSJdFMXeo8nORbOWiFG+FT9OBeQ6XDUogBWsH7AqoS
NO5uk05GfPAS/6uefbAsKeOG8BK6ca9xwcxmZsKcSHlNClnjTZJ+e8DIy3JzeGML
NTUVaqoiZWdCQnIfmOLPpBqaQiAWs/AjljJd064PZ3ms2QHuohxaz2gPpUndZNOP
yj1WRheH72yTgJFd5gXh2jMlCieyuwe1kcQyRiV27Qsvmxxr+AQCd5ZCXCn9vCsC
xikeuTuEsVD7nK+xWFXTz19d9w6Hxw8oMJY5hIz3+zhCiKULR/USFnSyzkUpaSEp
eIzFnsUt3aPQxaPzHqmkeIdcTxQ5fNO+bGOJVus+jm9nq/2fgmGxOT0JPP5HmwGy
+5o5pHCexf0/cUDpnkUDZXjBPXXLexE0Nya/SIntJfQk+L+csJ/lUN0OifL2ytSj
gl1xfe/7aO7iSdQJAgUu68sA1lJGRzkFZi4NCjHE9PjCliTH0ZCyr1Ld1JfSL7rT
oOM80LpDkaDzIRrMPjvLEY8QZyutUiY0qYr0bGskBI6G4NI1nXS2uZzyVt0peZ+6
SlN+egVdJI29c/TggaUvDwYiFNhKoF3z7UoyxXcwthVef6kZZPMjb8e5y0C1GLcI
F4yvfVWrP/6v0Eq4J7Eh1NXdZijePgXZuNcgU8k2rHpCazZpnsITxXbgXhE0gC+W
21Adhz48hW0x1oTNuhIf5IQllXHf6kX1pjT9SVas5AWuGk2K6tSgJEaKbS9l2oaQ
TwS4KVhl0LQpaVRcbjXAjRFkCwq2vOr0qppC0+YyRSMwn8do8v9j/QdZ+1WRKdI0
u8EQdqQ7kTqtzXESqO0ZM4kAyJSTiUW3B3/rdYQTwzoBj0JMKcPetjpbCSVI8/+B
VOsK8ZzC1KRm+3I2As/5sSXWgssgeMIfmYnTq8hEKgdAmj02gYO+fOOcOmFEihVZ
jr3e3lXnYy244PGB/hEIbfu5aIvrqsRdl5GcAuxA2MwTUYzzG7cR/on+mdYhIvLZ
zCWf0BWV//EjxOo35Tf4QIwAYiqsWce6TFv6+uRK7xCIbHgMKoJLdJMX9wwADkZL
vcRFuPxrqN1cDhUw1EYnaafkJrfSqZp4FEGMYLZLuS3DNRtw9xuM5HpZ+iY33j97
aqrj0RfDxJSSClyD3b7rFWFYs+/l6n7snmw+9MJOFFaeKsboUNoCI0kckS0IXd5E
jbfzaQQEaG4qciNRe3/rKQBKePvgAdAUlJiqUb/H/IlG/lgc4bhG5ppghJtHmz2P
eTS3HqRJ3q64I/TwxKX+tJhCkrax/mWEywzld8OfFZ6ntrOFKGRmSNjt5/tvk5eD
WFZA8aZElA46FJ/GaRI9/gfhzp0jjew0h5Ph6cdD/4l627rtIn11OGCdSgdaNAzZ
bgOcz2Dx37LXidyV2GSEg8TbIf7cT5hX8PuA9oeUOev18PkEqrU6WnGNbJq3qYP4
2p5mRI2X5YbyCj/XKn3gpROlWt5rr5M1Ed60rXOnXSjGIDGB6nquiYuaMwAEnkql
fXISEYWIFER1F7HwKHDSF1TvLdvceeqFhzVw8fD8ux3n7VF5mqKzNe6sDZEJuyQj
cnSus4qWzTFuBzS9/hMsSei+UhAaMo+8BqpMwNHVWDfCjFGT8XzDKxNfCUmPwxRs
WEJt+APxPpqn4CIg8P67Csu0eMHWgpgZrc82ZMbu8e4a8RIu315n/y2rTF0ahrEi
x8z7cPy5YmoONuJLU3SXnqZCAxUJsgom9PWwEJ9BeocdjIzP/Ie5dR/N1aJgMIov
2FQ3PD2ro62vKKB51RyjcoDHXrkdhAGI+ZMn2peOa2c/9wgkDxUvBXsAWVy9cEXY
UJHRoZIiJUWH3xEmksz0o3zfni+tZPYk0tndQarQCDIc4QjmSN67Cl57BsSWJi8o
aHSnWohwUTkukJT/BTTMPyvNBqX8qnwMDa6MbaQiQAu/BRlb2yfpfLxGMnk6c6nd
SRVE6CaOH8TYcOAI6m1PFVI/0YRGRRvLWR0PRaqQrj5Y7nRY8KbCyFAnp2baG3J4
338N9AvQ0GgZlGQk/E2beS40i90Rok4lxgFIMQ0g/ivnU9sidwJM4mJBV1dIRZA9
42prY7LOYDTmyUbkKbAG4JvTaKaHLR5EUF+P3tHd3ZAFnMkUQyBbH4Y62+Hq0tT6
t2VMjbdpHRjoP77zOC0bdrn8ZS/b41YBpu/JBJ4c6WdZsbVLBVf/SiCVvTRQBSWS
T0+oMGf3wixobcCr0kSWNowjG5nx6v5RW2jnwpgBd7KQdol4PECeCu8Nyy2ZlMgb
7+XnLYLZFsaomBbvOMQ1npEnIXvXuXE6TpRrFztBrq5pzWjkn+7FXM7krCTCLpMF
E0LkWAvhW6ff67q8dPk//ENdzrYdD6oxfpraLjF5bNneaBJekb8Tvj/mfoXTmAjJ
f/zKCyl7ZXxGiFxn6DHqK9oTcM7OI9TR0eblj6MPxx0ao+kd+7IKG1EEhS9+cw9c
31g5SxgsefwF4mATpVPM1r7A1NChRJ+XDQDXhJDoqFnlLJIGwFFAOcen5YeprHKq
HBE7uvXzgCAgNs7aYVMPugridh3MS6CE+Dw6YrnMCvjiJb+gtvlUcMY2fR8GLfJP
XZWGYtzLzmHfnQTMESBodPf1PP4NYE0Cl1Lzdm6S2DlYR9kXs8CrwXRwWd76pSO2
LR1BpDJDWABr+c5T92nBLJgv4Np86vfIvzljWIgcwHo167zQ9uaywf7eEUgV3AFP
QhNIY3bybWrrj43pG4PLdVPHkldCMDFwScJsVUeiYGD/kY+t1Hkpvvp609SFUqlM
F4Mzn474bee9Adccm1x5ULBQVxcGcR+d5IfD+LC9URcPHoKSmL3DE9sSC7jGBjWo
+1nawSji45zFsaFygvwe2aDcQsfgC9mWrg7hkaRoiXE3taCOlsPRmSVhqTQ6sD4b
/DZvNpkkSlJYeNCJFyoGjc6PodHwjbMnbobYSNXmaMpeEGdcCb0kID9SKFibLruy
Ha4xFbLZMA7NJXQzsgZsX09QWg7QFGGodt1Ys1yJs8KYogw2dsHL5E90CuUxvwb3
tKOnMeo0YrTVNKbU25CEp5xfcJZUeHdz9tJVpKDgyHFYi5zcM4oUqd26wTrHA5Ih
j6b20A4Q2KXy3IiwsmwN4p00TFOK61TTFWnSfMbCsl7gtcprwn3g9GUnQ3oVTrPI
9cgZCi3qIER0x68ZQMbQbuqY2midUTBKz8tiYHXmcX5mzlo4IhnLmL88+6jSbRXt
WsSuMuH2Ubphj0HudIS2u5iBn6j590tnKzOq/CjF4a3FNEls3wr+Y6L+CueYJbs0
kSt86c0qYaIpFkvDan/wD0wrjEPNLinXACFpQ/5aV5G2+LqU8KrkrZJQQdDocmsE
1yylM1XxxgGvJewYiTK1ZkX8x2ZUBuMh3a2Ta/2hZsSgvAWq7tDFPNkOF9wpLIUv
hKM37Hf/r/sFD1QK9I4iLOHaZAtrtIqsl5vS2b2zRknueQ3DqPFnqXpn3zhLAgTt
7BAryaF/kIANvPRVL1ft17g9BhG+Ew2so+42xtcZs3H2G3eSGsRHBrjVD0ZJ/gZx
y6dpQvBmmp9toyIE+mortTQB2HpLGzQZJPBzOVjPjYATCoCG2IOdMum2a0MVpOS1
2mrKTJTW6CNW08VCI+YbgQ0xJZ4K2HV7Oh1rVjkF//dpAaeiwAz4p8zZLESvbrmS
C+xzWybvgz0+bLu3wkReb7Fxli3Mmiuc1JhnPZGSj+GqbnbnijBuTFSPegS/G5gA
BZMs6PhR+HW4QKmQEgywpiPjqL+ydaqb83gHD9TIvwxBUwZ59Pzb1ikKjKLYgjkp
ZqSIxaUfvNPqs+R6wPyaGvGDRyWG4mjDw9WepLAey9dQygqs4eg2fVpNCGz6zKyt
9mENP2/SP21UkE9mhw6LQeZ+Eg9mCI0n8/aodgbdTz1dHHtITSEScljnA6g3GEj0
Ggm4g0impnTxgpmB+/rTxGd4Zqt3cNY3SxI1H1cz4XqjjlvOYxFS3rHB75eCr5LP
yJwbw/KmcLcRYsLhMJC1GPidmdLbQ8BufFXSZJfO9BJ6lxjUW+aaku1X/QFqB7Vy
SUmu/g6Mkc1UyJYNjkgG9PQ2ynhU2OPxr0bDL4JcxDXiHz69MZEY5A+M6g5VMW1e
ONVQwV7xWRWdfUWAAZXZGmWUW2NYzG4o3GpJee+N3XSyScFUvboc7zW8rWbKz5cJ
yeILZPIWKOpdBlTP6wcwOkH8gKn575bHQaUL8RLa7Fbqd/2L8fPmcGWaq2C3+G4Y
S+0E1X8iOp6NtY6OcuUjoD7oACnm7a6n8MIppdTcQuqRoZyoMHitKIyqrnphZK9N
H2E/f7rogkCmuk4hdWxJ3Xegz/pGDmS2Jp4wAr/X6AtrexLtXbhRcIaQrlT6MzZW
aa4euuXPFUAzrslXdQEYhS6XbeCKvGyeHvYFFNKKV5b8oTSb1YrsP7G/CX7LDBTi
UUEi5Kt9AYNgTZ0OexQfeyxZTte2uhuOAJoN9GJfxljQezP+XDRcbksDf53XvUDR
/0TW8qzHYb38n+I8V+QrZIwcIEW3rDBORAdm6LumyMH0GXgYnPvP0JOkNM8koaE5
t/Md82wtQDnLSGQaWVtLE0dAtYEb8iXNt13ON7cjzknRLtgK9zjPFlwccqLsK+lW
wU837wtwvFsDxF8dIhDFYtYSkyeTIoz3D5++smVtTwklsxtxEBjP2LKJ1T5x3VRN
6hyd9gJN5hYHjJMtfUjkbu9ZrvDF+MwoMjFAPB+624FYKn7SHRXFLs1taILCHFwn
8SNDrAfimWYPy8M/tcla4f/VOZGV2hzE5D39fsxAGSWsT2JU9PdWNiasKU1uTtbP
fa1P98A1dzzR2rS+WELihGYMr56/9fRItX+QgaHqVXBm/feDqCGBWwT2Vfe5do2y
9aEyguwYx3DoEYUTaUwt+35s8crZGy+NDUjofMaq10r5KKpTihPQp75MGBgeWYJc
o6+y5gdtSD3LJyBPHZgDzT9sFwb2Baiq0t6zTumMrLpsOgN9QOKvhL9q/7aFJb5w
rZgdGsRoTCQvOAh2ZCONQsbhmpOxq+gYhZTonj7Kkzb1nfRGFeSW7CiqGCA9hgWx
U+Y2lKLABlWRJviZ9wPzQ+bZR0Oj7WCve4dNcFQTStZ845l+aG22ncpme5V4lANH
BHhmVDjB5TjpmF12ZapkkIrmWXBJm0g4reSjVi6hxTN3Irj8fJcgdSUKZknPCJzx
/TN1t5NKO/dFVWn+xpMxa779nYuIFDjKBTk2b/DyGjScNXrGkiHuG4jeL1w1vwrA
V3KAxWtqWkNLagml06J5rPyZCB9QRSrx0aP4mKZQ1fOpYtnao/jtm5/2pgoVZM2D
bZ8HhiK7P0W4WIAqtvF/lcQ4pou9SAFQQ72O3v88G1rnNQ6QUXDYJEoghKdTacbL
L3fb6huBdt9hwPPc2WOVn/DgqMj39OfTP2vGBLUW/RZ3vw/YGZEWwUkQ/bERpN6m
rCFnUYSsug16r9cNbI895qta7hS7pNEiprWwNrMeiR8a6Vqq85AbNQLfVVIqBOK7
u+9FnyDfrTSlLPWKUMV9phUq/0/Nx76MhwxD4UiIvgyVUbo1/rpGaxPYD7WiGZeX
JTc08Hdbh5l4o63aPytaNy84BxhiZd1XeVoNvmXF5dCiJ4XW6LD6smkNzq04Zp38
exYLliKC1cbXRAgRQBvp0MicVBQG9x2HHfU26s+XRWVqpUlC2sKbTwmU7QZ2a3mf
6/vKvyyq/PBtKJogedECT+KID9cgDYYOTtMC7SOfutufzwyc1NMrlEP3ufUpa0ZR
BwfNUqEzT0WWR2vE7KjOiOX1ZFYiJQt1KEEwJKidKuCG0xrUEW7iJB4/K6rlSXjq
lOevUTOBsagKG8B7nzXO1gusRu9H4tWzNiFmilIXiNwACcBxC0cdxS4afHrySYvo
geqV8VSozPlatOBzG7r483rfOngLIYCQB/21zHN4K2J+0eWKOo34K+/EA8vk5R/9
oFBmc38HTkrHMjTwG/xHPuQg5FUCtds+bHMw+yy41U3RuN6YOgoecz6ZNazTzovu
W0052JRyciBoygNUftJPdRhBmDa8v2NcAf5fOIozm/yaBaoma6FgoBwyHAqGMTYY
h0GG4KpC3ih4nm4cXtZjn/FlHYF7Wa9EcAqu6PiuAWKCIEEcuFviNTN3Zl+UkC71
AFJKGI+0zyY2yFd9356HWV4VpVNj3fqolUCMIJE87Obnol9lvGoJutVkgmXcrQ+n
WlBsblbqCDiFTUy0ejSHATLCP/Sn7vcxlPJn4ogGCITKK33wuhG1Pi8jy1kP/Cod
r8227QuHHHfAC+NGr2VNCcx9aM0Fn2tVn11+lIbkV7L8jOwRXqz760uYgH68UhwD
vqi+qJunakHbwNfiEFmiGebh07XKRdwLFFLuHrBiwsWfd+OUEx9H1OmEp4ZO+dc6
ctn78kjQUT9+Yb+toFdh2K0lz5GUFFMvnBcADMDPMiggVQ/NlGz8ATFyECnOH42A
VQlIycxGFHFUoUZLBkfV0OyxZaOSIWfupVS5kTRg/1icnm1WtOzeoBf8j+TWtyGp
i+pnjr4FCp+S8PJb/WgOQAG8aw5aFcL+HgVgLanEDzHy9gnee9Jhegios0tO9LaP
IQLThTCiuHsQ9ATidZperd3IuwNO9Qtlbf64zZlLInJW9zG0dk6kQj+LuyNito38
U+EYw9y9a+boa4zsbfGRmrChBVuPOrzYJ4pM6JQLKdDu7qKH8GWDcflhIAzqzYGx
pEeG5be/zOr+UAYnfj18q9WQnhcXL+jgfmWDEgjoL7VmzfzdWkDRagY9CR3YKZk0
MOP3K8lxugiitaqpYZw+K9d6QXslY8mbdFmBAnd7j+Yvib6KFgPExaPKx054Sbgv
P7R84aJcHIkzVvEJ9KDUSnaGCLzJdd83Ye8Md4Jex/1NATCZ/iTELDRDenXsueFw
/02fWXFymVYOBKWOK8OUfMIdVUN3scGmhpc3E31YPnrmPu6HgS/iun4gfkxYzPQU
2Yq4Jc8RWO9cBrPZ30Oc8E8jLUdkikxuTnxsNipKbk0VNVmhz6B6753/gVJQ05Li
xzR0ASSsfH/q7GnWVuJD7kRJim1G+AT9akDWktzIbvD0REv4quGaYQpoyw7B0ca4
Z/wqDE6TP1FXX9l2mug5wzxWBJSsjYDuoSY9GAcOSoOiQiuFyZptpQ65AbeI1Edn
OK0E+UifeKto/1RTg/JFvwE0/Gtj9HWvR1PtqLlDe2gDQG4gkVv7+qGhO0GoLO5z
dstQc4RyvoYmlmo9oJ0AsS5acopGeoj0SvEq2f97UjTYvdYqRTia+dHZSdTGDMY/
UwKvCqHHdaKODu65xQB/tZxXUicB19pjG0xSOo/eTeyiO9Wt2kRwhSgQmiZLi35h
lCNL1X47swE6f9iDW1uQBvfmkSOvMMEwfcc0w5bbKeC7fJ1Rs8PWFwmel5GwHV51
T2Rzv+N3Iag9e4oW8VI3NvQEKdDH2nyy8pQxGYJsdkOhTWYu9qz8+qiGQTD3Wt2Q
PCgR3q4NL+UbXDWnPWJ85FoBYZ0rKStMuMoz3xhCizCMjvTlbS3F0e8PltmcODyE
zkBaUrJnFpnO68lWMNxOrAvsvnzxnZAHy87AV5lZhbLncaCeLBHxGZmLA3/jMvcF
+RUJWxtZuzPPNNn21OTzxph1hjbaa6J5/1+njS9dkaHDG4tiWZylwDmOEj0TfNXN
eRCSv7LB1Jk/s/70ue/iRtIj66n1Jv+h78RxypKfTmfhqouoN/iqpcnWArb0PXZZ
C/QD7oG081/qVdyt3MgCt1KvX0o6N4LsqgwNMwGlNsVZ8ndoR1Nu/z1/wQypbbFA
wJBp0qBsaLukvU2fAJO2LuYuqTAVgta88u7ampQ+vUKldFtmLpO6XJaFXju1bAVJ
3acxQkQpu0Ru3lTMuHPMGeaNpt0WCZLNK1mK5eUe854yeBGen+TTjIANPgrAFCWS
S/tVhTFGuNtPCp/SjVl6SMiexQ/HHvzV32mHK41AJv1KMfzOafyw11ewTig3Sk+2
vjNpDBp9IDxdSKJ+5I630hbut1Llt4zQ6odc24UVGmBiBGvRgevv1KsIBbWUHtv8
+IaMdwtIKZIGG/QqXAegJ3FaGIATLgzi/YiNXTnIjetiYcZ6aTovFikqiyqF3ZDa
IHA+HqcagdyiakyaRp2LWxb8N3+tjeOTgQpJkzo5YAJlyqOkVuVMkkMPyPo8sTFN
TyPOWlpMGn7BO5BSmMRFmqdyXSAAIaiCYhdcz2ZtpCSa+Po++BcXRgcyKirWgQ5i
L5UXwGUNiajNbbm15ZzjOuFpdeD4v6iUIOv6xlHhiJM94vrwt986lECOk6dO/usI
BH/rHYvqy2q3xUguogPzFCgSQjnSAb3VWcO8ChXTce7r9fa8iqSdZuLw9Xaw4bvO
R9R2rrAS37osgVMURxD1EdWi8xBIfkf5q7T4iudpv2U8Pa4ASgyBo+/Q3zqAl7hN
KXZKiCx3xiwgLzlIrVLiE6IC7A7d4sX2J0Egv+TWiRVIXsplQX63hvExGrRsyBPc
QY73wwcOaRWdsN6nC5SRuJL+8IKmBuQwrJk4e92Ed4chwysw/lX/BCC6fIX30mUe
S5RL/wuIWuOXiw6XHzKvOvhrzI1Yet3e7/C53R3JrqpYXO/CKkdal6mPD5U1CJv1
KvzqZK9Xl5AZtzhmZ5hkVA2w7JhYztEN9Ptbv6CreEeR/byVz2SJfFUf5K+2Dy07
bBWMKgb54I9pO16XZmePHxMMGB6CbIvgqXElx0B935GX31sCbiRcWymCSO3k2ir9
G3DgI/dPoAfbr6mAXyBMZp7vFwW1ssVzL4ENOlBrsboC8CcpzEJUXLHQvSyXFuc+
lezaFvzcYKyS0Mg5QTmri1qmZzJr24L7q2PFXLU6ScSYFCdTWAeGhOfm6Y78LXd7
sR1Kvx9eX4wmJACHh8opxnHmG8PgVTq5E/znRgCuVNqUPnx702f4qidnDFi6F0eg
s0Bezj4RC7/sYi927LGx5PqZu2RpeI2dnZkhXdVXfpgb0BL2vfC7Of1DjCtIezlh
+vFOjYa6BP4gR1gwArr6shmoEQvJgL1PsCEAX70FTFJpY8zyVYdWna4PuS5OsBRW
5Vqa2/FY4mmRddj/n7RZIg0kHO8f/42WO84mm3KhVuOgauToV8+G9mQnLJOoX0xV
vjcqYM3ePJrng3PVDL2nwaNmND5LaKlqcFV99eAV9Kf/GWD325CTHPsk4cKEWz/g
WmmEGSU7zyMWI2IjycNhHfivrp3KLnvTgxeMxsNitoJQgXRESZx8JmTexsF0PFMl
PSGSTf+NcMsuKHA49u2HyLJ20l2aRmaGpz62gmdSmK6rzLMns603ovvri7y2bxbw
IeXSepiYrcKucuE+gCx32xC3lrIWY7j/ye7CjeXX5a9k9BhEHCKLjs8NTc7k/nsU
mYDFcxBY9vXDjzyJFhmNJ2beBGFSPVtW08advWmxDcGRQ/BN/fWp4FB8BWTJVC8L
CQ9WCv81yLsy8jmKewG71CDxAcsQEhRIvZ0G9dqpMndXU0Nw9jv57I7IFvUXZFg0
9Fk33Oq4b1kn6cXowt/s/8IQ0viNhiOvJFNn9kVM0HdAzL4/6bRBporerMA47ptp
iWscjjwKadUih0qWmNQObPZXWa2pKKISoFAPb3DZtqiEhRJ1ybH4ybpmdp8PbuQd
UUoPV2BCqM005a0+xOy68OZ1rFX9JQoXjR88j7NC2sHAshLrBQN75hsYVp4UxrWf
iJZ8+29+zYh/6IqXk95MUj5hB8UwhbDTCY1PURuSIut8DyPJ0YyIcIS5fvIRRNBP
PZvJJkCnmWR9zp4ZUej+tcrhDsXZ1xaaWD6u3RaRNOVavbOW9U7hbKn0DpRGdcNi
9JcFTo90EqmSepu1BuH/cvq5Y3Qo5pOueupIt50x3P5UQ+wa0gHy/EtHTy17R3OO
94UMZr/w2+V028JARJjzwWHVo8k/OsWmnEhORCDrPD9eoQfc75IANtLCNJkw+ARe
r7kk4JBAYFiBjH9l72CXqxHL2xG8EiNiJfdS+WrrN7EC1ds0saY71hz3kk8bsCjW
AeShuDswN2rh+0iJeNb3sJNgfxpZug8iaa6zEztmQs6P5COmSpXKvJJcHAEf29yD
`protect END_PROTECTED
