`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
claEjYPUl8v21MJGw9f0hL+PdmmoPK+My796EIu9Ewnx3ns5hhhVa8W6lsAw/QFw
9J1MJvSnxhp9HromiA2l4qxcacmmAlZTsvsDlPwps6fS4GqrJSnETivV9ocHxMcw
BqsoFvVTn++31kg8K4GYavStXcL6JvqKhtzR1x6usayK09kSsH3+dFoj0DoiUz6P
N2H26Yy5+M3DMRwxrRgoREN5HWHXJYmCgtRYjZ3A3xWvglo+p9gCBu9J8cqYLsR7
QHYdXwcC/WjrAvYNsflQoXf75wWObp2RgzsmHJyWnbQaP66Gca3zEeAaWI/+5ypD
koDOWQfKI9QNLNYIeWya0wjZisCXEK1HG6s/dVEiXzg3qb4icm+r2KkVNWht9FvU
nYF2TS8y9IcvsWFlqt9kp+aLnd8Tuw+jsx1EuL4ip9cQLxpns6gu2kb6swkZkWE2
SDVzFWNAV8leurVi19CT+1TP8wsFd76aZNdbJj/FwKSQHciuq2IJsjNs+JemSuIb
CqNoTOjs1wfupR1cxeC+io+b8Je+OuDpTtdI3ocKqvaciEZEkxcULN870zMJSYPv
+H8NndvecpOisAqiRcAVYC9lBeBQUhndugiFeUZRGVZXBwjsobtnSepLwpOE1ZQ4
+H591ZfORpBKgubmQEQyPSmpyDq90qO0naiuw4hB0AvXY7pmvqfuQejr4qKP2KaD
xSQJYQoIjOWhtGdy6mWUnbdA8p6RkyTY/wvX74uEiMEbtNX92bkkR6dR9hUzKjqu
YEcM5THx/v0SVlYg8eyChcZD60TkkJbZA4bWgx8x88E3VwaxgO/4rGWSSA8d+hXJ
TjYWR1WOW1kBst/vgxskG50CSGK1+kbRWQWHZzVrrXV3BSNaf406VD8HjryUaHds
8tSAdMA3eBS0uJNhmNcJ+KGziLdlNjiH44u3LWXMhKsudR1y7ndoqCpQnIylw466
p4u9nzMtLL2swk3Irj7Q2akGr5ef3aqOpElGd+/oB572s+zAcPrMakPpqWx/ewAr
FJm44f9XB0mydadxYaYmeY3pHszE6Dc1u1s8TJuvqE7b9BH7NgLteOs1CIE7oMfW
D2lhppd08SX1emQBUU6F7s5M64SdcjDPrlLRO9YRKBDTtln17l+m34MQHuG+fmOF
FrRFxkFyuM08pIFIKTUJ8JMxslU97T7EUlLyJCDKA9S9QpBh896cDsEiJ3PNHCrR
U9zQw7+Z06Qhilt6wTbks0udMiZMkaDUNupIsGs6+T876fYSDIerOnMm84ZlpkWT
Kc4tif0E4BOfYbOSeUAZzCFfvh9s/P9oWBzDIl1XVXIIsTLL1IRPBjdzb3V3p4Yy
MrEBHK+zVsBvBODW5xrDPq66vzJv0mgqMsZH+JVhcgwbIgKzWPHj4WfBNDoqWmxF
yxFRWWAO/xhcSNcRH5eGRtbFu/ISmUCm4i8Mz6Nv5P59PqD6CJUpQ9veWzc0sBKT
UcrwQrUmceK5qMJ7RLXGp0fMhjhBKgm9kCWIAEPcKOa/tHnk3/60Yr6/NjRjSZHR
1qiFH1XkM9mppWcTNuPvhmE+V5vFcP5VK8RxKdqK0ODKceWKqwqA8qDwtJItUYie
vifsBy7XqfaHj9h0v5s0FGDc6T7B9jBukiR2PkVzolCfwBr0WRe0UqUuI7CMGnJ6
XZy7mNkGajP+n6SQCpngbQBY9UbQxi0SAn3mlSTAS40WBSdnXS69bwCiStSc3cnT
`protect END_PROTECTED
