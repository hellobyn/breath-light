`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
132Dfum6UINsoMsSqf61Ic98Jujv181WnjO0sOjXhjCT8XbOYMGHkF8fVjJyVNB0
Jps0UWRkwj3TjKy6Yxk+0Ika14sXilndKSjub2WtIGPcD9hoR5sZxAVwn52fdc7T
ddCec28yOLwjOA2YKpT9j4sWvoSIvXeY9oNtOewTSAvG8XfEKAHm1K9sStY1fzXS
9kDFxAGSjrew6MZQ3P3ICAczJRENC7hf3iYxVFYjPub9PZV0Ajqe5n4YyGCugVog
yOU7bbFAvQ2fj6CL/ltrLhnTinr0uk3qmu11qnh+rBXEQZrmbIwbX1JXcAi44Kgf
y/QVzRH3baXjXyoltNh1tti4ctNeyTA+mEGGJEtz8SiIsYhKph0ZkNLE0f9V4Jf4
YG+E+Q7aBSutWVWKjbbYk7glyL5Jf/CQjVWEUVMshdDnk3vYcXVHC2sl7L6WjLRh
eAVpteyeiOk6xc4s1QZVs3/E9yZK5svSjQcXGDD1iyhSFuuf77Dt7C/JxKTxw7P7
11cePY8JRt48RfZc9iRuBa9+xKQgckxpCKLtBSgPEaMXNLfTgXIcLeckRCVvxvNb
rNX/L5wa7q7KUoINdLbyCX9qrNNA3B6w32O1LeSsWKTWbb6UMWn1jtE4XYkpvE18
e29PETjYzukMrzKm2eVHmVscOiREOW7tMvDVmHfbZLn90gbeXLi9lbJpeBhLFfk8
GpeGQDmwOzKpb44jhL/aabbaIrsy9d7zzdOVhMbl/eUe+gGoPX73BSpVtU46Dnay
diFpKskWKFo870QFOdQLWy/tvXG9JAMdtEtpfcs17hfEua2oEUpwx6nNlOwyRzoq
mNuQDr+AKUrmlZKfZD3AH25vZB29NKV1bdaw5Ub0uYxovjAiKthkJ0C6U2TReKAS
m8wfCeicCh05jpbExPGL0ooDY1LVvxABoXnMIfdgCSOAb7wHpt4oa3ZVz/1Aa5Cs
/giAZji3qJsJaf+83Irsr7POHVGR3DMCxVP5X4c6i0xf+bA2LH7eHNzyfFwyO1yG
rl6zzgqjuJZXrA5A2aMYeJ4HmMnL7HQWU9Q98MqZsFbKn5RFDvqq2oE8OxLxTXo4
aUDFHWICwP68k0HqvBW1ypzt9+3hRmwfeMNp1FGXQnh+dSS64mckeQ3BqwG2IEQj
dO3lOibcizfoNUUD7mpCFFsnsk0a12hg/Ooj9mTRn/tQ/5AAl16362X4NRqHoj8T
RoHbR9MbzATimPKxiL/I/7381a8kaGjzCK8E9zfFtDMm6FxYEMPDbaxK7sRTaVad
JJCx2iWPq8l7NjywhFeRIu1Vw7T2DZZ31O+VxG9KPVCkxJSQIsJxihrSEpZokgmH
ffZxFf5MuFWkiq3T4xdEx+gR7e7XS9g+u17nHixWh0jR87RhsuVlWaZZlhzmTxWs
0Rbx0w84gstjEAktJim/8a3pVGjYCSVluY5HEWi4P7cgOWzqfQEuLJ/n/eM+X4rD
aoKMt1Yxuymfk9D9yvsmMYj82OmDO1+bDHgmseuz0EuB6E7FPW+3WmJukQReAnlz
HBhH1+V8Xp79tHjrHIKCMF5PyUgZ8zqZMKoT3vxy5oiWuJafBiG4rJhySfG5qNC5
g+NrxGXCbJt5CKpwU2jS0PsUWZoK1jMqNmCM+ih6xPI=
`protect END_PROTECTED
