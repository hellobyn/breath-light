`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfekfKeZ6q7TdkhvSmoV3H4eNy3ewRXBTtS/UPjwU3wgDoyf5yEL6KSLCg6XLFMd
anUMLPKpXC5fzqzABAbwrU5Jqy2DvDlIw4DrOR9kpBzTJxxiSm25K+RzKEYUytRo
uOs8AqtwuP7Fu5YU2m2FhAOk6qvVcb+UOGTCvIsg46hRGn+lnpE8QvQkZlNivJn2
c2KTAUK9CaTKmy8W2qosHOVgj2hoNZV4LEus+zxhhZBXFbOCB3Cexzp84tszjvYG
tMQ+O72EYu7wID7vpWEuv12atdGI/pHw9xKOg+ZqwXhuYvVXNwMWULj6F1LIe1Jv
fDskj4sP8y9hJkcrDwuXtg9rwa+MqwRmzMoknVQ46S1RRoRmvFG9Bct2YA0+zigy
6cmBdsgVYmeGvJD78x0lbHagA4cjPSCt03yFhqJg+wAVLFzI6ynvSHMevmCjMVmL
GyRtoffJQ2lq95bHpl9yPOwmdSeuT/fmTTjNpIkpcCLHcPvPEI3/X4gomozmSRBV
QsRFqeweX+O2QuMVLVml/Jp+AGjiK2gVuTP6Qwi6DepMDio7NVI9Rt2uvhm0MEIc
B9p48MFVgbnfo67Xzc7qzxpADthdNtoJl5RGTU79y3xPgBF/HXAHsZlzXRjnkorv
Rcd0aVsgoN1Bpbi2g3Wvp42VQLzcbZTkYpBSBJ3+DMkpYNpZSbjVJkaB11LE2CCG
id6qAHc1KjHXcZIgLiKPkaiTGYLXrXxwJ0jIh77Hgw88bC2nK0fJtOid5jjUkio3
6FEccYB97tLOBET0EJeOTbr2ZIV5EqN/6zwJj9SGakdi1kUeAK2Sf/jMw96Jugj7
w55GGTc6Srng+a+2OszriXelTmhE4+mAhv27lIP9Th9cp4cPtABephFh4vHKJ3fV
PAo2sn6Z76/wnNO/OhY0mf6IJzPIvkcZ/gl552d9v+JIezcIPY5GUcFWKWIBG3Hi
pNebUrybMhwGMAJBDzBslWY5DBMGuLRcGV60pQOH09GZ178Fhq42MMJI4726lLMh
RgvcY18yZPm9KCuKw67ajp+YPrV4dk9d8cGHczzD0mEtlkMcH+K95K5M4T8asTl7
y3RsUghUWyKK/YrKJ0kwZdDJhoP1lhK6ZJZfzCViSuj3nj301cNaQi5MW6K8x5KW
PCsIkIJQWKWVj03fRQjCqQ69Dl6SuTEniR4yY5lOHca6fSliXLWzHq+ivXWgbzSM
KI4ulCeSaXb9NCEMlqd04wAGtNezhdDG3o8x6J6juX4ELDlshBzRJtHdCXxZKQ4P
6ZKVDc+aq1+fCNmEUMks5FmACfOPfaDuk4V50pSlI75MT9rw9jjT9/bVJt4QqbRB
zmdvf2D8DD9Ml16pRphU6cNjaeEvfS+/vInyEnfRV3untFtp56GhYI4ru8ETA/Qq
wssSUg0cuvrhY/48y0RO8DO1aTkF65JqV/pfI09JVjwM44DJ6hwiNkbGYLIuMZ3I
CNCZA8G5qPDeMA7CzSA2lR6D44Gjs863K11nb+fk3ZUG2SHX3dh4dRFOd4eB5Xab
ckhc4AugQz0M9VuuyFw0T2czKcCFC1a33CIXk/yEiRTNB8DRTEY410f00DlOrugi
VkJJjjunXMSjpjezKitfulA2YMG/LhUpb0EtDEBvifg=
`protect END_PROTECTED
