`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+iCqAN4iWFwa+pEJ24ATIbYNatNFWwX9EOmxaPmAuZpAh38Exos+bpf+sJWHti4
5jms8BmosE81mnmqXhclBP3RrWVcduZqpTjzSEaa7xq7cCRXexLGY7Je7tARXD+v
79hg6cWFdIGzTkZ9mvXRo4GxH2I7xGelumEtDQ+2jX92TtNj2QUNsr6g4yCnEwlQ
0d1o4gjBmm33LWL9yWlRvGCCgJuRS1OrqTF4zHDaJu1PDIjbnRlqQzA9nDU5iIJ/
ADQ0PdUWY24hltbON2CwsZS1LXHlS0iO9MeYjtyshXBcw97RJFCTNsHpLs0tg3TQ
EYmhoDlIehuQ7QHb4G8fv68E2MNpHpqexT1Dgu3hnWm4RLQUeLV3OO42gbKYeTr8
GQ0HOH4VN8X//T9ME9xe6mpZmnvyKAWL6FAMhz2H+cLIcAbp4xXemwZ7u3pR5kJd
2Ga9K75d3o/7cWjnrkGyI3M7huSClZi5GrM4LK3RWcZtqH7TDDTIMMltrf252jX1
imdP2hK07/gSXIXGQkFmE6diXOWYjVsder/l2/lNjhplDBfuSfYWzwvV/a4kjQgB
q/AD1t7ex3YckD7RYbThFK8rE7ejGPjIEri2QcHquVaDY2bpS35b+MdEEOn89JjY
jjX3AtBFiuCHFpxOuwR5bh/OA0UfxVaL6lfSJ1Iz1dI4m4VRl56BynmVgq/t6gsz
XLahfhxe1VyLcZeZRPKbLqD3hhIhfBHcbk/yWlIZUmpCX5Jr6nTzLsocHIfQvn+6
UJbbKQfrqZ+q7VGG40M9l+DJAN2oOYfzPnPpEyBk5L6zu51/hA4MifxdtCyt5kbo
75sdHkE1gSO8QQ99+hD+D6MxIL0p5PW/5kzmb1wPsBlnw1O1fUlZRnzf1DXIimCz
oR0OQZIuQYx6wXASOrO3e7UnII/1MvMZm6S2Ga1go5/R+YDjk5hLItnXYIfI342Y
t6cZk5li6PCzjdRtNHKZoa3X4ZmTYFL+oHsXurgTb5taJDwzE9HnsPGnF2l0WtIj
1vj/RvLYaMWigHB5kU3lQTh4oAZqU+yZbVOOrV2Jr7owztFWpYDaObvJ0tBAtulx
JKbuRXgb0rslyK4iHMQMrsa8mfMU55r+UhHIzs3zzcOgTmll9m6cMabAWx3fbeFG
1HfbC14FhlEJ499N+ATGbSNoIyhlJF5Vu/drpZVfzoP3EzRVmIn7e+JogiLdHl6b
LaNiSr+RWQTAsnuSwWBbRqCdgRR3l8DSp+WJZYgVmcpDkl3oJb426wdPE5xhp2ZA
Qxkj4esgK5cdPx6646qs4HHm2O9PaL+fHqBXfa2Q+hOZYxbujBRNzEp0WRGO60yz
Ju1daGDX1w4idShoEzeYPpQ8rngts/tuKwe4x+ehqXCFQEK1NsdVg7LPVQ/SxkW6
AebzwEV38tgDVqbniz3DBwNOngkKjZXeGBdYIlNj70JsWFmR+P/ytGVirfFX/2rf
KRqpmL/h9W9INwzmWinQn9Wt6N/xjyhPeXYX8/3IlxzSY/obweoztnXG9bbF8jLa
cD+fq23KvIRU5NtqwhHuCWudcLE7en6CU3vh8PbuOskotzfm6xjFToYLdfNyO/pa
kRNempwIPigGGSMD6ojcZoZfcddlamf7OgbN8qB9MadSDXFVbRG80BMQqfxfjebO
DpBuw4tblXBHjvfSbBkyVBV0jObNpcqYdtnzlGkMf1fr6qINGPI0UC8e9n9V9sm/
YlR2V5WQnjxRFLLDviCchH5bhQG5j3hygwhiqMcM20DaXhr03Dt8twr2pNbSqmRE
Jno2TbazgR3XdxjtXkjMt8HIuqgeawHRShnRId4c/NHMrdliIXJjG0vqSAWeTakT
+0HNx6bWLRIBl8+G00eOaqSzdZJfEMQp3c5YdNwkNYyX0lnryRe6Qqd7b2CG1NhN
gRJa5SQ7xJZjFK63pXS80yfkrDlbvCrUO/1nJd7wJiq0J5yvqPyEhpqZfJ5m6KYi
x+jm7e6EPvgs/vT4Zu/oJLcU3OTskyF9YD3XW80sCKHdtuNX92UWdIWlCYXSVwyY
K3wek1cK0qFpO14RaPK7LXjpORu9oJOqYG/50nV7TTvaQ8u0aWuixemgIdtVZk4t
i7NzzjR65eFUZ0J+fvyscMcyifD+cogmf6XxJfbJKNUUlJ9iCNr38/H3TNT6tXB1
WXqjIzfK44DSA4SYGW7cLaERgvRBuFd7CO0I7603HZE7DiZ3m2RE8euKlJMH/C1R
VcD8mZpqXtcdNwlIsxHywvJ3Qbgz+JbJWEdNKn9ZbN7KIwHHNvLdOGxCJxra2t1C
A/LbRB9BATsnu1/g7I3cXQ8Ch3teKyKV/nBXCNpn/xwKQNsh8v9Cp3AZsYL0TlZH
tniBR+bnJZQSMEYVE//OnySpdmzA12675DFiuFsg0QdTCYRiRxNUypqF5U+wXZaG
GV1vPdMFUNqYhEv5IpM94cjbWC7qaVSZFCWjIR3yuAyhjoETmZXKjg14hkJvQ0+u
wRMQeo7UOGv6fJmXMtiT+JRk5lKYsBIndNyEX7H/Al5NNdEMkCSSq2ITYXHX9E6k
VfMtRjWSO5Dhujl1jQhMhuLdCiNC36IZ5AAgqvZ+SuXbZvNJS6upblOY1kq9IhDP
fHFW40qLlFhliiN/y7k7CHEOJzPX0pxp1xbcVxE94SBg26y799wmcogMCuc0DZ49
6rHhkpicUSl6Nfmnq1wW0H0UcmdlGqRS9GNB0TrHb/3BYyzJcU2ryUcw6dHumQJr
SGrCRumNH9fKrnuVSQ44CkkH8oO+e+RqhBh7IS9+w28Koky9LAkF2mp2h6Rg7xVK
B+6YUHrmV7BxttNhciF+ldgb8n898QoCVRt0EIFvvaTXM1oORH+SGs3Pv24K7v/7
7zHaBG8BxGU/JIpTxSUf1A2eL9KPje+XuJpIhaiEN2huKa1cRkBY1qYBdY0M7WW/
NGltgcPrbNn6Xh3iOfgIUigdiglNPSG5Z+8Ig8S6rfrRRFKffMPI0M8Xot+ccxFL
Fqszy1KhSJwzT6/SXfF9kKfqo7IfB9OTBVKPZqxycut6oWqfzcph84gH6o21krUd
sKYhrYuRgtPhvL6//tUV8y1k/hoesbKpBhZBuN02DqZ2nj00vW7/y9OF7CeVlMaK
v+EsH1p38uv0hvN7gpT9Edhmp0Buk0YMefxbbDUZJhUBuMwC6sb4YvdeCUNxuEEK
SetWF5QngCCtWVHC9S1y4tRApdOa8U6MfPeToy05JQfPW+znyKLlNA5MhuoNQ8GR
LqInzw9v9FKsKm6ns09g2G3+GnUU2QBWiTP1lEmZPKZmJB1FMWI6imotojpHEzzW
dGgqDE9PFTtOJfG+TIgkWA==
`protect END_PROTECTED
