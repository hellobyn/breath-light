`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RLmjWA5+Zzd5dEXUHZ/b3AlC1/JJ/P9jN7hKsAvDYvi4/oAqVs2meiATtJewKM5
S2BbWKp1IeS+tiOXh3JUiKHb6se2CJhdAaRYAUH7QYkSOdAErw1P7YeY1ghGMoz+
kt20wYeQ9DbewqDZNhJCmcENRsV+8rOZBCJE1n39S0c1Z4Emx5Ew+Vc04EujCm91
XvtTsSdynoodRBAHz4+dajmByKeMLi5yCn2A1X4B77qWdH4dyjBcjqnh4RxvItw1
tbfP6gWNE0GGMxnY0z7wuZ0TOk6rq6aAlix1VdmYyFrli5C7oEMC7trhYveaSrFH
eKW5tqV0SkWWz0oJz2C7qp+yoIUhwQhb0+4mhUjnkOJw4NUZjmsWtCR8AFQf07q5
j3HEfOwuZO3aIIBfaYE3IaQrgiRR18KSZZbmAh2QsQRackJyrt8xK8+3Lf26iWj1
pkvVa45SDwO5bhtwv55sRZAJZS28wQc4Ny5GAkeQ8FudNo8J7hoTC2LQMGa2Yhes
g1g1fqeKzwgYCPturnmEbdO8rRztZwJzmlmJN8kdSVg0z09gn2D1Q/5uv0Zzuoms
Ws1rTtsdqSM7lJRZYemuBw==
`protect END_PROTECTED
