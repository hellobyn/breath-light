`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e65ZJEwKueEOWYUsYu1oO4yV+FZLQ1qZlScXSJq/r/ro7pw+X5iO2ZlpcB40aDnR
weQ2dx/fYqW4qXjK97AyjMEfmw4/ViwnIeBoPkQ8SgFWWEIEnwzhsT3WMFHIJo9V
vBPC8vOcqZ6iWBxEttKnNwsQGOHqNykXs5JiPQLm/3tnCVO/i9M8FtMFF7grFVaa
U+m2hrzVABxyghqy0IfJQZQAD/kE0VYonzUCNTdeyV5Gk1qIIGFT6xf02dPl3L5Y
3ETSDg8/XgbU/M193SKljMerdiln1Ooe09iqU+XmtUm9WTOgZ9R7ojecUkQmwsRn
jovO93sD8JBW/lGkiYWb/WiNAoOqhtR/BaPexMMYhLjdDom3GBGS2bKXQ4JBJZFJ
t083taGE8+sTAQenqJpS6QaUHaUUrddIpSun2G471Nc1ORNjqmtoJphV0fD53qhN
W+3JY/NhLO/oAsWcuun9K9ptQEqYbAYo80v905zNubEeR9rgGw1mr6eqU2KGgqDl
dIHGp7kPSwG/G/QV9HlgFnofVVrACoKp1qBBGpskzMnsG/8RliNbScnpbU6YZzv9
qPYvS7aWnNvzPxD2NA7BIXmN4jd7cyWfDIuGM+k3JUXjR+xQa+p9FS+9ZUZRxJZ3
/bBzMz+MJLLnMy0gIwcc3qPAy7LNIqweiU9KT17o+FxlV1v0jXaAiwmprRHD3ixp
s443V3Na8TbwhP4XdcfrSPTMmD+kZ7xEDfi46kU3s/htfJWybc3AOFICL28+8T9/
swpZplJGMK9Qe2YsWXv2dEXd2Gco120xBzE0QIsBrb3L4FPWmyTItHIO2iHWEMZz
ej4wBGxjl9ajym2/QKcSevc7pGmoBZAyRs1WKD05iqqlQoTOk8WQZcYWw0bF1+FC
O5EQI4/ZSXymGQDy2ZrPL90BvVpuMXVRuELo3S8OK8coekMQ5CzJQ6VsOs5G+k/8
jqUTiToPgyeHwrIZvauuSeWgjIW26iwecELhUlsn14qsbnG8zQV4s2RdAtD8YSo+
hwg8xGwtd7iJGcYq6hHuWhOngLxHAhTf8EcksBiR3SoULbv2DWi5VeZjSzaSZwVK
vYkNsP1PA/Kn9d9dJi+Kd8ThCtAORHM96dwfQL0HCrNTbO2cCZ8lFpn3svE66Ubg
1re/J+uZddV4kYG8v5SnQf6NrQr3qlVzvt42ZUQArQ07NqZYuv8vZ0sVh7aeoEgn
POGqwwHV5rUUbVBcmCKhRRV3FzWYgOFAR8oakCQ+uoQoRj3ouljBCSWRmQ2p+B/1
AXZ4RlRmUiig/7WlaWDVOXvyfgYRp27Pwk9RGsC9o6EbdvPT65zU2+NVOmUcDNp9
Y2G5TGEvgWdpjHtrn2Ns5N28UiYDS+5gUm5jDe2QjZQrmX27iQCb2YcH7ZqZ9Vqp
91DjnN3Ou5wizYzaSQ2NWl7CNWJURwzqIdO0dGq9l88LyaRghzTLzWwRzKtJGqmR
falXkO9LblMFkdtB5piElqNkSzNYW3mg2kdNAXTqYaDoXk5/yMi/8ZugwOgLPEl1
fWj+cd8tO2gQSxTjrvYnFjxv9aQ6oFS+o4zv4OVJGLsymYbRFQ8romQy74Z39NFY
2rOaIRVGDVeSibOx4/lPi/UBicV/aCvhWj2tYoLFZ1UKiJv3hUQZe1C/m7kl/Fke
7dFZ2bFe1le7s7a9SV7qbha69+DaeHzmsWRg6zK87gYjSjammqzciq0W0IKQBUvg
D94pEUmmwcXbWOSKYwI/z9X10dT63YAVEm0JixL6+zprcUNHJyPcwnsfybnj1Dwg
iy6gbWmcunuEk4zjDrJFdWDI+qkHC5CUb0p7811wD+DwBbVJqtZNdOVO53gUGjYA
SVxErZ0RKIjzEf8bkwGGxcAprHSyevk2PoykwGXfYi/F9eVi58OXsKMhvHs2ZzY+
OPP0m5gw9qHqtFlBQTCaBBeOuXT9Q9lrTJmNvD91ECV1lGQituYi/Yppm1y+9aqV
bvxTFoTOzj6LPqW3tGnjyifrrYgOmAeA2j+gO27+qXi7JbUCJHtxUVz9AuqtfI6p
Gey9K9LcTey6rLopmkccAHn7d7AzxIw5zDW+aKqBRajyL/EUDHktag9SqqhxmFaW
d8w7Ni1Z2P0O2WhkHFc5mNxR0OpZPqBOmR+zlXd1PgvoC68PrDloyK4Bh1QGYQIv
2h/CmEgU91OLjrTfnsKClDEks/nBH/Y3gwjfpEhVb1METHx+aRgxiXBUdYBO16f3
S9yJWGntVPLC1LUbNEgxfSsS5Bqs0iFF2lcsu0f/OhSp6LCANxJpRXKF2tri3Dg8
wDOgJWBA9ghqyLlWw/VVBDXjgfnG5UpyDcYeLh9Yc4unYiO5+hQNsvfig62CyiUX
DIvxHrTHU1EKC41binEk9EpQ6ltrYDe8hS7OUPmJkiNldO2EROYG3b6g6y29hIWh
LpXY2bhnhO86k+Folj6wiP48rRUe6ydLC8UsotfMdlFoz1DrnHANrb3navwFLCzV
R86x0+5iQA1yg7LERZGgabPPQVENkxvKcyk8gCoB7mCyx59V0L6gSPN6DS+P4duV
jfxk+pq6ZVq/XUjoIuwR7GBuNkCCFb4E5bsqq8SrI3g05kFOS7HJU/01CbdZkSsc
8hUmwwTLlK0TZVEVPmJQrJokroyxNZFI1aArueyTHkT0hAhhTVEXYFfHPE+C6hcR
rWX5NqILqDvZkz9gdAqhWrtBX4zhY6tHdeiw8H9DUDMp2d9ZTGg3XDxIsFvdNG/U
`protect END_PROTECTED
