`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUDlq9QfCcLPSfaW5r5yVOocRHK7eTWf0tQabSHSQ8le5UM70LTI6BojX1bB625Z
cpCgvI9SzgM0qGxV6PZ1sUrwu8pNhI2Kp5+JRtko1K+PerE3pWXN49bmdteh/iHj
Zl+8VpR5RWq4xcehVcfooFfU5cXxCJy55eUzwVvz2wC39rLqtLxETqdFCDDRdfQl
Dy5UHi9R+6l7RdYNc3v+guLwon/3xyeQhTpTwcuS2JFAwMppRGDWdsM+lvQjQ+Jo
pP6cIO8nZ707TUXLc//sPVlnF9LMkslapA7vaNojocw3qCR1+Q5MQPuRy8cdzPMD
6ZWXfafGL72e0gakwfkkrspwmnubT071gWXh5yoqlADEjELdgw7z9s567woPzuIn
b1Us8VESiChb1mKL0utX8dHuJN/DzBTyyo4pcHrEpsmWyE2zbIfvwbZFxfF1vkI4
xRI7tx3Qob176NqHVUKkgbq4lI6TEnSTAaqRRtXKaUIKjRTfJTgWbEXbL/ZiC6DY
qE4Ayf5SJG81KEPuXh7f9Md2a8wjEs/we7eCxTfx83VtDSmPtNNhgN3XRr3+KZ69
XJ65w7VPxP92AFQ3BiP/dyO7TUaVNj9mye9fFSZq2yaZHtdZkSk4mgtN0rR4fz5n
eSeEu8j/tCgoXZW/A3TgBbIZ4CIO5hOkS+w/SfSm0iB0DNMQiehj2cPKZBq9zuJj
zFZBVtMSQ31ydlOd01jYNyDi3CG9H7u2A4XL2FFjWLgsQiGtZnanT5AcE6KzqEqI
8V+tU0pnw9Tcv5GBjAz9bi1d7YmzrkP2Ih/fwLb6tRb69Y/Et8y1T1oP2KldOLsQ
GlXRVwuqyHIYeTn8q7wQKjmoyNxMGDFf2VYry40afh500x4v8ts//ugsLd6RIp82
4NdLzHOLwjPJ0KmK7gtQue41kqt/JkLcDsNSvBxQmMUMD9ECwbdFGnktjjejdZ+V
pgOc93nuhw7xJZGmbd/IO9z6m7CgneukS5IyROel8BAu5Q7GxgpyArgOho+P8rK0
0vK98wIL+UiUF1qFLcVHliEILcQzRu4TI3V4hJV7d+o3n3TmtlM0wpCJnMoOrOqK
8V8CZEi4Lit0v88W3BtBCB2M03xdpAqf8kHIg1FjxPZjUT4KLdpuOlaf3nJXw/VP
2/prXU5nZjpuSxzjdILQstWaz/kJOykwLG1H8bwZjGzTw5qohM7fPVw4CJyQU3Qi
vboaMhrg8mFYnBLeqMTkq3LqZUohMEvfMKP7Nhr0nr758yY+B+l95bQ40AUWvxey
eyi+R9baG7phTovR9uoGNcR4F1bi5XBPaMypr3f8W6so3su07xNYOocI0som9hIw
9IyoLp5IzaoNpVLpmoa0TG+sDDpV5G3Y7npRjDneyRtq62k/FIQh188r8ZgP+f/j
NbYDEvWfVFoRPVHwoQFZzVNBIeVyUkaWdo+oYzDZjBmM+mJ+UJxqpb73V30m+EY5
`protect END_PROTECTED
