`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YC6xWUIUGPlhYrrKn3kkQtXJrQhhro5R6A63qARzZ+Qfag6NS3R5jUvwxPhXmg/b
kuSt8Ar2krxf2gNWFLbnEabD+IUedzAWVzyNTd3cts7wW9M6MAxb9RbjIdIiiwXg
GwqkbWGEanid4NB6EZfys3YQ1xBz84ooWqTHsyISlMyAvtiv6DSjRs8FLlpFrfnd
BV89+Rr3cwVfrrU++d9H58CODnZBnF40oBzEFc+zqbYQMLH5O+KtrMESSYoEskrP
1qCRvAbvfwYZsVmzKbGmA9MbwYFzPzr7tekxHuJ2AgOizkVxRyz7dLWqVlyZ/aV9
pjopAhD68DLI5lCvRo85aTgkJjLzCBrO5NTA2xVgCE57+/aAftrKcLyHuOxfQvYc
hEjOQYzlo1r1npg12CE6UmeiNFlLQ7bpiBLuXaNeKVOXCBTKKgh6HdVLwnY3pfmz
iZj5tSoEV6OdVcBYSus+rQ4Scv9BXWbddt+1uAVl4lz5t+Z9XiSNsUEmJa5EjRon
vyZThY47+P62NURwmKui4PT3SnY5PG8ovD4JdqvCxJ25iIMbZvifmrWK3DTscKxD
SJ37jSTS0DDdO8sLpHAULjyY/SgZT9RzqaWs018kokusFMcqaCsaWFGkDHSc5tDm
1AoF7Vz4KB+jE58O/MH7Y8uvFBrNU65YolBsFcih1YMTRrOCMkvcYmP4pGPXMCAt
E8RcgDlq3a0Mk1bFXnNuh0I2HeC6rVCmtKUmIMzM0ULQS7fZSpo52TTv1eVEgPyY
04ZwO+TOL0dhySEkjhHxEnsMenPfiwIDJlSrlzN93E+kpMp527T5fmO410b2g0/z
vHBwCw+9ECRY+FDospxl3CMjcuW6jzk/as3GHuPvfj6lwGe1ed/IRj/qHtA68JH8
fFqAYlQ7jAnGxpBAidkMJixWvKNpysMM2oW6yy9rmfOz2ZrqhMtXhMq3vvRececF
IwwmbdL2Axd1J43tyo+uTCyKBoEmC6VyT1jyUCdinMiNTdUGaDVfsUJHrCsSj9Wt
a9IxScArGh+NWgFdiZQXrVa8q3gcZHOvcILx4YtKPHJEyQOQHh+7ZQNETiHNjhUh
gXe1Mc9PVyAL7cFiUu3qjH1uD6914XeNqUU6sGfMnR5SlyLSIXYMdl4wLiOB6Q2Q
/fHftGISP3k9DQPKSDiLE3KDCXy9lYmklXF3T5aVcrnQXMGe+Ui7fn1nh6xjytU7
78mbfkEUPAMRrQINx7xLHRx2spvU0gcdRc0tYH9+fixrxH7aDpgoDDtxRE8c9n93
oMd6JZe+QANkFcfQ1JD1lnLNod831y14X3n/1T1EmHiXldHcdy5/w+szzJ7PxjEC
XOmchzo3NlNkLUV8mcjVof8yWY7JhttCf9GP6qCMJV+KSAKFCR0Y9pukH4MFMVKx
HFPYfNrTvBeIcE4NkItP26jSfbfYPqFgXqwon2jfOyY=
`protect END_PROTECTED
