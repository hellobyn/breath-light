`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cosWnMcwwfOlZPI5kGWTffn6e0rm/+7UtLmQa4L2mc12+N8sLjtAoa9KPKVt+aNt
tSIfn1Uj+/cfYcP0qiH19NurIftxGAJtbM1loK/JadW08ZRr74cH5Jx9P0sV2606
p1102yxJgQrA6gJ6Jz5EyWMixFVJqzgGzLbNM4yEK6bnLdc0ZA5OOsyvxyf0yIvJ
KkuvUufncfJK124DJbC91zpQgyEU8htukvkfear0eBBgHR0XnRQf2aoecWMwgfKu
anT4YqxiA2K4eCxJVduuZHWgkhthz7ZdS6AIMiDdhenEyQgNSo9UELVfPXOf2FkX
F5x0mfJ++dvWXPeuV7PJRWxA3lL/AadCTp3CbZLLswmdZI3prD+gdTbKVUkw3qUy
jrieKsE7Fcnib+5hMhmrS5Rp8b8T+Jzyu7TS0fvOnDSBw9EKE26T6MlEBYZOxtz7
y6ykt3I9lUdmHAU+aUZ4xXeRm75d3FME+SiFN5OOH5OBBVzOPzCC+qfQouUIcyQr
fA2NKw/p3GA5xC5r44MlEALnje0kfn4H7blBZrLa7u/rp1g/YtqSAYpO4DQKDpI2
xHYRQk8C9dAwhvKCDMripGS61fdRQUYHHkKmKmeqd6deACZDR19YgkEpxJBsfOV/
O+DVXsiG6jBkd+yvhOPtFaMsCld6LbCvDA/ugVmUVPqIqjBh81sXjzU3xoB1+RL6
GhErnDb2GgGUEwXrqnR+EYOvpyAKhEqOiS5VImeNeXxUYGsDvnWj6CyRhjOkkbFN
jNcQhZclq2gvJeTTQSp4zV0Aw1/FpkhoUPoGOVppSFE=
`protect END_PROTECTED
