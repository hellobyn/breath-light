`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDPT+lSSm0OX1Ndn3yjk++mblFnmkHbSY9lgWTmqw4K7vGSozSrGvis8m8APrmPX
z+IqKY5EzJKOXL46SFmUgWqgZbvaQGUaIAHh+CDwfeMxbF/+F2d2cjXRSFz+fjOm
GdLoWLN3KxDLYJOOyDQR+xaBiIBOzZlrNPJbfO2Pc9d0mMsHGkAkSUdNMwWOdu+e
hweJwDiYmRcdcEh/gJkZh5VQm/2DzrVzm/cFRes6BZbPzdHnZBcVmRgyIpfd8xUA
mMXCdy4wuBiAxHB3pSNH6lDnrya17EiyGOHAUSrxu2SoidY2gNv0EhQxehA1i6lQ
CcAK+dArZSQO8PbgTELVtpQTIC0wylDja3GDiEClsJRLq7ysN/yjez4BmXSCgiFy
HCdqZS1h4jMEMN9c/jyLbO3HSugFkf31e+fklIOQgJ8p0cZaX01NxDOPnvDW86e5
Dt5k+aivxwfRsH+nhdbRfOKuX+ujumdQvwppMCV+ptPklqsXFg5TfAJIGgfk5rTd
4Pqe80DticL1PTwtaE6wFFFC39+EE5G+3a6mybu2uYtSo2TR5xoUocUknMUjiNxE
s9c6ts0aXBmDXidSgiB25wVgN+tEo8e4jEa/pWAGYg5ISCOuIXrvhXR/O5zIaUH4
uePnQrWpm2+Qdm4stfinNR4UM0gPTkKTR+KHYxUoVTbBFQ3eek/ITBJHP2ox3DKd
fJ8i8uX209zejLpPJgZWs6h9Pe9t6D01A1ehg6J2sIbxFd5eEmoUdUJ5bdC7gnAj
POeBkVqr++tvvH213GhfFwkbm1F5EcMtkUjLRBJPI7AadeAtM5t4eiP8eKjktu1K
L6zJq8YibRFp5yaFhQiEb+SfHcMNPYbTxcCjJqpS8Ada5I3JDhfzhXD1KdgKWIKS
PsegCvhYFeyZB8526nG73OHv75AodRD7c0Y57DzGwsQ1tfN0THHPdFAGkrwxdA3p
eQxL7C3F24X+WjU4wiilwqp2yh3gZ2p2pfqW4OsNotvn10cy6Ar3Ie0KuuVEORiQ
xc6kZrKzaiCOwB1KjfjDxL364m22Q2B9t9y6KR4qVhCp1nc+L5r/EM9jecUTuHAd
FQTUuV05xF/iVx54+cns/pXkDO3GWRfSHa+Kdl+/oZQVMRFdTLo6AB2dY3ob44iT
I+ANjDGGeNwvKDNFBpZiyi+pJk9eOPiaOGxp4TamBkoaqCm3t5zg1KO4AHLUP6Ha
M4GbjRn8okK6rU6W3BRcCsLHv3PTS/Pjv5P76P5F2WjBLyw5E71rbqaMbBZNw1X8
U1YLGslRJqYLZTIwV1UQ45DD14S4eqGBp2Li8j63LXVx6tNpuyYnnKqPd58t2yyT
cXNbJlcR7EcsJ9Ea/yfgat6FFsf/hFqTQDB1RSp07DH+gPUbLRje4G13cfpskzFO
QXQvQqB4cz7TXouQcxenzcLMsc6FsIytfyyBj1Oat8BoJEnLlO8rdKBYKe5T7WsX
YHT2ffGVXYNF6onr2CtgPKl2Tkp4lWuFE17pEv75LIsgwGu9qWbgw5aMa+jhzOte
ZAAG3dxVSMScWVidzFWEi/z4Mzb/iYRATN1LwpDiAO5N253Pn9rxBX9vnfbxE2ro
j3yYoTQTZto0xJfvXic98W+Dp1sYXx+RhJjU6UmwyM4lD3fCKKIUc28Y1aeQBseu
arDyllXXa5sgX+ocMjw3TT8QViYmdyZWwQzGwtIfCAIl6E9dM8GylPC14/2I2L1u
U5gRAzy/xujA0b3Z9VJTmQ348q3fArRo6kgADm8Nq4p4Uk4nMI6oJgod5o/K/Eqq
0ZQMb6vGt6CH55qEkBzeYBhAvQwS5FW5ynAyClfTDze4GO3Gxum0/o42wuVM4g77
L1VLLTvcAHX1Gp4kmjreSX69la7+VYl7geHzdQH35TQJyiPP//bZvYNHkanojG21
J5KIeivntcSpvYVAWv7PMsdIKpqrSxcU2Hr9XtZpXC1GdQsPblvL+wlAlAVjIWap
tUBNYOYM6jug2DRxc1Sc0K7FbPmBbE9MzFU620FvFj9phaHCveFn3m5fTe+DIWY0
XwaeKsTx/cGTWi++eU8WyZLdLPjQPNjnRJeDABAqPg6sluQRBOpwtzNL0yaZYDAx
NSdCy7F9p34DVUOUnEWJpDgNHlIEXA1YKknjZGVjcdUIKQNmryOrlAi/KPI/agzP
++yC+XyoSDMX1drgxPIbgcU8XASX7yRO5JArjlK3eG/BkW/Kfvoe7yb8fs6O7u6b
bl3Yu7y7L0ERVuGsqIqp1blnoKVdbbm+ftJ1xBYWlpy+WC9OynffLOqQ/7FqwCR/
jvgJhniDdKiDGnOnY1A6i9k1I2HyfRwQTs/YQvp83FI7laUbeoOYnSGGB64PGZ5D
1zgww5KLfdKlXT5wj4gsq9mhWZ9MwJ9lnedh20lkG1MKDU3wvXMpflUeM5e/XNOW
aebfEte2/DEU7Qp57/L9KcE12Uj29LG8Z4Q8JsH2tsGiPc46fCfuJlPF2KKERPL0
rn+fFYSvkvoZWHaXW10swMSRnBk+LvKZQLtcH0zJDL7/WL/zMc4dO8atF6cYC3TN
o/RXuT7Jn+eAO27hLllvhXJig1p6Ni/cHwMJfWPPxzzOem7KeNWJdSiLTLHcW6Nz
pGKnWHZDlFngqLjDEFzsdzXuJW9BRGssSV5hrIkMs+RbAsnpIkat7fm5+YbMLZxV
3o2N5CHxo7KqJXSmpF4gIlfBJo345PL0DMZRdkU6cxcKUsO3eIBoQNnIzxT/7Crh
2BJY1P2RAHDZgH7I8XzgQ67I2cXp+aSxz3IeSPaPeeNeWIIr7zg8EbL656VkkjGG
r5SXVCUx+fLk99j2v7yj7u545+WhO9vL1kBHFkvZ0SvzSxtKPdnegEzgRxP0ps/a
3nN/MLWDi9OiS1ILSmOX9RWfB3MYaEAgql++AtQEiY5yrIIcwsTOBDLaVqQ48doH
ygUue9nfchqU6yfjd2oCwGyhStnZQoneltLp8UdjEVbQrs4Q8KDp1tu4JYJs9fdS
i63enjTv7DzR8AshXfdnS3J/FYCQZacJ8EWhDk6CYYPkL+QSCEl2MoVnXGRfc9cR
pHHwZlVc4WlOvT0G5inFjEosx7GxNmcT/2qjgs1F/ys+SnlkjeVINdZWOxkTwtkW
V8ehwOuxr6zyGIt16Ne+8981A9ssLxjqKXmzrUg93jdIZM5oUdmFXXBFJ/9n2/5w
tdRSitmK66xU4Y1kAZlbxQ/jMrGmyoqOqY0TgqQ3HKA9Asr9x/Nx6chaBd5Wv3lU
24icILGT2e2O5v8xvRZBrhZTGrhERwqkIM0gGcCOXZoV3lTnv+PpKcCyFH3N5bfL
d1YI1fxWu7GOdxCHIfVtWkjvhnH6bSQp2fvkKKwrj3st5POs5NVN/OiLYmpWc1BB
JyHgwy40TK0NLF/B7yzFrOqfGZxAXzmojbH2MYf4OEPgNVGpPZrHfKbgR2bGv2ma
GIpkYaGEML1Qo66NlU5wZFzZ7V8bm0QN5ePK7T8ykuTKwXeoImrmp6nADLJVxYu1
CrgePKIAGkTIpGip8Fn6yCYNwItdKhKrHnoOLTG36hSBDV8QqWdXzQImIM4Qesmc
5Vif4EGFOunBZVepkCJrGwcZVFY8Tlhp0wQrHaFD8B24pS6CAwE4PCHfW/dvvEAl
qmm3XquzqO572Pas44ooDyr5+Mxe349emcPMsdFd2R0JK0z8x6y83GaD8hOAFRuS
g07lHm5HZMIR6c33OZjXFskWgK4JawvCdhtWSlkyUfRakm1olrNvyx1Fc59oGctN
3cZ7RVScjTue2gHasI9vmn9wF5wUDjSc4a26f1d0HZN5qEiQj31HhVK/nPxISR93
ay+8fdv6bnQ2b3QgVJud5CQKAogszkTjYPIgFNgOTFJpsPK+j5Gp4fTNknX0faYW
7kUSvZE2QxFwlTTV77OCqo9eDi77qo5J2c4OR6KkBy3L07qnUf4G+bTAHxPa2vf3
qT0F9WqWec8MdNNMyfKEDgHueewFQWgJXMCac9VLaZFy4ZmVL2zlFZAVssGtfLGo
VwUhZNf/t42JRuBffVivZ5gebxmI8MKUjJBYdIKQpD5TW7nXHuJZkky8G0OFaoTZ
PDtevjuXjrfkOKIPiE+s54K6IKjm4ekROWNi2NTjDKsEOkQateJ8gxmNr0/xfkBV
NBga4nla95duEQGwn45oKdw3Pu+eRgXIL5hjgtDipFPW7eqpvrak+0Howt1PbxuR
urJRTcViGkTdYvHXJk6lQzPks8sFayURQCeDMAf1pbG5LMKMqSdpJvX1YzfwHh/P
xbz85c74yCQtucD2CoD3rWMAHvLF4P6tnuJjOh8VzkaWrE0WqdkG0lanAB9X/bsj
oVn98U2obY19mltfPMCMAQup+Uphmfe7A/XBQfbFMWlIvOpNLJ87U76k5rgnVNqT
KCPPGd3doVH5/8NzXSB91Ac5dXwdqmC30sCWw1T6pCGmct6TBmOmVsZhX2r9QMyF
VQaWxIcWWD51SpKmk6gz1bzaJGCnDsy4iiIDrZxIgLV3glVL2USbOHtDw+r9mgVW
QlqrcXL00dp0UzozHr986EUPRoZLuUFktJ0DpmohROqbFLDT2eM6dWaVPYGko6Oy
D9zg6E9HKaltpcCAgQ2uqnwfdBTrmTyN4L9QSaTJkLrhCyiPpzqeQBlGzwyPClUD
O2JTcxXzkiQDZRmA6hq3afZNlDbDt0D9TjasBxuzuefpjzIcNBvvoFktcqmlhRdK
lSRVvWoTDFXS60JN0wDIOGMCbJwiVW08pav8OhKZsYO90dNdIc7Mmo9Zzuo1D9IK
8ftjCnWCOorg9N0HzYdtN8a5poKSMDM6XFj2qSRqCyAvdf+MKQrLu0IBU+8PmFEY
rlafpjUJAv/qU7AaXJdPDgabZweVnlx0eqSs7qdp5/3BkqAcDWEB+u4Xt/OuOlOh
MF26w1UwpEoNVDiv/3khAtH5PH45+FID4wwyl9adZ6uQcpdS1NCz2U4u58vxxLxQ
Ivg+dU5sXMaKv+chIS4d5FYdM5WswEnsyMLNrEDForWWkZUqJwDE9MSGe2zTAfUf
2xOhTCBHstd2Syacj4JXneKvxPjNSV/wctSh7S1g2UfjSWvntPXWjYwqloMIbUgj
t+S1ZPMt5BjA0xkMZrE8LvI/Zwu49TzhHw0aON0P8cibu97C1DYuTV+yR6HTGDzj
JwKiFzRuz114zL5go0wVyQkxeRm6jZFl9GqGQopWPN16fWI4ojU+mzW6jlxeWi+g
qPEckR0jpDyN5zM1u4y+o4qzHXhnVMEkqZdfZVuSOyb4Q/IuO9Tx8p/g7Q6KqE2o
aCLXz8UN/vUhsVP/+0Hu2f2zFNvk6QCS/jTurE6mY02y/oFe5njFTb1hyDTFb+sR
s7gNv7pWqeE7WmEpZAaW127LpjxtLEuG/t9dj+oqByMsye5m44jn5I/BWowZ86la
X7onsvzfCvOf1S0MT+IHzvyK5piQwc+Bh0Z76ueYH9K9VZBmI80DTUEgENN/VZns
fSSrgC2qk93LbCQijUF/Mu7RM5vog/IzDZwOn8TyDBvbJJitWAIVBSLdfdJKcmon
Ftm7L/rXh+TsIgZu4qyKA1G8UpC6cIujeD1MD9/oLZy5uz8sG2kMAl8/Ftw0mtQ0
43QaxvbDGTJIIALq4dH3je/GC2ytDIfnmVAVoIOY5lsRfwyeSx9Q4rM+JB3rQpiv
QuG+xQOtfwi2TVVeDsLoCIkM9GHKsAK19ZARd1omps8V0MzuIjuWZfP7yARS1Sjr
iUqFyZvxO4gssSuFQ4Mje36yHyuRMIgm9VX20VRckaWbrnTdy0fmU3G19uOFnL4l
lRSLPJ4coWegNUhth14vR6q7FvTBkOo+jQGEKtPo+McMerIrCgvRssjh6y2DtJtW
l34ciVY2ic3llD0h2Jwu41ZXE3FVVCQW68JXtlCCFY32GfZAjBm4koOMgFozPFLN
dMJddC5xmD0ZrkTpi1XKMW2HPT5Oqsj+OMYUfV0jTOmNzDP03eca1U90B/yrGGOf
UT/m5be9+OV663lMWZO5Jbboi3mx7ZYUBq6ksHLaUlch0vDzu5RbZ0/VkIRlXRta
0vfuiMD4v20OAMd1zvEOWunZTFAgSmhRX6dkJ4ydg5jjRN4/1IUyWlp1PQpoWAjf
lQr1Qm5dNS0cN4KGuqLFVT9HukmE5+S+sUADCcvp3wueVY28Bwiw8mpY/j5lU2oB
UVXxRwS53JQCjSscmSk50Hia52AxfkwFJ7XwmRuXcGsK1DnWwWVF/66dnsStr2p+
7kwi/fwbXN2SruDja/E/ovZ0LEYEWOJhDXqrawIHD2c8J8yH31EGwy4XOt8iel4b
6JSNZGLXVQ/WvG6gy8yghMmwT9nhdnO57ZalDC8/g+4+fTMS/WjgjQxJld9QMUBk
jh8oPkhr01DyHi7MUm59zpjymWjlEw9SKgj/NiQHtvI4SpuBEAdM2AjXy3y1S2B/
7emZHVGNHOqBdrLAz+9UzBSWh7x7cXgMPabk6JXXJNNWsXDAlFBOl/eFyWyTgqF2
iB2nFbxWQU3SHHCaK9NlrzxivbGuDGHweecRR4rUlPzZChuaTLiicsNVtpi7kqnP
L40BOFp5hxrLqcHvx56JkIuqA7KLyKv16wJmzrDMjcTRR9jXimCxrnNCmQ40kL3P
rMF69/JqWIGfIZWbq5IsygYaL4xsJvYbS8iGdCv72C/XKgUIB/QzwYe93VtpcrBv
f5KsQ0MkpvjXuVSvK4umZklII8QPs7fzzrpGvncO5gwwfrvYs6gCgt3izeMe3HNW
+V1zV/qQDib/aPtUpew55mDpJnm/5aHi0UVJ5M28yaPB3bdBWg5rFPCZU+HtylLL
eJ5Nsw/oi3wnYz+7qs6EW+ORUhp9YpjHWAPMZtQpdWiKXyc2J0vDWgXGxVb3KvR6
LnTGraWSyqt0KLI1l8wKwKQfUl+zpyJ86EEbtuzPjlof0Z+T0XHudTFbnwhixqyG
Rpj20pWiK/KLUCfZ9SzwpdLY1pu5lr9tRyXze8b7P6ZGvx7SKCOJDYh8cIfvnrfD
ywf9bnhGY5F4Z+jveaAuZZX+UdA7ce2ghwo5+2YtAF6cVAmy7D77pKUJ6WKbAULV
CH8Gqrmp397KR0kR4NYDFpLLC3wbbz7p1eniDWQtt0sQABfRxhOB32WBZ6DO3CVU
46VkPl4yo5miGe/O3H5cSPTwOcG21vAgk5ctHWvf+fEldOAYYhhkroTQUmkPuUSx
VQ0JEZD88x8z3nTI+bzjcqt1T8j5VaExLYuTQ+Ubawfbyu7ffrHfxuZJ/s9US+nT
rdm8QYtgpRIVf6DQg2/UmKDexNmSarW+BKXfhl450Xj1Xu1MjK8077ThRu8jWYfC
gfalzSECMtdisJFedzO9m3rKw6RjtJmFgGqx0UyUf5NSPWi+tRXVZSS9X0MUFwGH
m0lUdg8gEvH/f4SOR8pVBxHITqcmh1CDIj7xcc+sg6YfksTKj0Q69s4GSaZXEtPD
vZLUgI2dSbRn/JD4ALV0EiwD2d9gdWUeIvF4anT53ulln6kkvbLDUZZQcV0a8Rg2
4J5FzL0/e0jRq4qEpA80NTIxS+YkrAIObt5T3alyLd8uA8WetSH0xXg0HSuSTbVp
Yow/0oLC4V3VJ5WcsOpAj0o7bOcme7+MLiObq6uoUomUR55XMZQE5CxjN9UkAVTG
7SsW6lsUZU4yo5bqk8RaZXSlSzlfYbQTRtkiPkm0vCe/O13wsFyD4SshVA8ztj/g
1PPWhNVpP7fMqy8Y+luLrevcmxls80zOhYVz4VFsgL5ve7koMX5KR3tgsUVaBDIv
IXLxnPUW96nqD+JB57txbGG834PAhzCmmiE3v3Agmk3mDJkf9UsgmJXl0LJdXyao
8ViPM+iphdgz5E+1bbNav69OgzAs7UbjU7+mQRVlyZWWD39ujUDp+4T+JLrTQJ0+
VMNnZU7tLdEJD5e6cVW56dZwyDmBsFV2puA1Mi8npszXjBMi/WC/UORGF7iMyzFV
YOAb1N69FHXt3+vt8OFOPvj5pKc5KOIgk4Sh5iSfGA0MmCZ3LIvjJBeGgbFem+PS
s1Jfi51qAMI+QSHvym9Il6Vj9VUGgF4AfoM4UcjkhcOoNM9TxHdno3SLbUpxWznN
9M/ySEVvTXP2hlRIhU+SLxSyuZ40sFkigh8Yu8Ux83qqifyVsvN7PwwDMIpYUbhl
JbPEU60MQ5RjuJjlchaYhDagkNoysXxggSCWuVJ7prDJhLeOsLAkMFnG7AWhPX4Z
juxOa10WAlHzW12TvXaOtC/w/wQCC+9OGQ2QINhZW1lX1cKjJ/nC1D6gKASw8a2n
d1k5BMHvqiNNz9rqxqs5/glWuhxlnfHD4wWsT9KyhvA2wQyBdTxU2869asZQ/ky6
kHAGDK6yubZGN+xfEufvt/f/+0B3VL+LnqH6DQ57WVEg8lyQ9nc7hDkuaXxfPxJc
KM22O6AdUDxH1HmRkSiXktzPCMjUpoeJbrr2DlOLZGgKNRU9fyh4/g79cBZ26ms2
M2ITPV7zgOPQXsfcStmF2UloLf3pH04esHFoGlwScAvUHFRohq93hXnU2wpwaTu8
H8ZZjrXOZMW/7h0Odi+j3uBVkVJDDXs1wSckdLBwGgHARJjx8vYr6pw+D2ySvVag
qDHLC37+SELxjC6qhOmhnxZe0+flIAy5oz6J6qyUTtGrnKN9vImnvSq26MrFfCHc
gpSFpnrEls5kAjc2ZENKV2/LG4/vII/NtdAGWnTOboPRs9+gXDJP/hO79nId4M5H
jYO+jqr2p6mxV61XwfjUiVj4LT+GlpegPaj5B229ZDje9nregyLHP0swQbY/5Tv2
Ol3TOnd5RRnewxJQQH9F6tSIx+azY1niTLi9DzNuK+ueaXASlwnUYXel/zXFNgwC
1JxFkj+4Odl6hNVmZU3dxS74CI6ec5dF6i+LhQpHNgIQxgtJS60dB6pkdzJcwnH7
WJEcgSM59mJ2Pl5omXs+r73Uh+25SMeO3QiShuwfROjtK3I4yBXHcmZdRYyBi3TK
ay5BFI6j8gPXY6CSathpxDXR3R8Tflhcgrg457Je3Ay72JLAtYJSsS6EJ/Wpft9L
fv4WLQnjG8j84DN+GjGCISmkChmIYpLhWB6Hp8I/MhI3EbDkQE2LLaDfVPOO4qhF
szIy9TgmYGFU30y9Kb0agUY4zADRhOC1oWAf6rhsvbpzqSglqWUKl+qLK3TqdOoi
a7fTW/Us5CNDa5iP1QLnE1IKpaLH1EmrkfILuxiMHgoOFAUo+lw/TFx8HRY499IL
1Iii+WsBzWRA4Ya2fcQxi3t93JU0faEhF+Pmw97S/efbC10lEVepXNocAJWbNqFo
PGprpBeI7J2tjQSfG6TSatEDFhKzQwGDbA6Gu+Z21YyuYyaM4unxpUtzDXvXLI6m
o3ompljyaJ5+iPlKoY35YoCrj7XTG4FMAlHeyv/C7uBtAYxaXmw8bdoWn0g6UHKE
pXPX+5+Cr16TawdRP+N7Y1D4tszldczTmCKbmSk1gi6X8DXTO193s6ccoznCq+kr
8l0nZrxzfz8xoNVyBavB+B0Lb6h2jao7Pu6ct7+YezwyeUqiTQIFXGON5vkBWsP6
TJyLIuTRBLcpHWFD7ruXep4aDQ7OSstF8ik7+NX1+tyCgPFci8RMWurJnl+jHzr8
SNZVqyBDhKrO4MdrtRA61gkIeJUbWZTtqJGoA2ZVghmBdqNk82CxhRxircl5lIZk
0rG1kJ4CalyS5N1+CLi7oM5lA6VYq1OCm5Q13MfJG8a7KFEX0P6aMCexvb7jPt7m
1/yPdKVqI/DVRwpcNBh2OZZ4Bs+ikTCG0Kx/gq3nucY+kpXtShP8lANKn8OJgytk
wXG0aqE0I9RxcjV/h/ZTNrrpLR2Vr1j2HlZ4EcdYmXBG2GPXR7IEOKOuFoLiYhSB
f/FtYZH+8J62Hivq+0nDpVkyU1/SaPQs7ocMFtiB0oJptORnk6XP9Q6XDfAcg/xB
zKte1j5Tb89ldLpGtborqBrFk40+2DlDS+y2WaEQZfqFUIG/bwA9a5xtWB8NDbVY
7sJjgVvTShEjGxRHAbtgmgJrjJD/ZPwyPFSIOWuJGUZZq2T7R6WBiuH08F+pzj0K
ZIKpbSBvJcXYVWP6JHEJc9sVq7th4y5LbrPTCu7/vqenZ2oXYZeKtshpP83jiIRq
eX+A95hzQoZuMjlCN2gxJEVcI1Q9ilfQIdzmKjwHsBBy+PfmsVnrsaH1RT7kJ8Gy
+nC7slbU1s742Hs/5zHDAcHDw3lEh+tiMLiu7oEipvxK8nc9nbL07ZVkfe9ZhWmQ
lsvo8L7+0DJxOGvISccVd1azemFFZhhwCoai/yEY0dquU4cLwAGZrxEF6O+tqbsx
BnLomvVyO3bt1NInDdHpUS8dbnkhS9D0xFaeATLPrWgGfEvn+LUTxJCgrNbl0naL
I4XSCDc5QZJT9s2TDRvE4zyzEsoewHw9Anh7gR9XJZbSkgx5bhHGVJtdzKRCzuVw
fgcevO5560ZlZJG2zhKsideP0dxqzI2gOwcZa5FirrKOhcIlQqaCONB0wmm0K9tu
ShUBBQNad4QrQ/dGCtlE9ILgqCU5Nx/83oJcvts+jHd2Z1/uWghPEpS/CVHYpg24
oZekjjZZDeYkU4IRDNRsJVqjfKqJQXDvK3Qbpxixe4fafh6hSt8/RdyC3Gf/AvW5
Ho7fv/lbH0YXEs+2FZAka70d6RZbbiUOaxncfoTj7fER3IwDdhWM2OLB7Zp1ssxU
M8lZuDmhvEkl7xqP5Y8Tcfyu3iztWMfasrA81WLWEQTz66Kq7Z53yDgr6Y9xT/bm
o49c+ZhYzce6dFCrbAmj8d/F7HpLK2ISO0xCsob/9dfzHPJuPR9kin+NShR4lvCs
2pvB9+EsbfgrXszwubU9XGh/WMZRoO0gjEtgUimfGHol6sWF2SXBxX9NWax5xb0I
KRpDVl5c2ymsnjgND+BMAGcIbnBIT5/tIVsUd+RXTuMnTNqYuLdoAgKfl+7jU/XI
CdSR3bLN0ptAYeGXxXT4jCY9X6oVM0Pob9MAb9zfF0VBcfW0EJd5lauF5JqcuIjk
0iuaTkRKfygq9gdUZZ6kFFGs9ZwhFEluaf7z1YehpwYw/ByAsEcyc5o7BkDAJrha
+b7HQL0h+g59i10noVJo5gXYfXpa0owE7Vur9Smd4W0/nzJkqmPwSBN2+zPTqM66
dCnPKg8b6gss2VWyDMBYnk8JqcBNUDoGj27PCqwz+yELgIhuwYy50iYgml2WLQxm
2bz3N6zmJ6lyuh8UqfGRlUXIjyH4N93lxtxcXoKoOvI61x34vGeFkYSSskIkWTVn
/H4Joh3EPC3rhtC1UGJAjiZ61JBpo88twsRX4oy7SBrWZHQyHQ9XKx7gEvs6KFOx
7xJlyafjBMx9nNaKc9GPpD5iq6su3FZE+zXAXjea0q1XThQB3XQH5dXIdkKGIcHw
YQBUOFxqwNjreCUhk7yIrAgNeozNS1CCbXO4PGfx4DYu8uBroXnaeKJPZSt16BxN
X6mHcUzJWUJfA64SV4BdAWKwayRYGC44Q2xdxPmd8yWAp+O17ZkP1oG8sZvKtNpa
uu6RTEcZ0uHGq25ed8FG8qOxogRnwTkf+ldUWx3PdWZFsSlkH+roPyjslpZyX/ut
jf9G3DzSOTX6hdzGB7nqxQf+tkivz2VmgD5pD1Ddjj7qIunMpkSro9RhF1tJ9MRk
OfgVwteuuGQC50cAeTI4vFDsCxdcHVm/iRBCt1QaH7yLovMqlD0jQpA5dbdiIhDG
LVHp4wQEI8SvjsbpAS29SPEGEN9eymjXrhgjmk9NQVHap1BzyBumrSGwuWFl8ZhN
+HYTEuFPIIm0csnpf7MMbQ6pqxGqL4bH/pDRy57WlDTKyqdN4672mHnQEuvSRlEa
KEKwojvoAdY7+JZrmxHmenyG2wScsd3MXNT76bY78r5Vg617xlE7/9T2hNCfV6rs
e3NBkLaXlDESf5lzeMW+Dsy6OuY7e1R4aQl+FMToSa6wm1NNDRcuLmrnqimtwGFs
gveDXR6AuLNuYvI+7pQNPWVlD5E3tdDsZrQj1vrmKoDFWslLcVB/LcQ0SwRGHnBK
vHcKQ3bsRMXMh8pv4DdkscnOLJEKfE1J3gIvfqvWstnerCzoQgE2HQbs0taaMWOk
n7CJNfqOAt8cH6W6pZgx+fhPhccOONTJBFVuR30HK6Q8trXF2BfQ5Wy3v3WTB4qR
1xWm53IaU8iid3C0VHusnmYSJ6ahxBfnxUYtP/l872vIHkW3eILCsyIQ0pnA9QDx
jGCbpuX7vAau58mXq58BS/q/T/k9O7dQ+EA4b+RQ0e9HfjnrbL4I8IV7VEgaZzAT
864jZ0xagUFw/UQlml97jnzrmDpue+ROanww48GeaSOL7gbCN+rYwxLh1L3j2LCN
CpPDmzTDXC3GiclOI82XcYC7h3w3vYfGQY005UpSyvdH5spJY55mGEoClhdcwc95
sEYfx71ZgqNn5xEmHsaWvEl2rTsfGqrlE85zLa9FpQozANVTrye9kSdiKmd3CyZQ
kNdin7EBMVnF+eoOKueL4mjeCXpzvgWVFsN4L2hOrYvdToa9X40Qry1xOSafYTXg
v9MQpCtpulrYSLQxEFAQJWkUFLIFwh6a2q7YqUqvwAIOA6NqPz7K1P5vhdXW7BXp
R6V7cwTqH7xAIpx64nIi3Ihz9veiXmm5DXH8Wv4xt1DseI1psuO/NDMB2mcAvW31
qQ4UyRITdPvb463FyXwShxnJFyELJE4U7ppluyJ/kgRXb+N3PI57eyYpZzwhtBJi
HyfQJMqjqJjEQ3ljP8lsLZenB8hmpmf7vH8b5thY4/6Mqn1AYzxAvDk0BCXvP6Uo
CZEIPpx1tNY92IRQFaENNjPdBNeV7O3UDks9VOTSHKrDD7vq8Ag0ULPz7+bhQsTG
j0wnr9Or4ibjcbLM+8jjgt3NKI3TAkg6WBYQcFSHpAlENKZd5VJpTF+0nP06DBIT
ui9UHOgPP287venRmakP1hKEUyXsCz5XqtZhkYYpfhjK3LR/uLiMM6/CtO+AcXs2
NVU0n6zhlRrr1O1HC+86WeFTp3I+LlrMxuXHT/FufMoc4Al7YiUU4XNnIFoEnoHl
oorsBINUjsV9xm/F4mB4u5d9UxJLGZRxpI/WJfjOoIGiv7Tu8/qLMFsPwkx5+FlK
CvRUc2WAF9QANg9SO8ejTTNEBufTQ0CJilKPTTsERTKPUkm3JcWoHNcHxi81OaC2
G7Wxh/acpYEQywAbvekSOg1HO/2oZTLhHTiOi05xptX/wix9L10JxYWNxHzOyC04
qAUz64wN85+iD6vNm8XBPwKu5e1ECTfIo5kqj6zygkWeR4qY1AbLwT4Ci7YFkLj+
emB67xJyT7oQ9sXj7cOpDYwIASkjxX9SpUjYzk5vueIelq0/Toaso+hB7F/LdBDT
JX2hTFw6+jAuC3IgevUZ9oON0zqVL6HExzZUPMBQbiv/KqIVhwdexknnA+urKUUp
J5MoJpRKz1I6caVV8pibM2sT2LVNuhKMwU/4jpNxkTvADyEtzSwdUiI3bEXA4kBa
lkJXgjyIYAWihclYZfp8spAsqKCl2J9pfnbViOYQsqxknnSKdofz0UDzItkXqdsq
ul4sFljJCJKo07PqWx9XvlQsw8iArJmHLp2u5mqHpNebOcS0WBEfTdmfEpikNQYd
YYCV5NsAWWl6w7uUY8EsXVpmx4R1nehWwy39XW23h91UaUW4dKNIsKLIlswiCtzo
SfM2ad2t+134lfFDRxQVQ3ipPDwA9B2+Gxt7AISpZX6V/dtBU/mNoTVnVju8U2sj
yW/eUBHZC1Q/pBffg2IHpbFNsOqX9YCfl3+iJWIzX7OMkiDzrcAjNddyd/GQ+Hct
DyIt5lmESVm3c8r66a3Q6iLT/xwJ8XunNDUy9nZNTTWJ3eKsELq7r2zIpEblSRuw
zEXPxqpLxNmHYnxjcz3/UmZ+FAItI+6Hra0OrCySqkOrscHEIufPiBh9TruKaclB
o+m+cz9lBqSFHZ6jnrG2SHfcJqIPezBF06+vlWkRWk9+9+ecLyQiRz78hTn2YadK
kycPBjtuuos90XFafmCc9hOBcEEkB4iskCni/jxR0sRQo3WJebLyGNy89cjyTJLn
/IXw9JnSe8wdDNlxxI2/PZNWFbIDOagpy6PfKG2/J3qphQTWwX2RW6gbMU7rd6XE
/9etgaEVaTxLKDKf6pc9sESnuAYyBqe9REC3q5IpqKCgv4FYBR1wn+RoDi67nIIb
f9WJKV64onE3GwKO4ExkmuFuSZNFx1jfA2hOFaiKFatV2DYO4TsQNJM6qYCUa2Nh
CUoDSZECWBy3uGR5QYULQ7NB7ahZ0ak91gy09Kiaioc4OYQ2X8aFg4LRts/qbtzc
LLkMq/wqW+WKfEe0gO9/2HUCuQHl3KfIdYYk36CPyJ95lWw4e1abVFAvLyNDOK4o
QcL197F2b7ccnvRyeUF8ZPeuWwnc6ABMaqEGd8cc/jZSSyENImu0SNZsAV6LMYdP
RvjKC+K4lz8zslOBTCaVXBaFsvUc2LeUGWNnQOQfVdVojl3tKgmIj8wOc3cxOPUD
9dRe022f7AqgCxPARKnmkVEQIqj0N01Z+ht+QRAbh9PYoksR3hNnsnNDNs8/q1U1
g1yv3NgNmcPY8IUIeHcudgcIi4zx7X06dyO/lFcTknWiZnVHsNXyx/LA+oEyYPc3
kwE5CLN2IRgaxf6CZW2ysv1HTXFE6gM4cJIE5gwDvWQ9Pp1V6oJumCIfKF/+Alax
ezkkmnp+AZtZLoVHjV0EOKnEwNCCJ6RFr7w7UjVS1opPc0TY5ErwHNNizs8ITWG4
6vC8H21Z4vtSH3szDmCstpQ/ODBhy3jikXmHkNfj2pIwK3BfaBB54XuJM+2vTwd5
qRIxZHPCTP06ByBxjXibQJmdh5SEqTf+V2nVqtW6hv+eELLkherOqP251ceragMl
PaoRvWSP2m4aiMYAPygjaSfFb/9i2XKEGQR8t3YPxYWYq79PuW8Mu7U0JyHxiKgW
9pEuZc2r69cT9qCmxkDEzU+qIEdmXshSa1umU3FJSk8ytQsWtfW03aUxnObxwmmr
7Iu+CDYCsz8o4a3YWGz9gs2qxEIrkL/ebSMO+62JbZDhnGXtirsu4gxHhnbfKfn5
asE2/kTaeOAP8qrleFbVSFFFqtGXKULP4p/lroGUo3xRbUca1ex+VWIQvYSl9UgC
qzxOEoN0W90ulPY+0FRbcoNlOhnUO4OgvdefoVeAcvfsLko+AfAwsRbPNtklMpgG
KdHtXHku9I3Zky/G+ILSBU+wn1J4J/4gltwRNqrHQphZH8MHROwgMNSlYlyemOy1
4HQRanOSFwIk7bX1KzqHA0sAFY05bly9+Ys09mxo3c81ybEibgqfIX82k57w3Dmi
0zy5q035ze1WOTlBF9hDkjgIhRpOk9DPepaMK24BsJnnbipfSVMYbtUxtklqjzsc
jNJo7LlKUtJ4056tF1IlTwre1yLSReAb9txh4EfFSTkR0hexaURwsfDaG2Apx8L0
D5bhW4qiqd/FRhUPE76/v7nzBl7qvZNe1QGoJIEN4n2F5o/vdq3+Ihlj3ZHQKlBd
Znc1PlviKBu6G1rYMQXqtQYXuOmYsSORchkbHBFWVuhVAkHC/Q3pW7bnfSlmr93O
FP0/hIQL2aeQp9eyiayjN6kMsbtWRH4+6DAa/IngN6yS8tI8BjmDU9zL+SFX+nWO
Z7saYpjov4IbIQssK2ImRoy0UJdvzQtJbrt4tdkKPs+iGVrVkXsQUtEp7YSXB3F8
PQJjLElxQMfinDdRMSrkNWwniZv93y8BAm/z0TFT8k3DAjqM0t34XYLad7ouwBkF
ZX0Q3i3te2wPJrHJiuQaHit+Mh3elnpDf4IuEOYJZmVyedQnsQHK64Sfasm47Dzv
Vi6gdJS/Y086wLyJCH/1hu5BaoCpgjpMyxv/VFnz1O6QcJlieXE/t1QRBQ6Pu8oc
Jh/dYHzIg1mfGgs6iY4rA6hWpy7NIsBFuBfhHFluzvWGYXm3cCpuyeA2+BsSZzrN
d62HlUT5lyUlrd5U9afYuep21DfpW3fKyKa0VLY/mCAEp0QvnDLGev9QN7jLE+9W
zPhrn5BBqf1mz4s0xiArpUwbVrzo7GDh0NL95OYw6/HE32OjUy8kEyd7d6GDsF1o
sku2KV6++bdN1Apbc1TcCxwW8+6q/4w7KngDfVqauUf7IOXswYTwkSoNNlHSendG
YJyDxARDPZV0hQk0blG4QbN5BpRi8VhrxEBK2iZhcem2QtlrgwFpetJRlvij/E++
JTu9diHwi0gE21A8FkuN9M2J+KxO2dQxfjlKBzk330Khjo0/gWaHmUW9rH1Ly3ex
Xm9FnWJDJAgCZAE2fsRjpChdNGXVArzXE1KXv7sl9TBYfLTQpGwB6/Z8pGNBF7Sz
Vb/dmD+G+lt12XKM82cYeh+uekxk/rmGCia0r9kQLel5B/LjLL8J5iCJJzewoLFe
Mako/s77oS/5E1MKSfn4WDUpsGK17XqZfcaI8BSko/a7o+fXGWQ1vlxxOciT3FMp
FczEQTe9OwlgjpKMOhoo2zF96XvW/Xvf8JlBKf/Zp8iWTpB9gjwNhNs26uqYjZJi
YadauQVlmMtBJJVcd/Fl7LI8Plh9u6Er9EMVEcP58CH0NRMIMMVyU6JjsG3SkM+F
T+AZrurMUtrqnwsXFMlvYMPEA149rOVCJU7nQiNj6GjCh+dX1OdNn8whkAItcwvB
xSM9gDsKlRI0IFXFgiAHWYxshc2DHCuUaos7LvaWUY0bhQ3+3JBDy+hqL+OaB3wp
dZOJVBG5zocgCBUugc10IgVvg27G1BG46cjpqB3gC2GIXit5gf8rVWQNyfcj9EvQ
RW0CL5FIpg5NdKXhOdQJYvm2hdpG4hQvGG9/CbI66HVbnJLr56nwn7pvOjO06O3u
Wt21G6rJuw5SI4X5IdfJbVIkr1eRzTwxFQiIm8ql5H0yUbE2ROUd/1ZeKaTrff+d
qmwfBPHk2to4+oEccsSUsW1Zha6QOOJ5C9FNGrYpEAMv0tYj3RC/YASgZxzqUKT7
R6HMUiXSHNYRPH8PlLUS8uWSRSmPrXg5KO3OHkxehBOW1Xo5cT2DqQZscaJP+eGU
8oHewtu7xc0KC93BUIqM/hbbqVcy3JfpNkStTmV/z/Mg6YkEF6YQwfr658aXHQjo
o37PGq4xHdiP+oAi6z/rYBnjDbRqHke7mAobgvvPAJc8RTS15P2SF0NgVjImng/+
UegmRAekm+PGMlzOz/3dQNG7xPOYha6oJqi4HT4q7zXm1gPL3R5Gn7CW4NhI2RZz
MUz11X56/wOKzqrcvVohwsJYEqM0PQCnDjRFDlxYkfWuWsgPCVApPZNptLUQ/gL8
yEe7Bg1BmyUiGkRREi4zXAmKxTZgW7t+XZSJSZOIi9xS+YR8MaaL2ElY+WbUG5PQ
KjE7loNHY5TpbvxzTG0xyNMBKnoUuDSdDmvbyOOAbjVI9bwjas8CqLUh/cmUriuh
GF21Lkxeyot/DjzeiPKr+/u+sIgAgpm27B3tv9EIfLChZ1U+nDNZgRQR/811dsPq
dboAJH0yMZVkIkzthv6cWAzeqIcGsm8BJK0tZ5iBz7islMKYkf1BMnfjalnRekyJ
W1VqWnNTTVxECztAEr0DELAd/JLRee+uUL9Si0WuwT1qqMWDQAftHZMNtpmFx5px
2opYTc+yHPYXNvaNq3ECwBmY/rRlGlkbGduTVJP/l+0kWhSPcnXr4mmU8Oj//uYG
Jm2tglYl/oUiWFsAN6A9aeBEsomK86Ii8PV4Egj4G6GPKLOFPvtbEu3RoAudhhZN
eerkpg9IEO7SL5noUPtdeoqH3htOg3lCm3Zohfcfs3oXffWgizYZPqzj8eEfrGRz
uNi7VMQVWV3eC1x+qcazkCtfyRCIWXH5lV/DlvlcBUalTdZ0mQSrxj+3AK54HvCV
CL8fiAfDeOAPuuGYa7TlLAJKvaMP2tsmsBa+KF0clxvk9WkHEWZ1rKYifbo3AxPd
9fh9tZaZGkxBssdoWcnBiyDNoG5f60qCozsg+O3gYJvpnmNoQoJUqEUu2SS7RbSW
a88j+we25QoO281tYlGhFymYTBVOFUPXpQry7XEWCPodIBJdy53ebHfmdkI60lUZ
qarR5QSEnHLsrBFf5CHm1wbeup/ccYftQIRb8wMW1URUwIM/+jh6qYpV3FPEw7dC
YlpH6iUfmfEas75+M4xEOPlDdW9IhvhGtt4HGtPNKMo7gLQcN2Ba2HJpduwhPeDj
iRwexyXM5iZ01x+3/1WuZ6RZr8t9HsyaiDU4aLaFcOAmKT4WOdTkp3ZDZDVx/QQL
OMPUciksOQEbVUK5OKcKYLJvAcnfkV/U8k0XDlD2EuyoICoi+XxcWtYK7MBshjKH
K7t3AboASvD/gdzgRT4ARQRvlUGoQBsn7MbwIcMpGNF/S/sbg/ViV5D6fjlkpgOZ
v9KGb+2zaJsPK0nit8XPPxeOjVPpaAZYn1GQbU0MrmxBv4qwnYY5tJKHl05sc6Tw
M1j6rufB9+dSCoZlG19fZ6qTdt3TAW5JVj26kIbQsVdRVgJQ5pO0wiB28CYdPhWi
KF0lwFt5nyQdTRIIa3lKd/dRSqxNyMxs2mmU4BtbjaXvZGm32B/s1Xph6xFgfrnz
V5fcGVjPRjIP2zV67cooRxrAUvuaOLxCpPGLNh9Ob/7jXwtuD6vyQrAxN8S/kl2o
DJ+JEYAXppmy0HmkSUfWzNQevk0+WNHwXsplgM5+rX1DbT0w46jHFFAbEg6/fC2U
lxpUtkZi0XbLLSDuJsEoQOhYl+YetrJ74ZJK/ZPknaLo4rzSUyshfMzzvO1VkrNl
fPZyJe7ZN3V2RgTJ9tC2HNdw5OQC+CBHAL8U76Z4OwxaczrVRET04JctAP/eYSN1
KcldLb3T6EFTq0CvY1TTK5cbTiXU2ql8n9hh/z8VhAI9Y73W2mPXsTZ+hUZUI7fj
ZkIaqS/YHLMJylNRmRVWcbFCx9ytD36nB5bDMz/BfEbFaJgZK4cPRHCxg26aQd/D
eCmpegLQxQf9pqbJY/bh1b4zgKcTCnAbzAYJeSgppMcP62U2SJFmRfW+iRhMYRso
5r3vnndLHAN+P9bCNqZtnEx4Jp7+c93Ja24rVx9PV4Cur1JPRtutRkbYYP0vwmym
ofuqI+UZ8Fmz/4igq00gaAGFqO/oUCPMJ1BIIdeskIBs2S6WwH4D7bWaBmcWxKes
dHOmrjUbqkA5VZi+B/f8VWCrAsV9WcO6D7AF7k7VIuJ2sQjJn5Jwyt6ZHBP5fNxp
DoEVKzGJGEfTV1ELoqw5EfsLshp9NYPRecdqytB0h7EZPYf1vMglMyoMz9/MRM6F
64Z94vFDVUhJpBa2F3FY7tvtmcZN/j6uMsXDYUlC0lRs0i9F86uDCg1cenodmUFF
qPEb/O4Uj2JUf9UMhmQmud6FSuVJDtfX3fVNuLofkdvfMZIWNFAvhITQa8kd/oPv
SdFU6KlETvau13mATZu9w1wUR47zhVpgU7wzQTgtUK7fwcUw2Mhwe3pquRYYmPBP
NpXds5TFylut3JZz3xQ3xOcH3oQY4+xkzcG/0OSmTzxPWCvSIV+zvMJRzIidZvXi
vxirnS7+6gx43ZsHbPsLf/Tku+pFFi4b82rLY+OOQnez+7l8M0J251ra1WW23VV4
34tg+IHH8QH5Jk6uCCC52WwrwfTWJWwF7yDWbI37/Q+vexQ4Lh7+hMAnZ7NbLEjL
smC7gaWSRxt6STPTickg8Ar5IwnSGOWYgnVm+xalmua6GUe7ryxlB+ElBCA21u6l
PmL7rnVU/K20BL3838F/kBCFYm11SY9i06tuVyCdsabaPh8CxHPZKiknB/fH1/F+
mlR8Y/0SjO+hmF77CybWjxf7A5NbBHrfddTsUa+0Ad4vRMHovgrDBxt3ccnf9hwe
YDDIA6oWG4TooNoKjqWf5Mdry45Eu5iiyYua7nESJtSrhH2wjb+DITKIn3b92etp
PM6Std1F/S0IbDRyZk1xtf7gS5nkJft2BOPiX/EMCU0Cv9AHKNznTJ9dzDSKcZzA
PPXUIulLFWzEvp7zMBDAUA0Bp9d9NH2DTgD2oXJghBjs2Tg3rVr6O494P2xkXfsS
U8N9qptp1aT0y7D0H/9d91r+06qRxs7+v1BoJ/LRgx0MQIkJsUDdORwdIroAsQZM
8Z/1BdzsfWj2o5teew+m+98MQMJMQKTn0fxMQ34ULBkzKuJknr0ICCEok7E0iPSO
2nj1YRxJ0SHf+ujfQBh6rgH9ox6hFB5QZF05PCd7fNCeMoUEG8Jq0n2Yfz+RV1X2
txLPgfpdZymXLPUWNebkeRTNaDodrFBHdZxQWQuGRE0gfAl+glbnfa014D/Fy9/n
Isn9sAviZkQ7rFHWwi2hHsbuyD6nBxB5RRsrLacMbx3u8yiS9VZ9DwLNGsp6/NfS
UcARf3NvMaYzWeSsGupoCfWl1G6uIXY9kKR9BsDWELTUleXF6TiSE7qHbbXO/nLD
dvGzZIbr5RAWPu5CQcTgXWSpsilEX0PmPF3QGb6k6rarFb9QbpSpmR0jxqAvJXCo
jchnkHgwRuNqDAnqEHMYzegQB75BEH3aLJB4v3NCUCokvEvnfJa9YsOqNmR4WiQe
uqfFX/LwaUoLe/r21iK1Ro6nyL2L0j7XPcUzL2n8ukfAcCSJB7zkj2wTzTsO6h72
P+ao8Ybh7ulQ0aWSdSDp4Hom6WYDu8HuPDrS64OH3RP6Wx7uWuUL4j66L2u48MnB
cY5eNXnhj6mA6qJ01etZfwCE+BYoLSV1JNMYXM0tUGpKn+bLohFTVPYa+Za/nY9N
4cA/U7rmkXY1viwsUUIU5LyG6Ql+g/400/PRgzlbXpZmoECeyhq52HA9+qbc02rk
51d5f8P8KWxhI5IVDpr72Q+zxRISNuNMOv+ZwfYYHxdiXLbdlPsuJ7LcwSwE/5b2
ZP6YkGzJUzDPHATrNIohC5lllLGwa+DsBu/XTEVcHN0zqIIB2LgZj/YMS3qIw1Zr
8t6OTHlSkcs//krktV7hv30isnc/eKovV8Gu7WBj6WeKon0elKoSMvWiuM72Tspz
OjUWphFxqntr6hNJBmjIc1q03xa+pG9784HKZ3Rd+vZO3VtpU5YvwSzLhKHnJylp
Y8ms/MQYLzNDzj6aM6yLfPm1UcB13R4H1EUoFlsu4xdtMQX1Ym5oFTbSgtHi9IXd
tdlzxaYlT/PSAdqmMH1R/aG3Mp3n9lLDFq/AypIzWIKsjqTQVXkwgK1sFXS8jbhz
2G79fZpYvgk0P69TtTuWoovRRncL5hCMdHHoCWVzBNu+M+SV0Zt6IpDQdGXcVizQ
IvO48j9CET71VvEqdvI+Olw5Xqe+DIsLbuTAJ3Anshrrc9PeraGoH0eqtnfaFEfS
yMwH/8iv6jRLsKFoB0fxbjgz1IeqS+v4owjHRXYO3r6eMk+H2FxwFB25AW+VWxbr
XZ832Y+FvhKtfB/aVfSFpEBr3au4dAQpuFPaQ9I1dIQXkUJr6Y9QdGGfIhEej8tm
jkjlm22NXuvKwgn7NPRs1qInZKOqn+vkimRojUPiokuxSXV4MdhcoCvhFM45Goh2
F5iTkF6B5pZiCrQ41cDcWsfSyDGb4QiuI1Gj4n8QMd32zjd6YQoIHrh/b0OQvJGZ
c3zq4cD2eMwQXjcKRih6bGPoCxhmg/7UHYPEqw1uwXO3XPOX04E9P2zuYsPMdGct
fQnJwjCXQgVyxFh56+57I8/5O6q3C4k6gzZXwM3si4yzeNi2yOTDlHbkcrDsgiUj
cMi8WxNu2ewtuDO6pAvTQw5q7tu2qfSi4kUMuSz7AofBXztSgngD2K/WHSRn7wzd
1UUHHQg/mCZ8qyISOQbjqfFWw+tC+icBtFB0GKlrbEYvC67moVZkfaB3s1uD/xhz
Ear007pmB30GBJtdkL2KJMC3O2k+eNO5Q3YP2NXbdqM3uBiNRF9+fCRIq6UXviX4
wFAKubiYKAWruKRr0NeI/ydeZNKQXZ0p7brCTh8Ewg0HVAud31HODKJ8yOdqOq/0
0g2TFtNlpJvnxiMZMcA5Wp1w0Hd8VZUOP+Jh1JcvihmkpD79TUd2Lfvov3vIq6bF
lRZksCue7YWUEpJn3/INpdi5lYABnyf2hC8NNUAwSM56x54dHlmSATPF+eyzq+6n
KUOEZ5rHjVFng3x77OmDJx0tw4GWC4ghAkURFLTQuR96k980jxjWvzscDVb506az
EejSs64bDB4CMPF7XH5mqP2QcAO62jBVxcYDpQja5deK2RBXFiIabKG+DKOuz3Ur
6tUkwpyMe8InG1M/5X3kur6OX+wZS3knrB6W3LizaTHWiZLmDNR7kpfuKG9FSv6j
f/UjvU+E0Eed/4MId3FOGzBswPzfoMHPM2f8emrX4yF9cPI9zp1YdjenfMEG2205
yK3kQDGshflqNx1SzkJ+dim3kB9zz3MavsFmKFYYg1fmKS7U7JLMHS9XzkZgolWa
qqWOFJL8q+uUnqVje30YG9pyNFYic4rbQ9JqumKBFu9/y7uTB4gPrzzKut24tx+S
34XisW1dQSYzS9yNYgQg1AV0ilXVEAIYdHZniOipZVuf8Lb0GRdkTrYH3gjjltyW
GQi5MG1q1tzfFYhSbAz9/DHzFMD8k5iw7bSRKt2MVYi015uSJQWqLNl4+7p77edk
hYn9LvPx/pXp5UtDQ5VU9wWz7yfprxhTswWGczEDRj88UECLV4vzIY4zxW41Yldf
YL+NUT+Jtt0YVaCymRWIdHOiJ19MZjbHPpdQ4Iw3oSTAZ/V3/rXOns/G6L/wk5ae
aIuVpHx45Noddb88G/H1rRLNczCOG9WiefSYiXT0QCEEcTTB6Cq48z3s9kzKtPdQ
o+bCoJE9uKESgq0gyQ4MdF6ABfM3u1gB61A5bXZ6yG0Szfr4EYBmdv2TPT+N2CIQ
fz+9SIPacrBEbx9vf2cVz2qSXFamB/nX3PpGmtyNWOlNdnh71yaTxMuwqBD0hSxg
0Wa2IfsKQ+41gIgPIzIWBaF0CP6fX5ozoU5V5VPu0NJuHVHqaQFzPf76YTx/POdN
P57To5aJRX5xlESQx57ORGcRP6tIzCz0mJfHp5DO7xbJplu98NwQHFCqAGi8QUjM
u8sg4XyYJSqhaODRvzDhGuOp4zq4GzcmfdYs0whG5jPvevy2x3Fg4zbMgD+xoRYe
BsAQQANixTXgLmP8Qjcmb0pPsEVcb6V1pZ9cFzuC+OF12kbesYBgSExu394QUe29
A2fCgKKSyo+LPeVrnBUmGfP8dhNibgulJu2iNarIgTNFSzRY6jIP1Eu494jEKZLt
p/AGJ5y5pqsXer9l8wbt+tX/JK1IfEcb+2XwUxl4jUyh3lTL+b40PNDBqqHeQQ8K
OC3HT4uyW464R9Fr7zpW6uwPn0zUw5Zxm5dbZ9/3mhcI0M4vVBYF75rjaGFICrI4
PfVQzE5GtkhmSzfFOrP1xOPrg/q0Y/WysmLuMUIsfyy2KdlxF/TlPi4yR1kL2bWo
KMxjcsCFiEQ/0cuf2gpGD13SI8jiLjwzcZClCsUOWGX0lHvCThWalvJSYjtfhztV
vX3DTb4fCtPc8e4d0/UA5f8xLRSy82F0MJr1KVozGpCga86rXmu14/ChH0BHPv7N
t4bhuLtYF8m8TK3NUT1f+eUlibe1otU9+jmSNeayNaV4fr5veGDq4uRYklJfuR/c
pTOEeLwJC0xgjLqWK5cKMKcPlsrIYTrgaAEwALMThRhebrrwJUg8qeOKiMQ5+506
nx8fMgIv1obYiTsAjTpVAYIBmt7HygWGzDUccXxVxIjy5YlUVFBM1vzDyEusCIxY
cmwm54wSxMDnszlawxLr/EMm22LYrNTTMG6sQWzcsNVnKzSpRUQHYKab8z3So8xQ
1PRA8eZ6aL8sEqYiHG3qjQvIafrYC/PO2oanofb0lgDYsRE65PozqDxFZhISVQG2
11+t7k2k6pJFfa7kSywhwVjxFklF5zlB39rUkzlwmqIq/FvZfH1Qhb31iH1vX15c
I9CwYzJ8iYeP1Vjs8DBb6mWfg5uli27IWwnab/mOOb5ezzNvM6T3VuQ9xunjgQAL
9dAXLbnS9+/Waq6E7vgpMSfXxTtdirLY4szdVedeKts7FfjdVgV24VP0spAiKshO
9GZqGJiDdf45L1a6AT9sy9YoAU8kvewm8f4tmdM8irfGqdiKWrfeR+1yg7Kx7J1u
BT5bBMNLAXfCXv+tT/Lso45e3Rr5zaxnueiebtdr2zaOG2++7ANiHmaw8UOk6MTN
xwR1UjhO+0hXigvRShlfznQwzCa28et601PA08Ti+DNjM/SUJBSMgET8pDRjnotC
kM2wwKeeSfvZYIj3V5JmbAIRRQdaaKOg+6izJs+uyJ3xFSuEvqIkT4HA8R1ujL9J
I5vgD6v8zsy1bAPACwFzsSpXeMl6dIXSzJ9EZkcAswx60YzmRNDWKp8BOL0Pkzt/
aj1e+Suh7YMppKxQbU5fvepMBE7BbYKqoH31Mdr2/rlrrRfJ8uCIAbMVMnGTSJ/s
kj6SIlIDr1Bznh/MslNeY/vzETv1yELbEmu7tkQD4k4ppBG3OEQsLDBjBucW/sVx
2imXU9ihDIwkXmHbnY7FFD952F35IjdxRS/GByTuUdvnY11UAXea4qz7LtkvN4yt
0m6DeIHSriZMZd/LFfDeNZ8l7iZ7gWw50U3VxZywSIzZMdQ2Zjnk5L18qzs7vkDJ
WC7fT84QI7Ghwo7GP3R/P74nb49sh6+PjnZsiQlcgEHjqL/QFSfNEQgZ7jCl8KNi
AItXrFBzx/pU3tC2drgyGFOsKrvS3pOnE8Vy0EpgdvCvveBSdgegRWuR7nhzic+/
zrN1WO2Y4qoFprN7uK5jPZY9SMML2gUmVNRZm7pKPsHBl7nxV5RiWH9YfPfnhj9w
kSuyVMwFy4/7RwKjVX9bjutfAOwlSH0GkxC7e2k057C0eIy50PR+aWpcZELPJ0ZF
Emee7KbStcurYPiH3Js9bt/6uX4iYpvy4KFsdIJtt7eo/WkV6WsSkuFzF4vaim5R
Hv/XvCG8w1pjDeC6Vb7lYv0rg7us5bWMapofF8Tq6vYnd9Py8FPtS0ffw9BCKYnf
kc+gOsP7841KrxITmElHq3sH1BNiAqFkena/KwZyvx1EQoU4BJr0gaqZd+NXCg6Z
LKcJbCofF6XX4yAx3xTp4/46mF0Ul6Xf6yo+L92peSZAXF82QUpMBiruZrWmURqT
hSowlAbqiBFts5QoVvrJxB+9bJIhWlFOVGEE25yGcFncFyo77/VTZ1sPd5Jcd4gi
0lmD2xGYHueF2MoIRE/UJ7qXCZ/Dw2Hg5f9j3v+vFqJiIKQ2uuPVwDgS5p7rPvsD
sIK1A+DhEMYIUoCq9Thql0Qbq/sf/LGWghnvCLRwmMOVUX/uhSocwT/SVYyULGx+
EaZHvfq3jIG2lUoBrlbv23upLoX2VP27lQ5CA0GCoo6dtYkhDh7/32wHcdifJRcr
VRFGayymiWL7rNxMTuOfGiCrZZGlM+IE1Tt/SLe/3omcrIL8fpHh2Hvhz/Z4uC9Y
lfSeqYo1+f0UnX6cv/ybNN0s6RUsshgpov3XJbA0uxImxVBBLRXBQUOHhtugow9g
gUoexVu8hYPAiyIlL0h6ZQakNiDV0AxHYToBc2rva+Yzkui5M/GZckTzITEG0tFe
9D3cEht4C74KEN9I7pfvXIU8OErfZ3jofgK3zS0RNPad+LmCbQmK5cDg+cQSaubU
2TLCNq2CNLJ3kUlAhLNJOQ5x0CY375P2yy6vO7PBqua5gKT4YS2DPYd3326PL3hz
2DtdWUKTgnn19NTu3acTn8Mca3A7X4Wbz1uk0aMR4AfMcWOqVZkY82dgJ1pKTTT0
VBTYEnq/oRhE+dhXj8evuxp2E4Y84/3/dIRtTDbsC2pmpJzurNGa0sIEPsrkVu5+
1HEqBJOxdfO+i0v5LsOZQReV7nPlaWVmn7DDnSh7ECsvC3/UZ9fK2t2gzVkw/nBS
hegksY2ncHiCC6MSs8ZujZHRFbbeJU4sEBHWLFr9KjK3NFrdhLl9+ybjHWNO3FrW
LrmQeVJSjmOoBKfI94iVbRCIzcNHRNIL9JxoibLaWPDosHyQ8K+RHlMBt13kVJC7
ak5k9cYqfwywY+8KF/YT6gJ76PpOGraSr7Sh3TzNbRDHsO5/GUvicfaGFlDcx6LS
1yU3xPbzUmTjtfQfpS6ZLDvC+KYfS16JOxnwGTn9Gx90PO1X+gjIv4mwRAcrwM4h
WT6PvE/X9jlhufEGwcPgFN299t3jhoJIpRPxWzVV44y+aaGZrPxNnQpFEq1dXzor
nCL7+WcKO+nvU5Rm5BPEygev2Oz2qsRKaoLihcpbKV1+qZ/ButkWPe4plIMb6mmo
eDRHOJyJswZ/FTQKXAZfT3LCyxmKCTSQetLCoTH00oi8qqlZlKVj/nMR4K3iVNWo
lsSYDVBIcSmxSrlFH3KpHlhP7a4wqr5wqiyzEJA07Dtjvj1l50oXrFxow7XEDPU1
Slzi8Hy3i29WoPa1aH1RJZLjt77Rqa2d3yN+g9F21m0AzuIjnssCp5EEr4mw3AkX
vnwNdSitorfzvoB77StpbteAdGheZJl5ia4Ev8BASF/fO3SAUag4GpVWC98bEV/+
pV1ooAIMtEVv+rrlL7A89rZ/zItJhTQaJF4ceEBT3egp6DXQyiEcIObMnLMjsxp2
fg1cWrxwQQGeZ1339XFWU6WfBg+VXYGSvxntJ0k4eqJTDeUEZi0ZDQl+st9nvpR+
lrj7w/zpaND+YBa3yPOt2AnPelFFjGTBJQI6V4eLJhBvSgyXb7gQzl+TjgyjPp13
67O6igfqBtH9amp3GmYDeZJI2/jp9nhdrCkLe9aLBbhJQbr1puxh5epJB179YMXY
jq3UCDy2P+TleqVfq1l4RTDJm6v2k/zXDoWiSRmfaTmYZhxLNuCc+T22g5rJQbnz
rsftyZcJKnVT5F/PGeWtlnUzq8uTxqFAeIbfUc/yl87dPnwAKcU3VuBqA51AgiwV
wrAzAWfrzHbFQfGvY1lSibgmw3hNQ0QcMcve3AvgyhykW0AjAAzCGuTeGPRO8elo
WK5vW2RfHCVAInEb+RVpbZwBQCbpua4qdcIkdAXeYjkTPeT66ldwpalHMgPJcUlw
k6fjf1O+QwdYCkGL3GPGO+HnG2zp+O9Yc1zw8bm4oZ6pNFcik69Q+SvT7Q1m43+p
ocAOBOHhjyPNuOjtmjGn6cukj06NfTxwBA/GdcYnnKu45sWZ0EOnwH+cLH6W1DZ3
lTJBJkZTq/Ehb2/WWQ94JRN2vmaka6tor1LVpqzdd1wnxhPAeUImCQMejm99GdGp
He53noqHxXc/gqiob/y0jNCX5tHgZ1u9NmTXt/5XLHaLC8Gqr438TyMW8bGgjbHE
SFdvXXnMKgp9pUWM1Fn5IcZR8ZTgkFyBOOuRcrEkOf4ddpC1XW8LBHizsyJ3NRLV
Rq00mZ0d52Vx0ZPFs0XQfIV32ynjtBZtsP7GQf2y3ARGq78/INMDuTyPyq5DOAsm
w+OCLczUxM+xCDZQSA84HlHLiiabKuLmQbiyUVp08kfUGK+CI9kRSC/d70FzHOLr
C/eQS2TPO9BiyuTVRhuMKxVjx38ehBdAu0qLYpOZyL3md4M61i+aWGuEi8Yb3edO
+sYu++o/tjhLpMeXsqwXvpoqcpPHBwLBJqw0oVM3e48uapqAu8zeni8d1tvT2Cij
ucpBluQw9I57PV+tDOFrfBJYAs7x/KC58jFvQS6QLsUTUkG0nl+8qvBEnnWzdOSV
AUsup8VhYUoNW+iE2BrxQLAB/61Kdtpj55M541YTokuwCYlcJb6jzBFQrXAT0eS7
IDSME2sZgQi/6x4pMedtfq5rT3tPGsvy2uPTXVUsVXFdeS7z5KfDgWYQDPvzOkbf
B72N8NMF41g0vm+1ybM3VIdvR8F8vn88JqaV1Og5IvmGYdt7eXF+KyegtwwaZR6b
0j0IRQmbE/UPHgqh9ToK2wiosBTr/CnMWbDjAS2GNeJln5ORfBac+yNsTYoIpC8A
KgOP5JWVY8kfo1clqM6xXCe/cL6eTyTKx9UIPSexmKDn5oxTD856DuulmoW/rATZ
k146eOspNbKHqtDaFZ276l5XGfHYEMcYtlZtDQ4MXhBIbkf02B2o6TFMZ3slQkJN
yABZmEyWWDf5dcmvYnM/I8QMFivS1eH6JqhvLdRcbGMTWS5rts5n7TKfj4LudoQ+
MiAwvjFRh8RmV06Qht8Kq+E99TaNvncKsaPm/As37SzZA1lYZNENHRtrruml4lhQ
lpy51gnyNbnyDyUf2vu5H4uE+ZpGWofi5rettHo2X1668O+sD51I/4g9ueXGYlph
wRPyN2Lms5YDL/9PcWROOsQ7vaM6EfcrgUP2pm22NDWc2T2zUPCGuZhxd/SGxEeB
YnMPwtXyjHV5HBvHgFn5/ctx9yBGOxeXlPV2HGnF7CjQD+DWg172VzZPp2N5SER6
kCAmAAcnzQhXVgGg4X9sKyfkWEKhfPtdkEg8hv6jqBm8ar5nIIFGgbrUPYmqyFfY
IvkIl8YnTRAbrCME3ZE0j2j2kYwcSl0AtmTuf5yvPSXp6b5zxRWG5R8xGhOC8T/M
Euut3zS36MEL7Ij16yhRQwGgL8q3B8/Wu80s0T0zYuHynSlB5Ae551pnLDQfYbb9
9ZzQjmZfzyjfZTAVA+wTBaghEtjSTKsZ9w1wa4NMqhqNkPiZXiZ+F0Czu/dxGJIX
AQKyrb9kxWxTaUxEAOA+c6TaQn7T05urg4ZI63qeV/5RxXN31C/CWXQse6EqgxMO
zhqmhiXkhTeK3idMEr/S7E6AiAmywB3k3dNXyotnzYkymUQ8akBTj9soluCmbph4
hAgAIPZc7GWC5VG4wUInshAQhMpiuBDXGw9uqWwQnbyVXs6NzEnWt0dId5nNGb5c
yrA+dhzVeK0kg8RriLFIYqM2b7QEIVSILiouV6ZZow4RFyLP0AbHChldqhw3nuvK
ocNM6Y3hPRQkxOtkeWAD4750SbIXyUkNKh/oO7fr0cCllpXq6q6ugvR2GReo0OXU
HLNTZ7u5KwwpwlZZaHz29W0tLaTUK1xw7NYtta03GaoKNFW0Rh1eqUn3uzPjPYsK
yVyslHBNXcKkH2n+yvtwV3WoxYuVZcvxZ0esaO6lf6Z44gNXQSNDwxSf59YVyO9Y
tDeelI5aSMc/6ilTjmetL0fZ74kNMtuAWmiqVej5yH+QB4j/Cqez0xJNi9L0oDpf
Ofe8lVR4Rk0YuNYFdnJx4muK/rBQMWmik70gLWt+SezWJ+Yo8kxAUcqXpW3UvVvv
zgcAAZCjVZPqawnLa7zc6sTT+gNDI2bES1zK1Qw2KZLRiJfmLhGuj9URnLCVryKB
w27xG2W2QpIAMpfzQHTwNBWnN4BPrXW4vv58J0trPN7eAf2K/ih5JFXdiuODYDWN
04Wgn5E0dWTv9MSt+/faEdZos4lhRQNSrdghhNEk4GhlLfA8Rn1cM4E3j5kx4EO7
D4wC4jFPPtQ2w+Y0vcBOLy/oD7Ymdd75yzrxjDU6Ha7dqE+MESl6izwFgvjiJSrf
jy625JPWkcKJlwRoX0WhXCyGEOlsMY5q3fFTBvzcJfxsMGn3AGp/Y2yiPsseMOpm
+yn4UhVA1/UMrVkMHeTKSyh6G4HmjPIAGSw+35LrsAXaegqfjzwdQAIjAo5dEShc
JDO75kpTf4zKsUkoWW9fRh9RWBk2R7Qa36Sle0wWlTO2CAvlAr7iNGbJhJhpVVFk
XBzGK7iZiqztpNtvreJeqNpEuizFMe3XRwM8tca2zOZJZ2niITRBlzrEx048zCQq
fqoxGCbRHC6Q0A856Rx4kHWVZiHUgZBQ3TTO/MZtydSyHhLFV2twnbbVhl/y/KcY
r9S/mZ1l+GzL1WWKAD6ANiWUuflmrHAp64O/L1cf6Ey0s5mos7FzNjwcRgSH20Aq
KpzdkYYEw9xObEnkETaVWHfGGeRAZce/JSZVglcBIm5fTGVgW3cgb54GiJGlsgBM
YJkh8362uFwv3RGDwfHlfmpO/5+0x5b1W2mTFg5FjSImbhpc4i7+RqHx2t+kSpyE
RmDVTsPUz17n6ekvVIn8jKdQo/vAST6DUesuc3WQhzxfIgkzCGzIElKXconoZGXS
WMbNc+O0WLYpZVsK6yXRDDxIeTGdf8pphCZ0SRhzhtNH6YJuDfjpu9MA1e/lwDvs
WgF5ev1sW0lHaRZ9e5cv+FCVixv3lZW0O3P496ZUDEshwVY8+lAg01EV+6R1itTB
0wWe4LrHkgWMIpjv9Yf8/f7KXwd9qdLi4yt/p1Lo/dfUMILjr7TC+5INZ4ysXr/m
vj5sig73q2T8xBLMHNwPFhOXHaPEYMzIXJvClY4pJfoNyVqAgxnoKdHRi3jANhOh
5VptpXMRnKdYCQK8u+AQz4ew4nL3U0WS24IkYRFcPqChl8PGjaqqIK+koYMZmgds
WMpN66qM4GHrj97j/es+py4JiR+ZXkm0sCpKG4RRrLph7slYKqGcn+VCxUUoFqi+
kAkd+b5njFS3I8yZWFNnlPkBoLpzPiGvrnhV82mOQUAwcOd+7qasQfFYeAPPjAkz
CC2eKEkhoyr8AEZqTRawb+STM9TblhlY4QY7qc967WkzIsCqOFIIJScM6F09+QKd
xZex5XImTSwBV7lNPkZiEdjybRx+GXy2EzlWGbvH4bXaUDSlQL5ZzmZ2naB9la3p
e/9gsedXoYCMlgdOpWjqsb+3vX07UfYVNHWFLSfy7rTeVhvZ8r4PiXs9XzwEH/+1
0jXqM0HVG4gSw02hxA1jf6EGVZN7Ft+LHFb+7wcV/9RUMFkD+CgWGYmQ2baX0Qrb
48DmQfkA3Vl/7qVaWUEaErAOnkuKK8PP+AgwLibXpHAses10w79QfGWKj0XjmBM2
9AABh712tTDbt6z3zXPGYkFacULoNzLOvhtjadyMEmSeZ8bzXfUC2gGuOxjMnN2+
1jLJls5VSGbI/SQdQ8QzVGElXoLoxiYVeiF6y+wrwaNLExo8jNp4CBuJbOLFbl2f
EBhF8UKp3PNm3U1R+vvPklk7UnhlFKPuRE+6j8aaUQ5S3bOufcFCzffDQOY5VC/9
PmdZsTXdKkgu9BgQP5Ov/suBzcPv1Yx2/6XkN9jpYx2rAFT3TOYUqU1Cznw3lDdL
rm6L+//nwNjYjuzMXI8QWBKDT30+ajwGeQ9n44RwTSRd90ED0oPAWwfLLw83Z8Kx
pz9dSzvshCgnRg/fTFLLA4sRLgn/KPYAHB9jsh3pAnLaiSYLL9OkBD6gbqTJKP0D
eV5h2/w4HqmT8vd9v9u4yg7hii//pqFmRcZOWFGo1sSHfcPCq45r4XNoFJ4tbPlH
sXyt9rx2hzyyuv32Q5ljifVBZa9MOZ11hVCxYczbVzs1hRTR5j0/dZ8vZKkBQh/J
/q5fzrlx7fGiccWw1/fpf+VUS+chdiwej+4zl7rlW7J7MCxA5b2BGApUFt61eJfk
UIVeCDulCnF+aEatQMVI2rPWRO8PBwc2TFN41zmUvHYEOHZ1w9obckbtUHmrcPjn
55IVxU9uppBS8lj2jZDQ30z7KGHVL/jUgy8hE9UmgRZUQzE9MGur8qJcpJFC1bvH
rn4vk5Q6vH3AWA0zuMAvRDVNXeJDupaeUNaMSlvBgkkr44NfZvEiWryC2XLOMNyM
qJJeQbEDu+FdtRXeDCIe9yQnIZRS48q/s4JuxA5fAqjnBp1lXQ1TxEviV85Fyoqd
CBsEesC6wHQiWW/uq1otFiFGFCDGIJ/DJNMjHtK9VigId18IFReI5pp0elZ76ML8
CqntTLSwxKSq1yH7H2Y3aLZu62Xgkkc3rI1PA5FgiOlHx6FSdg2C8c4FM50c9tfo
gIgI2LvIr7P1Z7dk7oydmLYZLK9VHLhN84kE0AVL4hsmsJaL7VcXzZgm1/BQpbOb
/K9HUlnaRLZlVfBh271o6IAUv2SC1z+ulpyCMfNWuEGh6FDCRHZREDesmNfgqAR0
xkgJWe0P6IIC949Y7dYK34Wzr4EpZH1EVICA2DZggQudpJ2cCXmp1SmENZpnUzoz
D5rvMrB1o4SO4+37O+IP26HO+qFG6YqVv7+E4X/hinvyIqQFGctSt4DDw70NNUw+
VsWVyGjCRlDuGlfpK/ByMxP11PbU9cIhesh3hwNOvKHIH4yns5bVsWKsFeml+i5+
IH2cPVwBqzqEVIcNrbat5RS5Bj6U2EN6/sRDkLydds2g0FSOEajQ9r6ktDtWsGGI
wsV7+0vU167flJy0FtOfBaoJsDsYFQL6C5b0HOvOembQW8Vqzlpidh6fcBvmcleY
01RznOl794VDOwxBSNaORmbYMW55Sm0TzQVXA1uJeeAa+err1HbYzgx5ZVhx6KbJ
n6U9W/Kj/KEjNq+NoJ+pS8z3lVDV2lH4HQk0FfT971YbLvElbJAia+Dtsyx762C9
GjINyiUB92TKCqcUqZGadXDQGLffETt+tR0DLYMgAJbq4oS9DBfWxorM2DsFfRMu
dJOpHaEZZ+aEtBDbv+o/uS45m4hjL3AMfdgxDSXU7PMMnmvmGBnaXcBcnEYPEmPH
L1AOTGcJGhdOUqZX1/BDaMyOek1iWogDliBCKRZ2KyKUNoQB0RasMJJT2SqVDqng
1Kf3nZXNdhaKzna9aczm2aZWiIse7wqfpXirj99Lf6nyZI/cUD0J5yAddgESBVI9
rO/7d/JeUA6E0ajM4mMySwIHbNoonoZl20EukmStJ1kvCQkvsfHGARZvm1N0szvM
HCB1mm6YOgBNKdpxw40ENw3ypb+YL82QfRb1eFazVkxwBGKVU4B5WIKYl1C1+Osj
tMCKmWrI6n2GcK+nH8uPSULrhdppeLA+5Y10WThMKMtgLY2B1lR1JQekPRCP7XlG
v2QUu7CL/b9VALcV6/8lvA/ccYB+ojOQfqG7PHHOBhTmVRJ5swFX3HU5Z45BTCSw
rxZhIheOMgTvdJEaC5YmZDr9IeDbx/OKV9Iqjgkh4WS4W4OEDA9y853prwQnMhCT
TFNMbXOmY23jG/fWdP9umxvMDNlijBdj5VGoGQsf31/0SsAk4QPcFGD/J7LT9/tR
nBgcQy7kiTwA2eS270nDes0qHV7z2CqmT2u7v6S9bsWT8ySpiWZBJV2CFrOAzDp4
CEUR5C55zXsATDCdJVX789Qg2Qb0udOzRMVJ9z/HxQbxzYwY6wBt1Z3qpmjwXbTw
UEQLpvVYcbOSJkKSa+kovBsrP3axKLA/ga0tDnlvaA3ULpDmYEb+HV0jnvhkYjrr
fD0FVolmj2zD/3MMJ3IwdZ6wq8wMBRczP/S6TQjEaIzeE7nWjm/IajFdrLe9KwWK
QSM9ZaIJ90XQUrm/oPXEH/mxah9H3OpW6r/Sk1I9BKqJkn46mKqm5Jbufh/ZSHSG
5Ux+4DP4jxV7yceCe+XNzCc5isv5i74vgdJRiBQoC8ug1MVMmCW6tHI1fzV6wdk7
oGMtsyVQBe5/10Aa+VVzwzuAjGZztma6LrXh04NlCF+llb2Bfe75byFqIxXMoX1I
e3/O3xFrefqRgaJrwXTHsfgL+PRvsISEe/DTIr6k5QeoOSquDi9nEp+xHY9jiMWb
nFJORO1QOkh/XQHXbxvwUp/opKRJLPlZlJknief7LtyRFTqzxZPMH87jDuIayFW4
WjFrwYcSk/Nz9tnN5AwVUoh+o4jQtXg9DG+ANoKiRERi4EovmIVwP55R++NjdlFO
MR9PeRZRm0TbWGe5YU+/Vwd34IIYJkHtWOcWHSUJTZkOUnv0BMKQnHSFRqfFY7ir
DHzF7XssrLmsYIVG0DpuWanh107XvwrYalzQAwSXSv/0XJhIcue09w4GjYdCzhh7
RHpaorCdcYPSocYILc4tDGG8ipy+vu0g9s5XVVEf0Rj8aARqusT60x6Ji0WttTVw
offhWsPD8nHdLo1VSIM4S5kO8BedRl+dlj8iCyEQZ8xuX9g0BiCu/QAU1EUierGd
T89SX1GnrZtvXbEFXi/TgElm/BhG8yMhF9xGQ8Dx9QS8/CAIbWlLeCfLgwixrXX8
TKiUf3k8oeVKpnRJyM5s31kX1gkxLP2zGKYBAhRLhqlSW4lWmJNPT2Jw02I1Mv+a
vmeFZLlpt5FFmjSqACXBr/6Cj039qrNarPtXtiLhNg6mXkDl6rlh1/0l6wo6CAGG
ivy2sc+HcjgnvDgN2El/j0BjpSuxANJCCh6oEqkhYYs6xYnQfS6LMCnT6muKmzhc
bvMqfbUS0ILwg20Qzo7ey6JbSwZrumWMigjQW0o1RFd44VKul4StKYZEeSXj20DV
h6kHaNgvjEbzRwjWFWV/NdC0cNpUcPfxS8RvIjrSAvxFdK89IsIVLCO8AW0hpZxH
nD7mVQBQWHZwXNBcHemAYAXP3WxDyePaqeWkFzGYzmahCIf8Cft0siAgUHvw5Q72
nLLhOhmx7gbjlGXJ99rMaJ3oML5zRMMihDE6UcM3kAryZbSXlNbekYjQ2kGd6PkJ
UoTxZTpKfLBU7fEZ7FZoFg8T+D9UzUlSwA5xPGeDEwTPyrwSx8VRilauLkfgQvKZ
Q5FkBlsrBn82KpWpPVADCJnCk789iGgeNrRDoXxsONlHW7S7BVkGOA10bcKiwx4T
RMcKU6OTNyrGGWZRCihcmuqh1f5nyMth6nsTdWY0wRIOoDl+ow1gRm5po+E45lEv
byheWGKLBPKUGCE1V606X/3BUeo5eEMlIz9hA7TUshwVp34+QVjKjfaFzXXSKFD8
mxAAfD861DGQxQRDplegvFiARM1ouy/Y7WaLG6ggZm0ToamtpY25VTGRuXZfz8uO
Rs6FnqRYrG/mz1Yuft5Xd6HmsP9yIrWXEbk9paX+woA/+XwXSb1ofsJXP2UejOBt
JNc4Y32Cnf49GU5t+fuTBmuwhis6ocIslvaNJqyguGapb6LFfR0rO4+VkFcck8Ip
dk6TGvpff52vPWUTLEwunaC5yV720/7VHKT3J/1/PoqJpL1+JW88HAiKRwlhZmb0
1aedXFOzjtlS9qhiVIY9w/4Cao9h8NZbw4kF9cqfnHbl59WxtvfNXq5lD12gRD2w
em7F5IVyJCBJLmx5SbZhkcdiMX2iOOUQLvv/o+Ia2nf9GdghaoZepvcxQINkxIZs
RmmCMhkutSj6rl3silZiVVdw5fzHrbKF50AddXxtUB62DBOmTGYn/pYPT9a9Zjc6
tQsYQFN+zvbnY9mw/V+0FmvknR9qv5kycjfbzXHZ0HOoRlGcDuvOhHezEQmWHMZU
Xd2sidNd1hnoi9qieXi+/mRFVlO1WAnIM1LE4EssNMw7uBA6CNOUBxQZFWR7hOL/
idFO5JDw575q4CEwDgX0QPvZLGYf6ZhEI9/wkneY4rT+GR2L/De8KqShVutPNU1i
0XqyzUIUcsnVOAt5sI3wj4jSIdhurR7f32p+b/eRn6AJZhJ/jXW5rXFLuEp4ELyy
UW4HUU8e74GN87A+TKIUGM9FCNabC3Dvd1EL85qcghZG3rx+qLUN31VMIs0UnikF
f4/UP+rhLDre6hsTXp7Sc5HQImBovk2Vq8nsqEyAPSwmJKZ7bgSAbuaNA+P7AvQ5
YToGwnW7ht4zkEvDF0i0e9ufoXU33vwRqtfeaIhk30VEA46cCdWrxgu9++cq4Ppk
awjookSEElVV/xiW4LaVhj6ijQffNpYD4T+FztWqC7GRU9PqZ9OTNJnGEaIi6bq+
nhG9M2z1iTJMTnlXNPnLJJZOxHduYzOh4wTDyHPaYrvhq9+kVaIp2OGh91KN+zdm
Y+IJW6Qt/FXHWGYRIJ+ahls+QavmPcOk8xSB3mGFOMQLL9RdSeXcGq2eh/U69qy0
uYTbHLcQXyLeu3crJnMKbIPPVwnoepQS7zsrRb89e7W6LeIvgCwQ0L4gVisqzIF3
FrxqUuaEU3p37xttKRBpCtAYCxzwAB0UTx8wW2NiaeRpeworVh/Jkt2jt7t/KFGM
o9Jw0J00BP2erxJKq9q+U+2At+hbsTWYU4g9707SB3JVsQ03sxIW9DtWEkbWhkcS
dJTSMaQfUm4G035tZi1A7WPwAy2PUdsMCv7IsUygDEA9gD8QPQeQwdQGXPDH4gme
uylEjq+RTdFkLn7sOkTdyz+ouEg8qRLtZvR9yQc46QYVxOP9C3isoKaxvG8Ntbg0
w79aErw//Sic/SMmBn4B+EvP0gOjUwMstOrKPwzPrQ+slVfsMrsAopOIP9Cf7B5d
27i/TxeTe4+i723njyLQN+mIUHwLKb27KAUbP45FCnHHcm5c5yxUnvXf15n9pc54
HVGA5abMZQyLraaPivZ8vLXTF3aWt5eymD7ev5oVulTpHAaUWdLdFHSeGJJVXbFu
2mpGM5+L3wj3JybGlgqN01ma6d1H+xhzC+hCOzyV00FDzANfkjcY1JxtH/aRUrup
QWRx44z/23cSksfPpw7SWpDqFsKFCnE1PBequSFVh9ljM1GSAVMcOQscT3X5D9io
nt6OozFeQWsj2ZwCSWL7c/GnJ36qElTl3qxJNkwBaVZOmZrv/IyoNBDQUCeo058s
jZICBEyx9CNWmgf8Wh7XgscLmfL1K8OuaFuPoYG8JpBHuTAh7T6xIT2qFTOWNyhc
DYjjLgRjqWxIkJPuwT1/T4EEvcBRtkYPhw1+iGXGDIksm8yG9rLWlUtheizyzJr2
yw9OAEVB7TknWJ08EkzKIK5Foe8vI3hyxVB3iPedblQ2+r9Xn/qkSNr7Je/EPfiq
LU4wOIhcb0xZs+ZiM2LzSw4XCXpz0wfZZHLRNXKfoOKJS+fmgC36zYiGoH5257Oq
ume4lDoyujI4R9ODcgjydfqj/xFzKsl8/Q5+cVNq7r9x4xP2p6nB43i6YwQz9eFX
sJA79umsgfdFbDSiseNjd+uydTCKDOlsdLIxeMZghZRI0UxKFDksYLlHubAHeDms
3KxKrTPaMFPqWEgZ714ki4cYtQpvC5MX/RolG3qKGpwPeEIfkBuLrakHIUXd8Qmv
qZMf//zHGPdAeH4nQZQkrUhv/Ss22msnUO4BFGT2tIpOT7olFwdMMbdF+4kvRKPQ
/1wramsZsClcjVwJusb9EaF6kMA23VlfN/aMjYAnDxkUGXczGeESJgGZFKEeoOEB
mnc/WOnls/yIEw3sAfQiSNo5RagCqB1jrRssXqozOPycR+Jc3RqdKuoCDBRtKWQ1
+WzDMkxgFO6L9uBkO0a3BIC2Ikn4cGTOJ4DHSeq0JMt7phjC0lJoLqSEmYGfQOvR
Bn08KbTKvPLcvWmE2W0vQmD0W/lvn1Dk/g+eVMziUhRzgbXC0Lw/XB4SAhHys10N
Sb4YveCq8VfhW9vUbfz7kMcp62B/8x/2rp7mZRgS/gPw89CWeL1HLZv2YCDyWMwM
CdMOM+W/5nl6AKnpIqV2SErYlD/QYRqlQ+U65EGcPJtG/3XaBhow1Dw3afAu1Zas
lILRP1qvrgitMsSpqDA56cBHVoFPPRxsNfufmwKxT3aDcdc+03oGwxaNdPzqPaHB
xjwJarm2VLsHp52ah3tNSB2qkC1RM9z3sBmlbUhN4XSPZhRUfLrdooTs6CoV/t8F
XwbNwekiNm/IKijdZHkjCjdMEU39gRn/4G9R1WwtjaL0QopS2RZOd/yHgCN4ltt4
fAo4lJQCM4FNGhuhUe1pUtCAkfU4bleLkgv40NU8ORZHA6dKvoFfbSTJ6WRjU74w
YHa76bAZoMcyQ/D1b6tZvZq6o5SKiCSP9cPDW9w/hcQxlLeEf/COmRkcgfFQRbKB
Jw2pRZhSOzvF/5YnwWApUxrGI4Izqfo9iWdcqQEb7AF/qcUuO58n7mlI82MKJigu
1FehcaptHBswl0YM1hoctsNg5hxpxVXLv7fWlM3hbjt6x8iBPf4gMwIS81sGbduq
wLm2NNaAJagC8ACiqEgu01Uacm6+GM+6nZ6rMxE7UXgOLKfug0xuIvc4BWRtRvx5
2r/laoTcJXXvfvxGig4vPZPCTDHu4S5ZECPuoQ205RJdOBoG7RMh3uDqGavuqimC
YP335LlppuqjOj00ASxWMHjj4F5tBvSBDOowGIFQEayMdKE0tLjuGL5nCiNlEbtt
cs9pd53/xmR22b1mRYXBryyxMQ6gb680LDedukD1EOP/4lEdZQmN9yOAw3i6nxIE
e1z24dpxjKORmZEpz+IeOaJ9EAkA8gSgPMeqv0pyAVtMrj/KbyRcDW7pme5XpiuY
gVQL6IK4wIuCi13t1moWYONC0znpt6ygOdK+tXDRzLFwgAv2oylQXFFD4x8d+aEf
jo/Siy0+1p4WSpSxrqoGhm+xERRcFkbVXHZ5zzuB9ThvOXS/7fxxtYxCdQ+KiBgT
eNsBKGXyl+x7qzZTKozA4VfM3l8oOxVjKJ8mSM05DxnNzsm8iSIX6ayhVv98v4y6
UxKpBjBQeiC4u+tPjEdW6XqP9HcIfKD3nuKFCuQXe0U2aspa5vx6b5z3IB7rauQ+
YekPw5ezYNGrMl0+B3BpnyjT09FbPKBDQU8KgPw1BSGiabq7LzudAKvcMQViRbO9
ymC1XS2JiFCyEbVhdF3exgvOJMH+YsLLfh4k3nNfbUwUbRlIKH/APUz580StkOLk
SOj6QmwlenkDu3z0zfKBycX0MIMUemzgJjSywfR9rxojVNDMkPQSZVfkcgmHLyCM
j/pKSK2ykn+587bxjkxOesHxb4PYfEYw+ODdLujqAcgMUBqZ772L+n5LEGG+pP9F
N7wDAZTqXuD1ADme0DwKsfDV3lLrJWBHoxzSptJH4JRLAiojZPkF7hcLaoPiAn5R
scINwkIHnmqiL/Ii23MNr+QEsY8N/draqKY0diw64O3640ERfbsAKj7FlokTBj5y
ww1VDR0+AIU4X44jxJgU5yOSW6QFlXnAq5AT964v9ffxYQuwko4zd6Oo3+X3jZ/n
4b3AmnNq77o3SAIRakaw5DoT6C4VNOsXr+fM2x0g6a6wifuktJ7nv+JE5/FYtrS3
2PvMV6zJZpvhoIxwDXs3sa8ZCP261QINm9sdDzDyxHVwdNTfx3anIquFs8YB7krS
GCZI2HP398ZwiafZfN+DJ/AdnJL+yEj2DiKGPwnWOn9jV+NNnkra/kWjtM+rSB3E
k5axyhog6UXEoJ13uAusixgccxLJl9Tr3w2DeTl78mihFd7h0HN3ti3BMk/F2WHL
dt/JkEsr0SUsePP9lYouySrUpOqxGlCq3xB/xQoVH3QWoFdKHZrL/LIoCmDSCdJa
fUVj4KwhqO0dFA2lUzjkseP0M67AsFQCY/EYvxf3SCbbZ3KnsB5ZVbvKK3mcH80x
psfjjYsvv02laWwjJQra30RCdGcCj/rSnKAOnlBKdVYuCVnNoqRI+ePxxG3jTged
fqaiVJxk/NsFQa1FIJe6EVFRhkA8NAxZVYII0XB/86reuMKdUg6bJ4CC2UeNAJZ0
zsSzYlxa6zmRdNxtMia7iE1KM/S2TOVikBUgtxkygUWWJ6Gy0nE2R3XX/OBMjhyC
B0vgb+3KFo9f8BwDXUQpJpLT21z6uzi0BeUddmiCYrBFOAqf11uOh/ny4Bmm1OLN
15SQzKCivHE8bwLLTPoYGOTDxDU1fziDdbfNd7KEYUnQNnnp1cCYbRlTXmz5jYhz
LpcLCO5fdpc+lEjW/X3m6/M9y5zVUTHoc4AoCkT8W8DksHwYl+QlpVe/aOaNtzuc
nm1O4XxzMfcqhP+QWGfPKTVHfCpyYPJoqjqASyC7mZl8ZCaD3sxn9LnbrH3kKuPs
RE02rQLpkRRKO7ze+Q/ueoIIkKPk1EyfDN8PUse9rIJa00fgMzG6YouYPxQorc6h
/8M1qYCYpMZpI3amI8c3Vb5XSMhbNzEKWo/Q3tWfg32fqR8HgQFybnsIpP5KYtNr
fXxZf+8GpMX0h5f5igtd3sJKcmEHKeCcTQ8Ni100N5FNv+lLPLgvZc9MYEUNN6qq
uWnLwQbBDn8Tz6wsw2Jej6o0EoGTW4EDqwPIIv+zXvU1CtuFVHF+Gmq/m0g+Cegn
OzdFYQX/wA9p73y0aBeADYJxb6ek5la6lCaLkyYCr+WEAOeMdEhsR8/Bvxk9mejB
0nYdsq6ciCMstk5PjBaPycblIqavZsbSDYJ1JJCqIqc6DmU5PHmamJvAl99GmDYI
njycELHwCSRSg2JfqVPnmEfxevyUPjhKuPi6ACeuwC/qm7tqW+vDvOJASamo9nmn
8/51Gf5ZqSk8TAvuO8dbzFIfE0/wG5QvBvX5Md3T2qnk1iPZV3cd6ZXzA6zRJrjz
vnk6rq7fa9syplp5d2GwEtBLt8cde7D7TBtXyDIon81Hpydh2gN+CiRe80pHRjt9
IchwtLGlqoUCDtw6uusDQuOr08xs2CRjAZYuamgCejIeGAyHBUERE4BzF7k1+JxA
HPrQ0hvujmuoUqwktjc/Ih/gCuXcM2Z59WADUJO0Y5VI4F5NFFdweIDd4pjgIFnE
G1Aelj3avpiCOPyjENPyy2A68U6Of+lZiK2vXQcL/D1gpYMCqkuLiAPQEzgvD65/
s7xnQ++labpQiSnuLbLsvZUFdGUYspR/M64XUVmlloA1ESPkmg6lj10MMFGXdmfW
ou0/0sNry74ZH8A7VmMVy5W+rrnxu6NAFnLAGhRCVWQAe80LWO91h8G0hTrNr0Rt
GbLFxq/YcZxJ29uxslmos8/abbecVcPhZ+TtmU2FCzsJikoX/HY0gKpDy2gH9NMe
kSQRAvSYWijJYIQUhGFJIV5Cs4Snc9EjyKVfKIWh9WiYlS49VSRMBENlX/1wt8jx
4CbUytOuzlBuIfqo9tR9gdGKF1DG13x5BjO4HxkEwToGRdMA/a8QHgSJcot2DgM1
iDFQf2LrTPrwFKMseIlzMGfajFKjxdQ08z1A0xLztcvXQxaV1Fv04FKyE4pjWLoD
+fVYC9EQeRdHVBT+5ftXz2c756rtSBMlz2kKbmMInFSmS0dKy0d+L2hdR9+P6thI
ywwWRBLH2fl7nqxFMiCB6GSlAN38Wfs8q5xXKJaF/Vk2nAwa0lqk5UEwZwb3YUom
c4tH6UhX8S6CJuUXWpJBwTZG9uEGty8+ufnzBb/P1OuoZ2Hi3z+rZ3YZNtEcCwg0
ZArzHMKsBJooWkBIUOsCd2+4FMeCTMRv1FKZZpPNRNh6IEC9jR7mfO2IFelldQAG
k63fvEpA0/JuBKZdBSo88CgkZOnRtJN2UpkGOQdUfQLJncrQK75NpqPSmvrlvlA7
rXxDf5tpp4bii4L+2Rm0JMj+A3fEUtROM84GqU8Az5kJ4b/IoYszWgzwJnSuwN8w
X11+haWu7ApOJBQZq7QWvpPnOcModH5ClacQ1JMBhwqygkg1YUEBoqkgM03FyfOC
nsu1qwc07QQ1gPcrntJbsOT63OGzjArPANd+uVFR42z81uV0yiWwA7x0w8XXCQj7
fiHI4VtWO/sy7HtA4Dmiw7RGPxyoRyoTyqBvM9fVO2b7dpSg6xS+YilekdVmM1M0
tlwJ77dGeyd3/PvG/e2VdjCKLLFBqIqDMDdv/v91dRoGou5Kb/TGtFZ9DfEmai5v
b8fkSRT01nL8Ym9aIdHVcMcFLiMJdSd5g8EHBnbCUW0y23A/GTAnx+yWKNSL5+gI
grf341JoLz67toxV9c/mCaLSntw/TgZhKrCfZrxCpV5f6Fmd7wmSCFLh8+uUYmsb
NUUThswuzsLl/6YNNEDSTYNoE774ONRjt9B0KkHz0cP7NQrAd0TdI2EMmc9/vo2c
wnCS2UsJDrYJKvX1C+O02nXhvmj2EI1DEmN+pGXEeOE/ZG0BbIkgfHX+ApZBWWgx
9xuUR8IsoEMjAQVlm78IGWVViNLV5J4Ewj2q6DX1JgKuX7LP0Ly3QG19lN/vCtr6
+Y0QxlAjR0d6DjJVHj/jmX6oxST6X3SAF9G/RYFIRaIQ7BOTcdXB6HtHNCHhOf6M
yJ1wpDfWxFprpjAo+0lVnAUFxjisoAht3BLMXZFmk32VxRK7xcERnaHz7IBNesgM
O1HHmVXknWtaW3lcyQ0i/fMGG13nx1xxIjbTvBB8JiiDR7AiKWpbJ8SRAAFNLj9E
hiWsOkcCJsGtu083CII6lADI3AtfuDxCmzm6qpiFd+eJh8kDRI5Ndjsj8xpUji5K
vq2Am/QbJWPkOG0xYFhKwiJ6swTXiYItP53nTnCZztZUjvZGEAjK/baoy4aB4eSV
o7kFFIq3lgTCSI1FI4ZwbPMlUdvtMUCk9VUOrflBaabx07ujsSiUFaLQXjU0dWFc
b0H/z1ToKzDMhqiXFrpSjLD8OmRShZ3l0CFs7CdPVL+q6DKWctu8LSJ4EYWCCU0D
hisPDEQqt42DQ3FP0dh1qjMTadYC3tXuztY1ul2yCNhupfUPFih8kfDqgPyIAub/
6LbUQjxHSLK9qWYHqEqGBz/aReJceOLhv5xdKpUBKCjBpnP+UO12z+/XsSkGLZEV
KthMp08mMDkTc1zmM5BwPFtqkPVuNv2IqvLlEEvPvOmdJ+4tCcw2W4MhbSdWbNeM
5fvKPUK1aYeYquV0xFHjKMM7gow7Uw+CxHrCh4d6fHnG76Qs0AntTYLMp6qDySW1
vYlH5XTaLl4faIjgTH8u+AonuYQcivJEjsMzAH9s7s3N3QKh7xtPOCUwzEBFDyw6
0NFEX1BNgS8GYMChn1/HS3OxC+3FqMLsUOLmImtyZ4VtfIr9BNpxgTexD/gj8zPC
jywZ5aTkIMAPO8OgU32hVqpXwA2qFORw76CkxdNMZYaYjHMCLqnqJv4BrKrJlyGu
kH2QeOUNsBAALASfJci4wEvEO7YeMaV5JrkQw2u9wslMGVk22dUXlenCT6E4aH03
MfWLgn9UvZamuSftcsYHPvWTP/Ddujzfe7JP+2xZFmRj7PxBSrAdU0X5gio/qz9M
nF8bEq3lHEjhBHKnjbE0k6nN3/M6jJYjKRio7fa29l7YwbUhapxenW8A2s6UbMos
7A3TO/RDjS3naiIM8ETqdooS8wGjNEhdJRdcSuK5RODCtHOV/BtEhFz+Qv3JiWRg
IaQx7+2DgBMI7ftD778b4hnQZ2aClJsdLQeGU/v5VOVvP8S5K0Uenj5s3B06Qwxw
jHVTtOluT0gveO+sSxXtu6NwU/2qKxONKy4aoZpZcy/BhtB7QNMYr37mEw4aYtCG
SCrmCrNT9avN+lP9rCp51wFzu2beLh16Hzk2iX2NJK3hFELd5RZi7b6kRq+ObeSn
JPJLqP9ZBeyIQmO5aMFhbR+8RAHU5yv/DZbe3qxKfVpnw4jeLVhfBpbzMa85+fTP
HyeJbHDviMSu9JcQKdPdLkvRdMb3XRebS94IwtocH/YCNIvPkwscO4PQ0HiiUK1N
XZA5fvtynYkJX5OPkGSOjv7J4DrdBSAv5Q0ghcK/DRZaXYU9tBgOt1SO3RftdxYW
4uD76pm7Y92kYDmw1L2uvB/SHfkY7VyW10cxvxaf3Ow5UCix5ntG5pgmm2r9c9Yb
p5Z76PKgZ0bLNJnkwUDcFzhhSklsRlzgKAdpUBatirCrDAhtInOSWfcK5PouMOAV
7FK5sA6MJDzJeyUXFkF8oQcc3riSuHUzOS+g27VNXlFmf1AUt5UhzKr6Za/7WTgl
uKftFIL2sEloqSIJqLch696T5Nrb+Rr18R4aQZhuTaNX5fHuqx0Ks8OKyu94X9b3
jbCZbrtyb0KnW6PDUoKwffEqwqnkC6Yp0drfIi30WXCuWB/sL8cJpwVH69mOkR64
SBKJSbUZRKU80mQjTJwq4ScoGDsEnyMPAStwEbCsNFNjXyNEjjNMA3AgZWVSSZ9I
V4mbzvDK0Kp42iP5kirD8S/mJaYthQxs+4fzOBFIEim3ka/OzSj0zjtX7dD6ef6W
JIqO1JFrjMmdjZhzgp2rq93bgN92nxfRia9nC9ZeBiW1GBC+kMw7VevIjyTJzmc/
ANnewi4bHyJZqyNeHut7IAUlHYTUIn9hP1YIRZjQva8avVWG6liakpTc9OzTvS3z
acwtlvcxz+v7WB5asZ/r9BxOvNkejA80oDIqbRIWaswkXY/ydS/uRw+On8X7gqoQ
0TZ5kaxUxp9PXPWps9Cgiv0Ko21AHUtZ5MD1ZpYoTnkAB74gL5nsS6uI3oz5thji
azMvCxg2ZGkTpg3a4ZdSd4tMqsrHle7iv2G2qirfKDwP/vTLxHKmkxTsvbeaxY/T
eUDG3y7oUin0ALHe4c2WoYhW4cf9zz5Vu5AqVUvCeRXhDqYuX2eoIYWi6BKloGR+
NxvxLbfy0TsQqkUkSKlBqj0U3KI/ZN2V8sKLDQfT8FqGGbfaScJCG1PRHlm2jiNl
5qaFHU7OlnnjrMli6XMcxtSJ4uzBVF4bptJKsIp3ZVOzMqKcswdF2t7vIC5M4kHN
mv+vDNY/fC8anbvKmhmEl3xrl7aT3iIftDfzzmgStV2e/xaHj1fBRxnxkbw33MdP
OkW6sCBc01x5IBl30/FAsNsJezQ59nv4N2kuigboo5b0HEWA/2klb1TaXMZQHKmf
1VdVT1OYqE6ThX1NNltdMWReZfvQkW2L3NqDtP1x4uvuGvr6uUDcFMaxGYlUiZ3s
V0NLsWq+5AzTZ0Ed3ittkxMFC2zvvRM9v05Cn/9SpB/f+ZLtPILSTtWSAkndsbtK
uUweqSh5yR5FSpPs4tA6C9CFuIF8Fpt/xRis+auab0MC+Ul4lgeMVkDnyg/jBhCm
R+O2PCdRnN7cXIutDT1bKZKFT/k4k2X4yzD0qIKPlrnN8DlHt7/i1fCHlu7Fnxa3
oDGo3koGgySdYX/UAaASnv6RQaSHDMIV0FhjIdqzB+y8EsE2cpdAxOm+ukl2I1St
fSRV/tpAH54TDDcLZptEujw6ObYZpU8rJUO2rzskcLQnAE7htsnL5RYKmJOUyEud
Zhrarc4+WxIQNBXCoY2/YUZYCe4yes/R0fW5QcEVh5b1LW6QlzHrXoQ/9ASgBmY4
kB0DHbvXlTRY8BOKRWkatb1UHdT9YzjwZG4My2Bv4FIahuJWweKzX6rGaULJnZEl
txry8vo81xJLoIAvdDgY+hYxPsGM166ZHsdNifcVRxXWCeaXqzcFEBiZh+Fg+6NK
2N6+T1V5fBgG/MVNIffGAFKTBiDmyaFRU0t4cmf7Am7DpNB6ifvqvOvEqV4cinnv
aancY5saI8MgQOcxRnuiThdl1qfuvSj8YtKdwgy3h2ceQ70TEE0ufguxzoVxu29+
+YktCAImsgT1vzbazZqwMYAj5dl5vGU4xB9BHlrf5B2WMYGODkl3U0kQMabQ8LUX
MFQYXU53Jc3VNJrM222rPjsEnDC6yahCIphLVWmB6pAwtp34K8vZ6Yrq3ryFJoL4
0E9mDAQM69202B9zh1MWfnIAkeP/+GOi/b+LSj2OHBnwkEo5lSaRdWR4JvzJB6ow
DpzllEiug8aBkziS7rQpMEYhoAPiwY61/QlhkmJxk+97vEzobZIe2ocr+3HNH9k4
DfcokebtIty/vWaWzy3eFBnrhZ2MU6/Z1tLuOWuYmwdSUtLJM52Mo+fNnKDXF6Z2
yx0ybQAMRhjCDXmjIXDdtHGDWoOB8tjDudbTU+gNugVlrPuk5et2xU4orQ4BpYQP
KvcUUbD+xJcMuBthcmXrRqfeSprwCUHXm6r9Vu6akax2pMS5bAV2vH83+PuYpgd5
qIVlyuasSX+m87tC/AqGWBuw1MacrutkvwlLi+lGXRRhUFVBbZFAQ6Bgn3FJ+EcR
2fCj/ojx/yqULqZOC74sy7I1sU1RKXTzfFl1gWjoR7I5CoaEV/SPJlIlA2/eKejp
BIhzw7AR9E7PPkUnwiY2qrWBn/avXh4h/LvYZx+mjTHPGT5+UsIFjybowgQqjt0Q
BpVJHnkwys/sWBgyCoUtZAxR3IkUiHKvfogATgOC7xlJz+0pTPjNYTWZpjQVFQRt
yCaG85IkW5hhPJvC7LtpmkH27zQQ2Ek3+Z1ijbuZhPNgtlZjzyvRieay5fONRZQ3
dHbj9I0UaJeopobQ+yldkZe3bP05W6EGXn45Ent6kQ0JYWkTsSQmwDP2UgWac+mt
JckZtvSj0k+d6JqmHmhSEdTpGv8JUWOy3nqSVPzsVwP1VT/da5TqgR6F/+390fzA
Hfv8eM7OfOgx17HGO1vbn2Fh1NUeUnTTuWlSMamQvwmsAsAc+2qSQFPKwuxDu2YA
t9g0Peb7L3xbma9iQkJ3J5DFmdVV8vl4zF2E9+2QsiS9XxoZxX0HM8BOYkgBvIFa
sdN1R/hCFjSXIHEDsAOVJpKlog8t6L4nBOioajYSnhMLuXr4QMuMDlN1ZCzzfdM/
vuWa2/wRIYA/+r23Jfo/440EtSYlbiP7MC8D2OITQ6o4QgQ8Qdw6RZfzPqSvotGL
VaCVI7eZocteJRjfsrQ6O0mN4KB7XQ+M6h68j+t973oYb/zZ8JFgsRaVWixx9x1v
SgCbW2g24+b/M7HpcklJ5/3XImh1B7BW5IcosLj7c4PMnvF5HF+dShUb7+HpLsPD
bUsiqud6fYiAxf6lxm66aie1QlfDUchxtjIcL+1mdoqd8loLi683JtAMeDx7RLJ5
mIPjTyUXjK4KVThSCFzrXuoDXEeRYdnHBrzaKBAu8czdslrDxrK2XvFKqEswKKUf
cBgItTdFZjqYHq/aw59aW85TCdBaTvYADBA2hVaKoBlVczwWaI8NPG1TbPNh3kOD
ALp8x8FF0usJZrIybtU6TE/QZB9s/u5n9crqEg6F80n/dA9ospIrKuF9o4BFfYTA
WJcielJW16jaajbcTXatKA8mWz30Uwf4G3bmEtW7hO1xmHj2i3F8tu359nEgcjbV
0llko7F2N67tLBldbr7A2lYvhO2hLfQci+kiL/+IBeFb9NhrcSOKs62OPkwG2eYU
dTknmvpYDt3vHKcK9nI0tYzxEmzc2aNyFp65LQWrAU2bhQwjrIUnwj0jvMP6JOlH
o2vhvjgHS/RpkIEWQ6bUbW4Gw3Km402vJoNQjDYC38K7e70fgdghCZk4x0LGEQn6
aefgOyj5pAaWzInWwn5tqpWUmCu7f7SRLQ7EHPpL0jxibhbOGftBFuY+KXTvL0OY
EMeVTpH0byojgwu1YrSvFNGnckFFx6Y4KralOta89uFt3i5JQa/e3gSm7RNNaxYG
UatnE/NLawL/+pvey6sRSPbLnd6wOxxLakcWyyeA16mFLxvT70Yx7Eb6UOvHgLJX
uKGqh9Bp8CoulbuBZFDmpPAb4Zu9U34/1JBYyShuI5yehm/+wI0p0VnaQPuknJVA
XPdQoRdKOTmARUwF1pifOCkQFOOjhK1IC0LsgWATj5reahUbBLoq94/WNiAIk2HD
pA1/oraZfavCXZ8V2PUY3MvekVoReeKcIE9czQAsWyfC0QaxkLjOtiBLj1oGnPFB
S0u3VLJSYR4qYze9xMqXP0Lkg4uJ8jfsQ6DF33aj0lB43/vAPJGx1Rx+qEiEYIWJ
+55LQSGTsg9MdiptAO+MhGv2fiyy9QDPpT3VbvkhZ7yrZWOky8pk+YNciABTrOEO
k8DS07gyRJ3wlLAhpNiIXqW1i2IsdtsSy/cp+QXZkoGtpqFC2jrXHM+HnKnqOr1F
6cE3/YHV39JulO08tH2NVbvtwW//q53T7KL/0Is/zWoqzF5LJVsfYKnOogG0x2SC
SWAzWxvUknJMbngpOZ0ZHaK8qqgAaVKG338nVDnmyx1Y4Z7ZNMI3bVo/8EXZu3w6
8IIdwF/NmAri9OrMDWduHjxF7zaPLhy0+yqH7Pw31oyqMuFKA9qwrX9LEj0Mup++
y2EDjTCpl1pJabiMCBz97oaSL/1NlxqmLwsrSEFfuuJIewjLp7tdhFbMywd3g1ZH
S/p8swoBZDWBjG7RaYVYrH2USmE6dPFAsLTyGvNGiZXaRSoBClVD2z9sn7g22XWR
eRBuS6ne+OXBgtedubbG7h3hYHE17azfLihCY1QXx0h49waNWGkGVk2qeKz7uMYz
nfvq7p8qNTqLuXScKJgs0EYiFU/8RgtelzmOo1GDq6sPzIxQ1HsS4w72MDSvr0dS
VBJQ0YttGKiCXVGFGRnOr0w+GMmxQaFWa06O9y/94PE=
`protect END_PROTECTED
