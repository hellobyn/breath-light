`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5yYYp+a1lgQhJfxP4s6py1LjGghGByIw9ELAFka2BJ2Yywz/CvMzPgg7X2fRKPc
SlpD6slIcEpSEEiH3nbftE+QzX7zHRhfd+NEzopbOxfuZZvU99+QsjlDm84r/9Yd
7N/yPmLzaOijWFCDVxnjAz5LFYbI7/2zruSWwNt2AiO7BLlmnygsbFkwhp3R4jmz
7P6cAJk+joBxJuU2RQgjWEy/Et0Dqv8SC56CU7eZgwgeKPCucNqsr7AMKhJCdTjq
A6NFUNodMjYej5N5eTM5PV1rgJ6OQfIyCIAXOyGfLUr0STOFwqmgfCdXIlR73mil
VG+cChdPQJejjP1SfdRNdjasPCet8crlbMteX/WrQhuN6Kc5Jjo6PThEkjA0l76Y
QXRNVflmyabFyRRS0oSIAJMJhu9FWELmjevPVK2jw9nlOHbVWeLLRTTGslaAS1PF
yHBeVi4vEiIkeoHqRSFw9eHWRs09AjevGHaDi0EqpDJQTDQNgQgBe6fcWO9e6Xuj
rdjzTBXnk5uXF/JDuw6wSIOVJBMcV2WUiuw8s7eGL/m32Jz4USZSe+qaky2iVxHr
AcMS3DSjDN/czk2f4VWBpEnSevK5pXJZmA9FfW4DRpTGSF0CZQBZTT+F/CzX56kU
R6+AMIkKZWA++z+j1+39OxWO4j4AseDbfnyARrQI/lY6DZRhFHDdGGdlVT7BFC1M
bnMifgpZJaHfG4vrY09qNrMdnSJ+maGd9YYltAyx3LkpgaBaZIk06852FRASiMa8
FNa8taGioJuX/TAmTjSFOEElCnsyRon+u2huQ4X/W4UU8kC9wxbf0D2TgoCxj437
dNtcVtPppHB/mrN3PuamKK3pTan+CFWHZNJ5wntdIAQDE24R8y8b8mh7zbjDqqGx
tDs3M0JHjWY+pvE0C1BBeu7JNz5W2L3azEFSaR2i2spiUpOwMw1g6uVKUtxZbjbf
83dz56jjuZfcrRlhI8fCVVw/v43T9S6RYE3rPVA3p3gAlwzMM/9vfjDJ/I4WnG7F
OSCC/axXSwMTLSpONRvhdrWa+vntNlGoSEPRoxYUKp50Ga0vT4XEWAR9DLUsbyfe
96+azvKnGboWhoN3GrQB/Igl+gu7/79fjVOP/xYsfuFQJiAcm1ApBqcaEN9txJJp
rvE2lEs3GEIVdfeo0T/AMO/2no5ZyxL2378mKDBZVnCpBcGsnsy5RheENYGDFLU4
Rkuo4usmFBs0ZUYnzE0o9C9Dvq0ZlugD8nvmdZjEBieAWmobNsA+IyEwDKdWpWpj
ybN+VsqDJbL+PXS7nQjet/V6tg2/sQx0LZt5aQX/JPz4Z7fBTj75Ul0M+NdQtQ2E
BnLqI5JXMcTQ5vF/wsy0xCLj+QYCxKbGy/S5Nyj40EW06DRbCXUjhzOAUYXgpsqe
JfYeW0YtTQtZqLDJ2ZgcFEa9sdT5DTJOLbAhdPB5pLr0yLp28/VFNcTDHWpzRmGj
Cgw4MH3mnPmKTmmaKLEdkzIPiQueQ5nWvK+W1tmHBL7MZZklxEoxcGrwhxiG4PuI
Bt+W0ipiXvH3AwMzFQObyKOcTes9EnNGnFTbSWkmnc6BWUoq1BH5cqCShIlq3rT/
kE2kewCeLb3WRXGa0Y+MgJAObBzgw2L0FGvWO9hJ1/mDLD6PbJfnwo6VsKYqCeUA
tqCmGMuGalxK1m8aOA2uJgGtT77/gMgkhOLjz+SRVzo=
`protect END_PROTECTED
