`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6h+BGiUzWItjYQRpF2ULsBUAciSQ1IPx8ZMP8w2dgEpdU6e7VR28t0O6ivDh66H9
mLeW1btc583BdhtfbnXKpmdp3m6eamrG/KNl/uEC3rvLCWRVvSxmGEnBfiJo6z7h
sKxgtG7Oli/JNNwFHqKzErLjk9cxWu38fk/KuoUzYboXN7ZlCuxdC2Hsr6FmRSrq
RHY0l3EQ5dWDkpbjwTCdzmyDulFESescM1OmwrgScLDY4+JUpEXv9OZvbd91kp55
38qR9GnEqTGavbnNin5Djz+VxoWSnzvSyr+L19kJwKqisNjjFVqJV6DJb/fNwETm
SfYvOO+N5Z7Q2CoTJ562UtEF030h4si7b0XRwGAFLr6ERmKdSbx6wTG7pHw5nHWk
OE55eQHjpdvxf9fr5D6lEYlDxtAI+/kk7xJbO/aZ22G97gndnyE9EOOEosjo2BhQ
ujFXs2hQqs3EbNgPxEk38OOZoaCcSaCQ8bJU1Y6TKod4RJj2VkX1vkETDsdMBu5U
+aPPbbIsiqScPMf2fXXYnYkg69LAPAfuJGZaZTTPS76F74NZLJHwdqEJ82jj29nG
IBUe4cK2BNI2A7bxMoCTEwsbcufXEikrWEoDuJWvIzRz/COXqpFdyXXTdC9kLI3t
O8KAk4RpNqPBPjoLJt+rWePPHHRzE+DM7HeQPehItGGJjx9ye5OZGFUb975anahz
Lx+gATTGcGyqYjZyslozaX3za5FP0fY0xAxKQ+AF1b/cCVTNY8C7eWlffHEUY+lr
lwnH7RZD0hZgIQfWczQdsOqHqPawgg1BP2frN4l0wXp55EVI007Wqpq+dHzvGqy0
NlATlCpPYeg9Kj+Bn6Vqjo5Np942UDzvNa55VpXrwXSTTtX6JgIHDCcBqhzjTOEc
HL2JIEt7u7rW47D9YoQe+BVlaYqBKtEn7Y9eM1SzPafFHjpkC687kHXHykJVR4af
o/CftrzwdwCIQeCHdHjZvcBSf0HXWZx8zuxVrsD7gNOl9+ut9YTcAOKtudB3eO7T
vcQaDKffWMhdYbm7wMOiKwwvpQXx+W3vBvY4vo4NIl5JekyIooypSJpd+gSTWNty
uIg45gIt5v2w5XqqFBKhGwC7Aj3JCAUdGGGSKpm+ChV5+eYbSaiDONCgue43ZAwT
IsIM4vca8eM5+Q2dVQx0ZYkITPWByJTiT3SUhQz7I3Z/rIxalOiMLG/uMfJMDWYs
VakVGtfRP1p9VztWYi6dR/rK86SxB9hqIc7kdHa47UbwBk3ELISUy4N5k/j1uAFg
4zCQrf7QX/Gwnukd9R36Sxxc73u/mEVzA6MrlDBaKdAZzSDE1GpAIFCCmqTxZtw6
NtC5vzLQSf6AvVt0+/4rqjJ4knyQIvLGUP6kOtaQdFh01dccWEBzoo4ri/iFyWWy
b8SZXb7Z/M5ua1Sga3UPZZuyRuQ1CVwufoMC7k79XWGeRtPVS+zLiLSeSUjxKzPz
5PLpkwf9Bvbp9Q4kTeXBtmxcDZS7Is1a7i2avTRDBXM7hPkauUDQ2Kkt1ldMzImt
K8YG1Y4acFfNsrNurmE9+sWzQDmaetKF9wFSbxTSopCVMp8qVe10Cy1tO8GIpcyA
k5hBgn6I10ytL3urAfXKXJSMJtwmcIMkVp9RieUREDoq/hXC9WJ1lD7GwjvYSNRc
iQ9Vs4tG3ENwOJ3HVl7/a1zlHKc0y55EbslzEi9K1Fj2XyWudoZMOBcw2fZWL1go
WjAvb/3OOyXI+468t6svM6/ZPed8kj0GV/huogEK1OZCcYm7ondSkRGu8SaU35WZ
3dRwfZV96RGtKtZ7UgR8xAiB2NYlVBPLA+42xF7znC2eoPR1Y9RZuTznhdXBjcE9
H9ATeqt/NDYdm/NDYNJ5/i5+JLVJqQIy0CTtS0hpi4vW8C7sFzWNeVYC3pLHpWbJ
XJIXWc16WtRA0CZRGJYkfsB8fQzaFjtp87Z8GqJR3Uq18L2pRIkpYQ9o1QFjR4OF
MsWXvl35lKqhbahepd9eKeKh7xCOnZw7Yu4abXZqYJD7F+jmVwT0YPAPPg0RuPi8
6LGWteALL2CalCi7HEP8fJCaQNegr5XL8+aHQmyNMEMQYHm4VEBzmCKUszJ8j4Nc
ky0TYgC34LKd2VhzGrOI4NMFgRf/QNF1Eu2aug0wsIUvpqwkQwFJfFS1honPjUUf
Ne4YnVtWkAtmS6Q4fpop7zzUN6X8tt1WOHO5JCMHoLQubszv9HfkYzmfWSVWOPeZ
L5/JHJOpY/6WXDysrfbkDZNq7rygNe2+ERAvOj6tae5Ael0Jv+qPG/tKqGOqFXcE
IVh1+HxTip6+M65wWxqSaNWUPkPaq0PqCqNKVWdmYNPIcGyEKjxj69HJGO9In7xO
rD0BvyQEfV+pM+1+KruOk6llVHk/tpJr8+oiHVrG1k/c2qX5XFy/VS69K3lkUfvP
t+QMzjpfkW3lGTs4dZciUgwFwExNeSYJw26k/1Om4os5B17BNKZK1xBOg0CrIQV8
bBeRLe3G+BlXAHM846Gh47hYAourZAoPO2VGDHthZZQkXZURlds/A1GElKaf88ZX
I3uen8xlWuCf4V4qH699fW9uBrRaW1Fd5syBncemGkdqxzw9MoHiAscrD1dwvDAt
iAqSMJlYqXIRVQ2OrBw01/UsAvtvM1YX+a5KDdjSsNQedlcGLWWPtziWyonACSu/
y5HH8VVvsE+/ZXhM5K4cLZUrJS8z6djVAKEsPfCpAsZOtA7tpyOkosatjAXhWFO1
8J7F/zZ6gEhDKTlakoPwxkPgNdk2oBkBelU3gkdtL1lib7/clTAm/vqRf9r0uG2K
VOPeNjdyfIa4xvvQKl9l0WRtUNoLR1QRjWzwhu1kSH6LlSHwxI9p6j4RqQ89Si4C
HbytgOUsTQC95UljC17JIwhDo5Mb0HmjfsK06RE+kreuXWuo1HKDajdjeCzWW3h8
xDbOAvKETe2aV4/g6N4KWZwqcBQsalCS7DGAy+ZyhXb5FTF8o8UWQx7Ikxa2Mluw
cof7ZAEyWYkyUF1eX17iKoV2aen0T/z8OzOuqYPqA3mSHVXM1feD2BM9zEo7oTct
NQR9aNnPHLKQY4lzUogP1y/amozbhoMYP6jMn1WxEhHMsc4LYo1ew5F2xlftgpUX
3ZV3UZpYsvpcgaW2rrFOTHiH3QN+G8Sjh3vbysf2hz6FZINRe04xq/ZeAaZv6Doy
ZCquQ+UR2KcWG+wCPGm6Oa9xrNJoc7dR0Ux+mp50velJrz1GBbjaFeoJBqIXG54t
JDK9hJonpMiWOzpIIkF6UdmsvlZ3R0Sj8pgX0hcj3Ds0DozvcD3RvjfK/7Zg0W6K
yrDRDJvAWKj24+Ne50LlrlCcHf5muBEAEzEmtrJppvWuBdAV0K7duQWV7s3Lk7C3
VLLF1QThVDo6PD4DyUm38Un7jqMmX4fnqt+7E8J1t09uEehPAvymH0vB/e9sZwu9
VKJwRLWjM4GhpO0wXYXjSpXZbds+ruGkik0qZPd7eohtTnalDbD9/zOXa+5bbC6x
BIslqvyma5ByPGLdk6A997Sr8BQiE2VenNBimi2nGM02Xd03c+liGT9XULj7qIfQ
ZcMP9GPSUN3IDsqGnmWzXgEGS8TI42UePg9x0xG38k49Xb++CfxlQDn3yNrEpsUK
GL1MbvFpQicNNqu9C5WVi/ru/gN7wIy31E7ZID+OjDyM+sotuDmq2sGr+Cu6SoQd
C3KgOfPY4gKegw54O5w2EZg/kOhj1eREIneRUDOCeRU4ZfYSqVienTAyn0o0hi1K
bjDql7jNjEXzFYRZmOmY0EvMU4powckYbOhW9mWTLzvtVmLV+8wBWxWGYzgJgDws
Eh+7ZwyRnyNPSLHT76ikc3OL2bJo7iGXMbd5OPXchLoZ8IzSpSf0mK3/bAaSdI5I
OJ4yLmV7b9DV7YL1B3Dy7dxx1rYJ2E8PGDD/DrJP7YgUCGAMtbukyBFhjbMDW3rl
zSMUvQfAUY/Iw51qet4kJ1eg+5iwFDztb2+4mhGOAmHQmEBcx74BmCKsB1Qx1iWG
INQId3KVVV5PUvzqjOgW/rXSEv3J1xYBZBfgRdk/qGVJWQlb58ahfdLzwoYLRNVO
ZDs1RLBB5AAzKZoXR/Mhkc1CuDSomMoY3AQWKRmCg/RdBlrfmceuYJOeqy0TF6gC
BlwEeUcngy7YSVrlsyLfvgjPKlD9JcSHY6X2gDqpLUMt1BbMUTZ3mL2Jq5DAETka
BKzS2Dlc0UBNAE+tKBUPH3jvrhMg6tUeoiozv4xNi1qA8UOYTWR99roU71poesPZ
smaQHhT7olhsmyPP+zXdSE8Vzm8+LyBomFb/UELPtjOXmTuRyL1Q4Ycc+GVIJRVr
zGpAwCAmbJ7akXvmB+bQo6IUP21IwPwaBOudAKHhNBbAc0nhgeVS5J+b+hmWl85Z
B1sMISD1S2xlwlD5hCh05FtC7Kfs/7/Auq3WTzSiOtL+zO8lKsO37K3/jHMeRBe6
ImWv24x7aon5hsTct6Ffe86OuPGaJClKYWZT3wml4QGakXGU0dGm4gVbI+eUhP8R
56ciEV3pgrxznFoBpI6lyPt+1i6FhbsGYl5m6sCceO3Qe4VU89sGu/Uk3kWIm+4R
eR51VtBjptkLhu2MZW7gq/rphLAuRAXE0ou+kyu6Yx/fkOl+9vBSpwcrDKUgg520
rZoc3TqFN/48oO7WU71r02QHeo60ok6VG6UMNhWw+7dhcZ6BtbVYGOHlG+9lsU/h
ZyShe+f4gUoYDvaAY235z9HLcIy5ON7DGjAkHegHokAsAiAKue9oaXRzhMh1TzLo
PsV6YmhtCe0cHFtKXhrCPe59fiLPtYiauYdLvo5jAw+1Hb01zK0sSXh0dvja0WQa
7Tz/7UKhbinSrodIeAlCRLdJs6BUtBViWIizlNekXcsf+6wJN8JcqTPRMqOXq3am
f0EALxRpaFHvY3CsRVvnL2nPLZGWhAmvRGxT6tryft42hiegRZHA3xDgUW1oarAj
Ba7QH7qHYu6vLraVe4SgfV/9OiD7i2QHT0Qo9FaCnLmMis3SfPLfnf3CbfbYxw8F
+6OKvCKpuB7zkoZw13jrslPvA5ygc1+BpWf3jwWRUs7sbSBGqX4tu78Q08raE7iP
5o4n5r0nUwsbJj9+8zTeT+CSdgryV/pvaxIWXBizy2O4OMVHUpH2zhSe7ddlItEo
6l1rr87n+2E6+ERs22M/KpZ+PJR6JBrXPx1bI6WgSS8uDMmjU+z9KP4+iQy27JYV
tEjNcrLBJf/8Nmgs8MUPLe132h3R90LWEFLdhedNUKxGCjPJUOFu6lcHEWMP0R05
8uDSVX+h3KdFoR3Yi9uwH+mNtWbDHctCUCUK81FZFEjQhGMr/BKHpJVXhwumUDFy
Pznjqu5LBJwMvL44qQiC4+xpRv03WTKdH0eZZHF2YmVKOVuT89KzPDyc2cCjZaUP
uZKFSNARYyQX6KFqYjLeyJFgCXmBQecDV/kV16RXt5mKSR65x8OJXACM8773tviT
S1Cbaw/a2vl3u8Suk0xLNe61yJ6MQ2U42imoOnDEunhfIvYkavcwHvvYKFqpVx0P
VbczCnaU7jEHHL0CbH7PFo/BCbV8upmryhfpHmfQUz7Sr4+ZUf+ogD5m+fWpxfr0
QUaLRf3HvvxHGHSLxwxtXIrEb5407xOvCDwESnoK+a7E5DyYNgzNX1TLfXkvlkjJ
vmGyP2uV2+rBZBVxo7a+I4YHqdcl8DaBswrRfhbs4d9Jxo5oWzPf6yrrhNqURbmN
l0JJNdKaYolnjRc077ZwjaV01nrvwO1mCnbvqyJH6heF2OLTWRZSysChmFH6s4r3
Udlo54MCs+guPoer/DRK3oCllgdsE41bKoZnR3wbs6C5SaJ9IQSrj1dyI/ixrrw8
sab/O1V+6uyGfs69V9ZFiQUvrHdBonPPy5L3IuOY93qiX5fuAYfPLgOoOGaYPStt
EMfq8tz+ypgVwWtEQIXphutsNNDBW9ers16NmZrJCEEgREs+jWoocdPXbDNge0lb
tlRY5FvTwzWOdDlpAyJCONtqkn7KeOhy+cuzWuM9N4tjzGCSSGM8U/W1BZubz3Ft
mjzCQiCLhI6qayb1qfUJJC+MH1hdHGIMOQR8mDrmvPZzOkZvHPxPr4KHV9AP9mhe
BCVcHNy+/CiHDbcY4lxwNwmcZIRafjOLpEI96YLgGaFuK4GpoIgQc93egiOqFZ1h
OfDyCdC4wI3isqU7APaxqy5bNNOwKduRLXWsxQtyyIOdopmroC2FgKUZluGNYT7h
gXN0rRuf+z0mOUu6UgQeva+c8+n/2IrzIHqcVvS5W3kZ3cYbcbeGA0K5iIpq+UF1
yTaTPIr5RZ8J+qcZHS0Ktsd0dav+ynvmHtT9a9tsZPlFa9Hc8BCez6i0va9afE6L
fwOyux0K4iBytcMfK0FwtyADE1yz7f0aSg9hFf6gkLv9kHoopjgV8w9xwQzqa46v
4t5pUsPAKHHu92fMRWFTVFvrEhTvYJnGlSLnXmrUAKt2SMSkiZ+J4kukj+njqkpk
bzB1DKwvP7L0Glv3LCVsl2RqqJDAMRIEYaZ3FTsv3EdAZyyI+LZXGsslkyYIty7U
1l5rzsIyYwm50uzGm68fiCTX7E+IdixmVoKP8WOFQ/7bTRtuwHpytPAe3xYVATX6
7gC2PCTmcNdY+lI5OjZ+t4kvOTk8qeSPmaOlNTxgVhRKXH7E7jRrTMOSJ1DTGm0I
4MbJjX0vlPAGzZo20lEo/Jzly/bCszGH3u546QwrowORNUF0kaiIViC3dpBxKRK2
p2LvFIaQsXlq0dJVqEFyFEIFLHjnAgqHPvQNh0LbU9ZihYUJzrMk95NruqOF9nJm
QJEv9cP8qtFSm/wAQfgEnfUcQB5MiTOLA9pa5/e5r44XqZkwGrP+O+0OW+oqNq6o
cwJJWDTSojRFdzZDnTdO1mw7vwuBddMMvtqdseIH6I4bcfBgbFzdSJCdJs49J2Db
JxZFYigm7bew8QjaQ3cdIORswmsHVRo+SBbYiSVDQjFDunYuHMfJEq9W0uunP+m2
FKED12yIESWpk1GAg7pDxH7W+NM0k1NpIGK97Tui3TeF61/vCeGsJ2pLK6AYFTG+
UzVvbBr2ZLqhK9Q0lNGz24II24JPQ7POQovmgbG+jf/9/yBrYc96P2FlrCU+jo2i
CAOXu/FqrFk7JupksGAwOXO/88O5g2AlJiqeV1kuMOBTN6m3OPqOOwQpbMKK9Fk1
dUlsi7cvOkKplEOIHEHrKbm4dVBVB/hwWpzYuLauzP1tQIpzMXSaYue0BrN6aYEB
9WqG3LgJTGabMpygwUrBjJ5NDrcEmErpjeDJCTXUJ9nziEzc0GQR2xD1vrfIdGUj
sGgeAH2VMmIt7fSqJiOoUNRn78gb3CZFLPcQNcFwv+34qnGE/IixT3sJu+HzBkUf
ZsrwEawcOLdD2f/mbmJjjK+Mbkm5S8U+vx36356iiZBDgYn8y6wyYjF7YkDmx1S9
AvP3Tvp2RYx/E7ErXDj7bXci5DG2IKHb8yvKWcinprHijeaDDWx2XPWiY4GmbkJ6
tyRY/YiuUzEx020Ez+w7VrQ7PVJB87IVkoAM+pdU5O2T+DnHlpzrRqmNwO+kMmQB
VOKip2EduH1WgV+c/6fjyQBmQYSznUYOS7mot9afs6Y64cKlJ7qLGUjjUxBoW1Gi
B9Wm4Xx9K+pQi7gkeeupnoKqrqvK3MifXfA9f03b8juFwWd6P/C83jf5aRu/h+4L
j1GPMiCHsBxOEC1CVj24vOqvicuBTKzaDF77kQ03IMeYBqq0cj0q8fYeqMwje3ax
eSvD4Pumx3nyHVPqkphWvfPSx4srerP/YndZa/4Yh5JLFe8vMlDGxY4OMQo/nLYy
EmrSHK2vzPqUIwDZ3CE7mIHl6KjQ9ZZjT+j6OsXRVgxYsNOs462TKdc86psdHLh/
E+lX3Ig0yI6mH4v6/NS5/KVAvzCGZTCIIT+P9RByl8QnMjAzZtWtS0bF3oCQW66M
ZUqjS/ABBHy6LdUDmvArLThmUYfMf7WjlpOfMP5EHvTJBdSVsBo4ZUxYa4BNJ+Qv
183fdYNpfKEEo6T93T2DU54VSGFNNnY04GdQpW0VOpm7+tFsG6bM3V2weRWvFfo4
DDbEOU+1k2ORKruS3bXUH026F8/8LUvOoLm1iswcEmaKXuXbcrmDILL8UaauC8rd
HU3SJrPNLAVBO/rqvEg+PqZ+xArmmCxOu+ItGChYLcOzsEkva8hRNctT2j5dE1e8
eA6o9TDTFtvatypyo7F1cuhNBFOhcWDp2a8WWWssOhyz/7ra+y0Rj1jYOf3Nu3H2
KPOco9SaSJgCj+o2xqMu3/oYjDWEBahFN/fdZad+Dy7dQdbwAQm7QwneBJ+cABdA
c7w4bZaR4ILcJc51fxfXi07sKe3ewZ6H2yGwmhhF3aXxaenJ1wlIyB3UAntpZqom
rJx0YzfXQXSh9PzZrIHUuhWZ1/KTcSIgGHv4P7uBJObRnMxMQhKp6DGJf2KhqHau
c27ueJq3tCPcOHrOTXeJIMJQXhHdvRHq1VyXOT9bUJcw3cxBWjLclpn4OFsLNV5x
hwivxXuqm6BfuH9NT09zvGQq/lfNiDkDewdnfIwscGEtqCbeVPcO3XwZYy0aZOyu
fy62Uh9T/yJexhszSqaPIsUrklM9LlDY1nnfYL2lr5rZoOU3qyMzs0QTHvkKP6av
y2c7TfB6zNVw4zOf/v2VizkD4LTyqZzHSnhqjGBD3kxWjJbPr3MFq/LhbItVbGEj
KKHfw6Uzkq4uBBz+u0I/79HSWRai/fj4vOUF9rP0chEAknPDMJF1nhzOKpp6jFDd
KceEcyMtxemGxNH/MhQ5cTayCsGno8DuBYgFKaQYvAaM8rMbqvHm3qQCG+tEY+V/
V64LB28VUx+3BfacR691CoJ2M09LMu+RD4hIdCgUbD3t2fCPt0p1NfLk99ZywyVX
jjSSbhumvx6iXWtiLQqr3ubAnT6Z5WHptenhzJLgpC9/KYIfO2nr1PZFIE7WPyag
KNQSiyrws4ewfibexnQgorVbYjUszef7u0BnIwBFFphYJw5fPRmIgbLh4JgKbcnM
pdjGESWiF+uE6CCBzhmBmNkxYCEDUqiW3XqkNmFZ2bbM2HOKUl7ZQHa4c8JKfxx7
UvB7F6bWtzyz8rxpEbms+M+/7WkQkidLbbiquUTx+nctbloYYqTCsC3x8coDtb5D
xh99LnlqSifBiK95u1VuZs3aXm1pryQ++HmhGDgQ+vFzAT7WYW40cvXk/pIiVvuT
jKKFlJu/97U6H9ZpgeRA9xxOryQhgpnXhraBuSWHSm+vx87YcQD1uAclu4bheWrp
3ilZ2UJUB80mQWnij8OLnB1W41AvxNkFgOrKaXRDiezTT7MYKh67aEhJ9ZM2+bQC
`protect END_PROTECTED
