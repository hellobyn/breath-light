`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YZs+7Y5CoS5T8yVJ7ru/Npro5yDf23NTJgW21IrFeX6Flti6mlWpr+SKGR7ry62X
kYKhARZ/Gs0wFnyH9UkxXnDF8uDT5Ezb6coDFEwKnceOAmDg57p3ZfzBXdW34716
BL7fvr5kBIhYympFg3t4FKkV/PfyB+8gRGUwRMjag76TctKhAfcb60mEJp+p4Y/J
s83InyiSEyVNbQOTejPsXjstKtjhTJxPbGbjeuES34KCyuqKrCr8jCElmaKvyFzJ
9nzt+j6QUK3cM8VwZkovMay8xG2ADRm51p+bThutno8hNqTA1ZoMlNISEZtEP2k9
lQT2e0pvqqGEC6tG0d6ZRRG1zye8TbNR7FADBUNgNfwL0Sy2gxPhQyeruj8PPkeM
GzgjNFpc69J1/NpmlQa94YPxYf60o/Zl9dI7//nVJiXkm506r54ub/JDpb5rHdML
nwgzAE94A6H6ljSJMJkbxcTRfdgEkQLO3O0QUGWzAIt5EA20BWjvoPhMYU0u3Z0/
7U49WOYXGYCm3fK/1kD38eQme6Ok4g9ep7a6poUfpRgVK2SWGqzUlbnzunLedXNU
uHeme6oCa/9Nfpu2WnWnVBQFSi6A0u4luMO4GWKp8b5LUWYSHTxXRk3oyH8SzFeK
YCn3tEzWNE6GEcRAFeqIcqPXw1ivFaBzmw9RuDilTCAzuZN/WTXo6tLMPYAXtZZu
UsW76ew8vKlcLn6kmLS9VrBa7LbkSN/sGG/6AJrgPH7EmIiWTpqtdhSS69G9CC65
238gMaKCkJcYwj5nBmXCFrqUkCqzc50P2LAdq4VUuJ/wMH+bgi5cfC5Ymfsh/3HI
matp3vAWg4ssU88NC5com7mmkM0Tma2/AM5tSwgJHlQmRAzOL4xpOK/qeirzT7yg
rk/Qvj4fkAggeZ0hzZuGeW82tJpVYznaS376AGoPYPKTYTJYkbFQmquHFJOXuBHG
fi1KxjtGf/FsM3LI39Plslvyq6FgXhL6vYGEQUxDlYjXGPCuVu1m6+0VRHDqfC+g
Hbl8W7GTlKVcrPuidS1wF6XM7M2xaGIJR4OP3W8p/QV/ebP/7Yv6jHWPwxTDU+/z
ftllRdzZBdX6E2d1MiXsTIB5JADQ1SHuVtqQr1nBKW2RcBdRUZnGmrrXlSCm/pTd
K5xbhtlV6bfxctSV8fpXbw8xd+l+1QhHgI0Zxr2E/vP3f2ci2lD6+s/LrSb0gT1f
w8QPNgBImGpe9sNJk3HnWbwxZmFng0jYPIzUgyjAzgZvhyuKuSzNybVScdopSFsO
ZYYCsRwhMWqbKyXoCGEUWz+nn4VMyBBvCDqKi9w4svzt3EQ57JCZK5avtsboSlrl
PG8rlh7F9rAWgkp/xuFHg5+lGH9Ty7S1EccIuZYp9DKQDpq5QymABeGQy4rdlUmF
FWflag7t5oaweCNSSR6oIHRZ3UdzbDRHQw7h1IBL/aYjpmPNWSQFOTR3S44md4ga
31wVcqn5/xPZaa0VU6hXBnIOhAQ4CQARayevnPljwLjl2YWDxvF7ZtBIFeNg0HZS
mjT+G05+kw+imrWdGfoBzwkmiS19F1aI9HPRQAkER9f21TBYKhijAVDZ9R4B5KxC
sCen9qy1t2JrQV6X2umBdD/SKpffBIkD1ayLKfqnkNV2dmQEWF75Kt1W+w+EdzBb
I+wE8gFlD0UXdslZLwc74JK4aKjPOKKAMv9e6xLtffd1sF+1xQrIE7UrDN27UV1I
+OiX6+rhzKe5DRUH8IDSZLQsXRdnGtlyH7uemDAEStM7UjuMgkFMUs6J1M080Pih
t1vS6/bfm4ghqgwmskGFOhPwMgdrDMY3vPWMPA3xGJV1PCnC23xX6r3Jo02kRD/u
Fo1Om03mfFRugfCleQkaU7CXv00Y3HGT8v/4i5KBTLogfyGvS1i+MLYgCCbjJHxs
RWomuPJXDZ07/g8brCDuDk1fSE5/A3xv3ZtIwmTBGrFUktHI3OafXU4gLftTsvqX
zyM6jS3dpdFpZcGATZau1vyRJETu+HF2uLvIDl08+bxwt1dLKfH+IjS5Depy5ojZ
Vp92Kd/eRIiQsawXL5NQoEYIQJJAdcZ7GATCG3+8Y1iuiSLi5IS9zkV2EAx3NydD
o5Eio6QAA2pLPwLQVdIQMs2MqbrqmgCj2yzQMxGEgjNLwIeI+lZCYWGysb02WaKX
tEZPo89LXsLvvvA24bHTVUB6SchITWpnl2+al6TLdxfjvt9XHZpqLgKc7B6/+tFI
GwrPGXKtJe/qFdnG/vVzmUK6zXPpKpwi+YmV1KmP6la/T31wlCOE0whVX2VJHKOg
IU56g6iivm9Hr8JfnlOYTBsq5tmH8l73n0K8VP9qsIfoxDiKAILA0CfFXMbo6k2l
GqrGfPqcuO4Y/pL2oNCQKZTfXqB4R7RV6GisKNKFa6R/ecIHVdD+S26OzUEI0axT
3AsVJNg3z14DKVhYJklQa2GGpUmNc65KNcaa8PUyRLDmQ1K6SRLP3Un3SO/VjBbe
xANL2yNrtf/uZCy/F9pnm5+PEi59V38vmH6aQfaS0tgrOjACyMtPUVLpo8E6ITA/
FwkwX4fIJdvfB0EA8d+PkTpVBxlembAqCeECFH6WKpLJGiSrGx5FGYhUg6ZFwtRe
c4iC3W1JJ0rkh/mk2CeCG4VspH3Vk+a3uyRTTw9Qy6b/yApIsl/5kbtaYRSpabRo
TZG0sS/YIHo3WNdL2mfVzSYxWIVOo8LldRHI3XMgTiBaJiDDQmAUzz5lUDYv9Nwj
p7mVO2WveMeaDFiXbYYKZ974Vbo3qFfV2Do1E/KOtWskBLAnRGBqL+OxfdQ6pBkt
7MUPMvBTtdNkcVedcseSTSF4EqeCG2AtQzMkYnEc+7V2mzp+DTvpIvk8eTprpKUr
yX92OgHs5oQUuHHVKKAGZRjrHuUOHj2NQzH9u8HxZixNzAADmvPNFB0eim7WvaI2
wuFmC3dTCnb86GGnALriYX+myhMptOfgbQxerCaUrRXEEDk1uwo00gfIkUeAu7pO
LolkKKXLFWjDocgWYNtkQd5WX4jfTxdmq1UPRt4cjFuA8UX+9NrnBl8WhCPSDxBQ
9mxmBAeqIFFtadEMLnnAggEMl8t1/KVyqLV81EmE5y9yT/LfsnCQLCiv46C5GC5p
Vy3U9q5kqCsZl8QTk38omcpev02fEiT5uaT0KRa45DXFPmcNYCukrp8iBQR0+cWv
7SFOKczYr11CrjBjxJBI6lI5CSeaMvifgNELeKCPysCXRhN7UT7whFW7MAcTfyVq
8BC3yBFFbq6FcAy3XHFZOI6dTGvaaMDa2HADMV8AXXs4+GlkfjuexY4DfTugErmz
W+GwwMXoag9GijBn8iisOnHhKCvrhzo8JnXY/DxT8zb6J7abPsPaKCrSrY0ziIMJ
/BJSZPlD98WHblPNsfUMfAgEWfm5Sau1NDNax2bFzT3/hBR9oebm6WE2oSJfH8DY
VAHJsZBqbQkFY4HyVjmL+KjPUND4W6MHmAJ2xf6EkegMnAiSIV8AjiDOqOu+p8pZ
YPjw5DV4I8fXd0IaA0NJbjsLaFIAsk6FcieD7qLXgIMud10S3yKdSbhiK91hNBcV
XjDxaF4csKuQPZc3BwMDueH9gUIJC+T0TRpbJ24YFDt4o4AubVaaCv/6zG7srLF9
4AsEF07o6nKhekowo9DDR7Vo5SAh/6IEBbLQlZXO3+94ziUZRbXhmpBHWRlSKn95
rrzWwtegVk8JCLTPJwHH5H1omhih+iaCcqkv2msYYgkRGRDFzu7pgXgaGrqF1loR
lfHg4ehWYu89j9BRkkS01PQEAmTnUjmamhWAGFCGSyHHQiDVpxZa6N8bhvwjTR4L
dVvI8vBAfw63sGo5i9500u5bKRtig/vpwFe7ZhLpF43DwAij3AME9eRLy4OLL73N
SMR+yfERkYq/K+zYW87c1T+tBeQLXHdh1TiWHc3nLi/aXIGh7lD75Y7fJ4XBdu0v
Z2MyBQ0j2AodJqs9uI1lV2oi/Pp+wk6nedmSEd+d0nxozMvxDryE282decCs7hVI
qIRM3q3lgJ9DU/0jsz9eCGmuhf1vYMENjhck1YTRRD4VJd0T/bF0wjTa+RzM6PnA
7o/sm1R6IGCGcueRxreHMpl566Wje24PbV08haFozr1PN+CI1mjP8sUXYfyvD7oK
gRqTZEhVSh8pva952cL2sSg2UMv8uqZRglTQRBQcDCf/WmFAhu+U9jbSbuQFfZMY
T06YTl5VegJSb0sfY2cSZDPoVwIUK/M4veWbQ/gABCsLlSPf8SZN1hHi9spca4v1
9vTyZ3i2ceGRSMYmhzDrMrUAyEbgHk8Xh5dslPrcHoduWwTJAR+d03jq6DXJneQ/
RmkZ2vCfmGO+7xBa2vFkrZygu48t8K9qF7BoldgUQh/p0BcAjfV6rEJZkv3DKwXo
QUmbQBTOTh5TBQqyde5Lp4RA8wklKZHiR+LvXWfARb9eC2JEVZjGd25f7GSnm0XG
NDX3iha9tDnWk1EWDGnby0by6UDX8daU3EHrsMbUK7zR/MkzfHbAicKlLE9/IXCb
p0j2GTtgmmART4xp4fZtYvq3JL5sBJCiYkliCIHlJmSqUIj1qckqq3a4aUJN9Pqr
iBaUpgWRPsgDorWZUwWOzvc2UsGfo8RW5pcJlzukukzYs6J6lozNPZWouvJu3uVF
QkHz54UFZd2kZHO2fZPNkA+ZTs8U5Sg4GSGYIjgJCe5fBCzUWpsu0RglMZePOgnQ
zZvIrTM/z0ePzeJfmmeYb1p7Evvma6pahtwAaVQohvhNoTFM7pp6ulDsFO/rTwrD
fB5JB2v4ixlueS6RliDjuvlo+9lQa6MuWEoDBb3q+9zQZWuOuS8RCbzwHiBLtQs7
ru0upCnwPNCtYAIxDZvYI4EMzlCnMbzoSzFw5PgUvlTljXaTWrw+75BEiITthTqt
wT1qjCLYQBUyDa/nZJsEWiHIEgK13G0e+4ic7bFf5aXDe1LwDyKtIXpsLveQztrq
pIQRBflrcFOzRSdP13529qk/t91fNDJTQo9GKDTDIRfxHB6mHS2WoZVEYPPcsaaI
ze94opQxaPjtgQW7MTlvFX40NjuSTHzJGnrfJDObBGCdgEXG7T4bQdbioVIF82gi
nP3rmWGS6GuBgDXAWVmrvGLHvfrc3UqN2uzflgknPQWM0ZR1lwv+EOReXDwj6wgQ
EQwkhVLLwu+M/2wvH5Aj07SDWZVeTl/2wRILeiLlhHqikwS1xZQVWG+UqB14X6WN
XjWaG0S1ku0VBhGI3WkHEYjiVlA7+DP7Wy6IWt6RM/eYjF4w8tRsDHVtSzftvDe5
SHWr79f37UL62zTDrA6RrlYT2v3y8yNSn1+8knzLE+qVW6mC8l1jOvsge0UQga7s
zaex6FyXPAWCxqHLOpZH/SqlTK3xKg/GJsRmDWgF/NYV1OK7XR3rGQO3xQ1xa0Ep
j4jZwlBZEyOe2cU6HZ+c3MV0TKN8r4FrOEh/rqsE3FGOFqdVtfVEr63/qQWKXfTL
pnGo+TAvq/Swk018cFdrfRN8wWHgg3GoG2sjAOFdLQCA4lN1VTbcX5CDWnaj6CYd
GJuwgEIRABm7CgRj+9Vdf5IN2g488ccojiI4OktQYGnuZoVRpSEKDtGM0kaiGZM1
McLY8DgkMa5OfKikNBmcIL0lxFoJWSVtRoSMz9nGjuHFR/RKhjD8dYFsQDbmVzXC
wN25Lz7dXp1thWyKpKO14Fz4VPhzwwi4gO5wsgYY21fSX/pqMG8385oXfNGjQSeS
FKRv8iAkdE3z23LXUvCoaxs+gqOqOhmGMlf2eC1JawADQL6DPEdG2NCAXhuOgJpI
Q62aEWuRvO+liZmQB5rIG4q1qSHg6jJ9moxpbWuya+Q4mhZk9qr16XiEsEWg8ZAt
XWrVRL2pwAUcOijdpkmrKdovSKVJCaOnYtFkvHEsMFXwlS4pGqdtziOXwrgqdcPF
HyhO9tiCqvgUuSEZ694fghcKzOTUiIS7td/z4b3T6E1+eChHKsff63JvMj+BiJL/
ruMOesA4h0ZQwZtXSKhP7g4e/S/Srl0NRlUTCWR+0UJquwbEzig+/HKfjx8Kt1/2
1RPjNlkIZ+cy99UbSfwJD5u6aLZzK17Lt6bKIDO62bsq/+xblXj4Mk8cr8ZE3CAw
iuUz1HoT649QiH2OWcjVpvstwxvl+HMnj2VxxqOAp4xtBtCtPX3AGNF5LpbXC8uy
mFfPo6y0O5BNro16iioGrvkQ5zKzeXCbOQq4iyeNxXvp1gmixVqJ03CY2clUY83c
sSAujybzf08r3Q/8KKulbrGfRAwOjdB9NqdHzVYLnXuNNpcdOys99GwqKRCI+k0z
GjJJM4szrvoEMJDWFOiv/JGl8W6PuUoeW00l3SDOCnp6XwbqaHnLe24AW7G8Ngj2
63T2sCSBgQsUejZFG8gRvJw1FNcnk1F63kLllNoat9HrRS3Qz9AEKE3KSiHKJspj
LPBYLRTEtQrC1P8TfIZmYmG0oLipgJ1ZhIQ4WaPIN0NPaso3dRmnSpsgDN5RCxJO
3yPCqP/N6fOdPbc100yoEQBcNj4Db75KQvUrQst4uU+BGyc7GHHhvZokRmRC32z/
0weIaXOu48uUg+oazNzYtfrvf9YL1UhBsY+fdSE6nDfc8nV8IFFHtxfi91/pJT6r
VprqO5mtEf4JiJbBiHwOiFtMtSghJGmtB0wJWl9YLktxd85mIiRdJICkH+8g23Z0
YFziFd/oaEYInYkhO1OMiMnoJ/ogf7p0cVgfVll5jL6NeqsflZ7+Vh9TmrFJjObc
cgK18mBJBEgvgxTAEJWpZVqavUd3N/+b9IYetqQKjr+fyNmuTIdP8+L4BFRUdT6Y
U2E+bGO5xX4POgTbhzrjNBY+S+tiygKtzNplaQ90PYo6agQ1vXx3Y21sFRVpJaYo
YA9IuXXjMvdoIBj2eDRJW3PmSVZTThtssxg9/RfVej5Y8GPTQqPwzuVv44JY4xmv
oJYSLQIW6kyfkaaHjC1SC2++OOyb09arVn2fyGaeIRwC0ZWfyprX6tBEb4wCspZE
jS1M0u01vcqhtP4gHQ5wskSJfJE+90wvemu6f1tIQLVVasHnS2N6NyRUq8GoQrab
u+BW6x9dUBVc0NPxoDljhuizsa4UCGLAw8O+UGwdeNnVb780Poxwp9fy1A3tq62e
+kYGk9tWrL6EfZ+Po/7xJ5Zlo+VB4qX8A7Fj0aqnWkuCQW1RQv/0nPWqbu6vVm7a
jj8QuzQe7Tme3MAW0Cdi0HY1duv92J/YcVGbYp9DJ40=
`protect END_PROTECTED
