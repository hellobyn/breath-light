`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kMW3MO7eM0X5igQRtNEjNFzWSGpARlajJc18dwgc2IQPn8KIWGFxXvSbo0cqwOoS
RsMC/6AQaO4vQmSturcI3YnLIpLsKMEE9KvfgrZU8fzbrF+lvCIA+u4aPdivG0O2
hcFUABjN2j4YX4kjPvSDV7YxKSARpdkVOyYQYS8KianVS5XF4CvsL2584qav9qma
4UURkO5GNLSu3Lhb8oX3gDEBgsdf5+AIMrU1+1VSif+yR1TYkaoFLBsaB/+uwVad
jtQNKv0074bg23fLW03sDkpi9ugKCUn5g4NMo1V1LZXxhVd44ofKE4o+p+ryuzOS
8bqolGojcMqJgrp7p3eM5WeZJKtyIQdxQTudbr1H8fKgpNFIHbCaC3TH46Y3687B
`protect END_PROTECTED
