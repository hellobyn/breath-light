`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NsdROcWUxASOc1tugOvlmvy+s650Ganv5xL76fEY5QYreVj3INFin+C0gP8/z4PM
q+yYOe2/wXkvH3tK8p/LCjFnH47/Rs53y5S5rgrhOfajUq3bQBmY1iWMcAvR8FjA
6gbR0yAOjn928vD0TCz4Ajxz5gd/H7Q6XfkGIPmT6SXxDO7XgJGLb/PWONmwcQna
0r+yfu0sVaHpPfw5hO4QuDBAYR8GmOXxcBRHfHe+v9VVL8YwqIUapKxFwmRI2iYA
RjgqG9vpGW02qq1VN9ramCzRYohX2iUqvmsbKPadYDrN/vwyTCc+Jf5nlTNXzZqi
e6RMXJkTVlpAWa5qnLSM87/jgqaSW8LkwpgT0Gyx0xmZoy0GVyyx8vJ0Te/Qq3a/
aB9f1AHwOd+xPvf/igeNfxkVgU5U9OaeSU/wimBn1gZx4cFcbwFFUkU8/wk32w6o
rkWXZquWqjgLWypUOXJU3pvKTL4S6i+z5a860KmgsWOR4M7PcYVDXUfwzk3PgEpN
HKpsPS1Ggswxfc1xYwOfI6XNdMxZfLIpO4rbqeJTzlDEhM9stY/fyfkTM1m+WlNU
EWDepzMqPRjLf88ECmbvAo11iDiCNfof1OCWnEBQvzRhovgBIu8GwyZ0MPLC/cB+
yVqke86vqTqtC3ig3NNYLAevUl2QAUjfrux+qY7sI6RS/Q1c0bZQ4yLX2HaJ2d0c
gAdjcSfqGoHBHTGeMD8dFw7VTzDSX/xsBANmVBMOTa/auCAvPDklRf9aqePCOIU5
WLnGc9Vx0eqSkxxkCdj8SvKlsmucyaED5UIWIvL6JcLioOy2+137ihir6RCIDmlS
Xs+kbol66U5Utb6xvEO5KRlBk92p844o+PepSUtwge/2tZTzzmk8DHJHyonUNYK/
wgMA8Napz2TsWbbcYT8tiuUyK3QCvSqIACaGFiuHTk8+G/KE/zTKcgUSTB3E5pby
nS84LDk//MvM/++rsFjlN36Ivy0kipQP4LYPeMqksq8=
`protect END_PROTECTED
