`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iAJc79kGwXJFWTdV3OHEMAQf/p8ZVjm9eOrJjNb9yccZNWQKyA1KC0lbCNbXv0yn
tBCZqZ527uuC5BeJSEg30aFBbCHDPkXcHFPyox7pBH7A2NGwQ4PtC/Y2EmgGh8d1
0ffM/pSkAE+3ZTKjhg+io5fblxJe9PHrTCyo4jgIybnDN4E4usYdi3VmeZ1DNVps
/tIoZtwI13kfTUJtIa9BkeOX67BPWQ2tBbwxEXdCv5ywCPUeWJTLpO9t9H7XW+3/
6K1sB6UX4oBV0cSWQlrgvOeZqoeTBqb7FDAorAjHzQRtqT8jue8LeLm97LRWz9Sf
+2MAiuY7DSV4hI4T1mlAsgTE4PX7zbZyoiOIBy6KXQBb35jYQeEvrFNtKXpJ36IK
e+RSirF0UichXURwK/bDDso6WXQGEdxUCyzICp7MSvAIcknMEHcPXCrIS7dUK61E
NcdDeKyH1QWfn7cTZKc3Xhz43WQWT5KmNN5tPsYB+2wwP+WNCyfnwLTvGy8ohsoX
F81+l48B1pyvkzR/3gw+diXKR/omCBRLmZBhPsoEO6kN8//DJUodhTtHZyij8QGh
VKeKaRe+BYJmKE53TWSkLoleUeWco9HfrSkJNTtoMrqM7sRmoIeCOPV7uNb82TXH
Y4+45bLG/Mh6YOdayK9td9IVyy32Fv41do+1BLpyFRpEW/LiunNbIGnKYgMjOLDP
ZmOfWJOfDFO9c68qOohMyuTQNRZAArRz6n0EEyTDCRFrKUPjqHB5ObxLd9WA8y98
akCDMxzaEhui9bSg7bGjxQ==
`protect END_PROTECTED
