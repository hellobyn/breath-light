`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lY+qeRTOh0Y7ea1+/yjnh3aMr7fkTMJ+hL2YJ3/FffuhbzENM+oH4a26e8tmi69c
uoP61Ys1E/YhdoLuUZHOHTC5BRoMEo7o5K37MARREbiVrJCh2NPoj5bOXl8zkFeH
tuDFgfyOZGKSOFvU40gdLpxlGEF45o8qzkQ1VBIktP7s0Os4NrSVoEiAXzMmSNVh
QeUXMY3jN2QNDDwqhe9cTCMdJuCjoTIkQi47wIHLEtpdGlNX6687llHoOAD6DiG2
J0RHHYUJpWbHOAKc1X858caG6dxusr13rUi41VOC3wrsc8Ng5nCW+HFFGc/vfU+p
bm2kWE0e0I6zWrl+/9wDOuThfDkz+YCK7B/eFOQE0J+7vQkYqi4ryK3t3c7HLtwV
LfecG0m6vhNWBr8iD9rAPpmmfBPaMfOutPR9OK015l4c3rc3U6iDTJDBWuZlP7Yd
8WSWnfuUVIZ8UXR9TDzgqqc0O2moxeRt+iuDxTAmeVuiT2QZRRscsltPgDB0NzMM
fheKF/o079Pw8o6cSIWa6lQnejhBsa1r67OwByMy0Awub2TxIfz1vO1z5f4g3phj
SWfe0hybWtyErycAOc7DvCpz0pp0w/7bG50yFiDdMoC8MzIlrqv8Zv6Rb71VE0V5
FtUZbPLd5vYU0rOGhN+3XbAYGqVePYzh8awND6xgAc5B4ZHYHn4sssqGniU2wpRD
Vseo04AbITJx8+uhChRXhe6tZeyF+fyKqpZjgNu6DamZsk25cWzgoEprYGkRQNqn
vPkPekS+gkztVNXt35YGGVKyQ8wNu9pPhbav9LK3uaWoBEiwcR/9d+OM7vFsmkm3
a6qbuZjlpzyoo6GAuNgfVHKCiAmuwIOF/qxq9RpTzTVWA2IMqU4zMwEa5WKaDEaW
RTYXXzeUrGaZli16tZL3BQ==
`protect END_PROTECTED
