`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iHibP0gC2wq4mbyQeipzAVIxvEQyllTRm//QrJr5qrQtXmUr9P4dJkurggscaLe
PPDwqCPjUIUBfes2a8VCTqOj1ltR6JiAvyFBGA6nB+L9XR9l+s/hAmF4F4BEopxw
IMSzl1T8vRHOO8kWLghyIFEmaoi47w/qEWEnQAH9Jpc3LePVS6WmX06ydILoWJm+
hZXYYBx4B/qfCgiSKREiURIthIiaOvV9eS0y3zfUoYyshLdOj87zoOnVvwxaM3xq
Al8MK67bXMWSSSu4BsNQcrwgZPXgbT39qfrbybzlZGJJ3eghX58CYNf7YJxO25vF
DPVVrdY53Wwx74C0H2JTqcB+cAm5qFfnneiUqzXJpqbqfQ7Hkm0Tpb6OiNk9A1ns
eq6nL+M+CmJtj5rEO8/gv1EJHyFln/ASNySAj03d3sIal67Hh5S0akqnwnwOGftD
eNEfx5eev1stnIsqaZBVy9lBTPcVJRfRl8CesDpjmebMuk5OEa6ZmowQjBJc9abg
8B2928TuxqVnNTIcs9+5n0VhTzUj8qThA25Px3eypYFCFJmzoes3KXXchwLGmFnk
gUXjORqYhxsquwaZ64KDs0HGzgtRji0ti9gutBtbVHT3e8Cuh+herP4nJC/9kzoQ
7WriuGqt1guWhZJi1xhJseJUNq1pMtkFHrc6OctSQKwVixuTcFnmLVpjNkYnERg9
G+nsn00pQkoKkZrUB5kbvioCsGXIitxeEetu4IdNdye9XpoZaRnUnTVp56+nyZMU
8ScQkZW4fBRsSN/V1XBy1/8VsLtaoSG2DWRkfEGbjxlftKyrCgu2HFg8Amb7hdqq
wiDgm0s8cihtZj8/blMrpMCWLoKBAwc+s1vAxuNx2luLG2GdjG1unX/Uc6nU7dnT
4BkZfLxZI/LpqyKhONrMmgysGk7c4RXlnWZ6IWzToy0uehODx2lhpC5CBPAtHanm
7hwZcyDd4341HaEVdtSSzzA6YE11PQ8l9kLVYeKH+buhvJdSeJ+oI9FkgN5tGMel
HT/GsoOQow8juBePEgmKzS34uKTauQCxhNdLMD50yUKB5w+b/bpGuY76r3go3Lo1
tmw5iErF6iMkNFC5vbJhe7hAJrrn1XaYYWMKs8vf+XUHs+2WfZvrKeRPjB0iEQRT
Cse+GWBieaH3yhZIEtCokUsugCHrnfuisijCMZPnXCeQdfz2sH0aGSJ9CHThdVxv
SylJzdNJRMNU3AH2X9Rq6W9saXptfsGLuCQkl1nKr48cHZmkfXkRs4BJw/bBHBWf
6u7W027Sd0BUtEbDwNl159OlMa69XKbduXrDGFG8ITnS9DKuBkh1gOlxwrAbopD7
zA9LHio+n0sMUOU0W9bGxw==
`protect END_PROTECTED
