`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJIcEY7Y1P4VKjKsyTD8kMULF9mFazRAJunvyT8+0OpafFhWe+F1jbNiL9yBV9P3
VUj0pMJ8baZvR/o3IFPRTV/GPMU4jviYq5yVkeCegq+q5TJQ6Z441p3OONzbMTv/
Vgf4gsiDM07cK+WKTrbsbqnRzV2T7Iy+z+fZcwWpusl2cNo4GLm4kCtmDpnRmEtZ
WXYMKaAwTqxCdv037HbwQJvIBfO56GSXzY4XI2B0lG4Sh+Waj+A51k0wgLPLxjaO
XatpHRew1fyodlrLG9tdaC0EZfIxyYgWmAsJt1L1YpKjVvtHmFKzMTw+pcfpGTkq
pSE7lxnQ356r0hreDhQZ1cb/pcveeZSddTRr6nzv5TxxZtbwuDJhHJunYHEDK2pS
up9nP4v3ortwoharCuQwznF5MHX135SqDDV+uS0q0SQcjPBG5HwQXhf2AfZw6Ozh
UT2atv2/U2mVgcHayDYBwjNDx2XfBUkLEZlnSytOn4oYIXUgIRH9eRCFBRqkd80/
3b9yO0MWlCWcuPf/WZOv5m5B34vo6Sn26UYdFO6c8m5J3S7Mp5aE/ZpZQCW9xbTu
Cd0bQr06iWdr6y+N+Pu3/r0DfWzeK/ECjBCnDRBwzpUjjrdVcY5usszj4HG7VaDm
1ezxji+2islTRDwsv3E/ze2pKgfciBg0fPtZwiEFWO24jX8oENNZ+zQsL8vr6ygT
lbtc5YTM0q9AYrIin5/HnFg/OsCUxtTBc5LmwYZRbS4F3ELs7E2NJrhT8vAdyFWi
nRLbcRqHqfNObzcd587URvANoiKOcIyl/dHyYdege95oMUYgROF8wCRxQKYzhFEA
psCRzM/LcB87NdXW661PVSbr+Q64gGZ3ReO/ud98fRJky1aa7G4Im9rjpKGdMd0h
DCLKRsO5GP+xOxEE2JTFJK8uVZRsGt0E91RU4a7qqoIY5458dP+CdnAhx8lXH28l
Mov3HrSQLaSdpVuANUw9QptOTyFpgZw6z+Qq4sXPvH0oDh9wqOcoNp+8AQp4fMT8
celQ8r326X6HszuDe8nF78x4L5e3LXQrd05rN5SAs4a2VHXxu27CbKYmViN2kBZ3
P/QT5Om/KFTzGv1jl1fDSWZ6tOWBgAkmY/3zcMGh9QpCEbrspKOYzIFCMJh+kNOj
pLajyAB5a4wQi9PcpEb3s7dxCJKzBu1bg05iLlIJPUjH2Tr4cKvmEOmQrlbyrhu6
109SzOwTOjAD8pDSkdAD4oubdWoQN5N/Au9csBpJZO8oHaTjND0eCZu1NEBwnccW
J+IyjHoPu/zkYKzuQfd5W8ppeGjDoxg+Re5LOWpjS5CT2oJI8HrW+vHmNwNuqMm2
MDBUMy/FKPFDVmnT0gspQhMDIbBfxqUm6/zTFd3PWugVi2MDnt0qEAhJZi5ETmrh
DRvgmAEKnBOJupx2QK8Qn+lEpnyMfMSEBIGTck1+OdtfEDkBEBc3yAy19Mv32Ttv
lsmoI3975krqhkMMUxE0ARd8YCs/sJHdzjIgh9vfLXkXv/JvLknaI/LCwvpsRN5o
HARHOgA12SjKMOhzMIXfnc1c+/dCJISDlr5vHgPYLnJpAHSyGPmQG5RVnGmE4xrh
V967mI7z2RKeM90p8NiChsP/PSUHP8exZHKyoW/vwhFgkGsdk6UQjno3amYeNTci
TGus84oXmiPq0fNW+o9T7w==
`protect END_PROTECTED
