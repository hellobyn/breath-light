`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKwGfJ06AGwXd56SV1plQ6p4M/DEGGDQ2BNZ+BgmwYd0S8FCZk3sCH0Hajvtk4SP
pCaU3xRh5Q2EJ9FCUCgp1yNdXcOWVnb1pJ5BssV62P7cM34HF04aAZxV7W4EHeMZ
jwFprcBxKNYleH5OeXg0Mk81xDDvZE+yz5bGMdBCy3f9fL9b9XVQ89h3FOLTYLxX
EfSyCjiKslw1j7LSLGv1q6AKrw6puySvZZ29/k/LzJhrSijQgE1GsBXoPk+LFkU6
omCO7D5Ncy2CFaIw4pJiMOPL9syk1UmZ27Cz2otqCtSscjGZyb4onZ2foDp3g4cB
ZaHagjODAckcKGSrWv5knm+TwoWRbNKmL5XZWiA1EZXiWmRGmd/w1A2OOsntGmKj
7QNeQ7F5PvFZsZQrpDyrnTb4J173h3OzvAyAtEW437pARjxqtFfH5u0pQpmycoy5
YYDFkSx3UEO3JUwf1/wc5t0e0UJGyL6goUCYFSSDKbsVmAXIFqTCGyNxGbZREgqd
4X4ayr2Dtc+FSMp5179+ti3VQmQNG7NYDtAtVzg4RIGSfFz4p0QVXonPrL9w7A/k
+uhlKTwi/FN6JOuAerd9dYLcDMznTzLEE1QJHF5VjaNFtGsfKGBfTOgJl38gZmA3
WkPj+/JxmkAQxrWUb2LniuDMGHMPJ6aD8EnosQN31yt/TR2DvsG4GMvjnTAdvtj9
e6MFw8zeXO3lo4tQyR5KGYvvopyjJSJ++41KKkOlyji+1yAm+Bg9WPvXVwZC8a3B
ydZ9FycjAmI1Hb6O6lHfycF5+U6c8J7zqz8fyry3SCKcnUJvjeG/qN4pNl1FKsNe
Z8b7h6AO17FuoXI9YXsayAB48GcsYM5bvtEXGWjFbSi0Kf+APgop5Aariur9lenA
XPVDudza0sHvXGQ5Nv6igMHge/83xzQER0NUUbx5kShYGqq/3y6kNC47MP5BO4m/
zLBHyWqbky7f/soRLSNh9R6m8S0UcaD94a5t7phtsxWbn5SfIz3reGacmKRvc+aV
Ojgnmr/ybedE3FzapqCNk6DByLSOWR/pvYNZRQ1+O53ZNOnAqxO63jTEMpqFs1cu
MiArdf3bv8z/B5QUuWHJKparibuBcyJQkgK9eQ90ekRsE4gIkLp9sjwrevZpw/Ki
rhfuLJ6rw8i3LoS9IBsYXf3nUWb96kcm6U2W1sOXb43meazsbf6S3eJT+cSEWiVr
aldSANOZIXT5aCRJNxc47/eOglo7sexS6Q3ePQMzPf1HZ7PtQUDeXlsgKW29C+pK
lTkNrINZYX6qgK48PmsTDKSNlazEw/8Gzo/5hoZmK3rOru7n0d6YjBZ5OT5+WtuQ
03/xrN2Hz8u9zAWRu/rfmJ7cy7imDdQmCLEeqy+Y84+z0LXhM5tdcHy+1kwoUhdZ
RKiD4u55i8CchzZKkX197U2bjnSQb5noBEBpnltLhv6gNJmFdexPIoLxxtea87Q5
K2lMwH7Xie+JMgaCZ0S/NbbdMqAXmbMwLpjjFDVZNB7OM9ITl0u4Efs2clQcDr0u
YxIZNCAGCBoHG1c98L51RBUDppFysYxClO68ReXeghes/7VjkvVzStLaiXcRMsT/
uXMvTy0t1fcnULmmOa42WeUyQ/G5sqtgmOKBn1SahwrzdtiQhXOJp7jEIwXnJCUu
M6aJurjbbk3T/BNZHyDVzvzDSrkDG4M03UO8hs05kWfn7WRq7rCSDp54Z/4p7c1p
k/9BD9liGOr70l8ueUgFpO6US2WLiK8A5Ycr/poR0F37APZhfnpqNq6fqdbUg3FT
CjhP9HoyZV6nJKFfPuCd7N65uBYbmMWh9fSbwmwqCkY33ZwuyiXT+wefsKzg+HUw
hphu3Vk2KB2ufVDU4b8KE4PpAKYz+vDYCb3FibFLA/BbUq04iJxHlvEZGlhGNuD/
W2gXVe+ojGirIYzk6tQefus0I2oJYKEtBR7lguJMxl0gZ9MRy01svf81Lkeo8gwD
+9sVrCqV5XJ6hfzPxISI9I4WpJVJcKbA0tfCtAjVywRgZG4mYTuOL8OknsXjJGAM
q5ua3R7CDw2BlxIw70ZtJpL2En798MBa5jFyWDkv1/cdUCCIaXOqUWp48lnrQ3go
v71nQ1S4k7qp1Lc1OCfZYJqhWPCvnR03RyKC9wga07VEnWi0rHm1m+ktfQbuRMYD
Ws/1j5FH+QMKUvV4x4ovZ/ftavK7WCDAfX/xz0Xwv0ortLfqyZSgKLjerQQZdTG2
N3qm0RWaYJCH46mLlLjtbpbgEUcSyy6ybgqsTtH3cfsTSdhR8q8gNEG/UXBSnkgC
DQmiozpu+sIHH2wjcLSlVY14oATmQWRGmEKYByoTAZOkqouzywRw6zKzqNShhegE
hoTH17RhRu7Gozd2a1ipZSUjXlfcbNQWwHMRcbMv7e9/wuzN5+UbfbaBoANPeHn6
WMQKoilmJgRt+Fw+lAPyGJ2SKA46ZMjLgdcVshiU//DcvB6Y7oenrzNOFGnwpmS3
+rzzGZMf1Hc6/Gva7MrCrlr5DP46oSj5/rK8tsmsOJAbXDNLtuNnJF37+8vQhClP
apOgySS8OGeKXqDodD+auBMST+LpoMKBZ8I+i4LV787A6mCaN4rtBObKlMC8YsUy
AK/wmjSqmt/BYnsJ4J1PF0mfEgQUcGiUSFh4jOoJdRIl+lnSpg/6VR/k4ry3lumI
VJ2L32W/C6XjUx1wZdD/XBWqMjIlACSSFUR+0Wkaz7JX4/lfGXkLjdZl5+fT26zm
L9iQ69GcLXouNjLbc+x9JDxyYrfpyVRtitPXsTuZYIJGNRtSWCsTzePcrIZ2KaHM
JqoDrXvZLXZN1NDaeTmQCZyIU5SfGz45Hk/FVlsgOPDdEajMIfih1Hs6ZdQYgK9T
RFK5/2U1YAVpoB8paY1f7MdAVDapfzzhHWEI0zPrbGrrLN5CGz63+Y3TWUQH3RDx
qXm1QQPrUPGLMTxfghSn+OQ9g9B++H1Rid9F/baeYP5E6o5Eq/kRFyJPPfyC2pJs
mA6cnuBQxT1a/f2Xlun3Jv55SjZw1XR2ec1Yuf55oXfJbuzZnVw4qvk9WndKhpRR
rkiVWsvDjJH3yoso94Iq/83GjIAv4S34Bj/a8AQSTvRQQFiJSXKnwEvxppUssxh1
GkwjWqekMn3dstscdn9XxNh3pxy20DLdio/FBvwt1cVb8cpKdq70+kO1AvYBWZ13
xOPHVvNSIYrnZzdFPgL7VZMLoPpj1qo0mVEZ9GmRHNX91HgH3/buJ8ISfyGJ/HWS
RBWL0dW08FbDMnvj706Y/g==
`protect END_PROTECTED
