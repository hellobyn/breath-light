`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBfuA98w28l+mXrZXI8iPJyI17/uAcAhrRRB0zEY/t/TUvZaZpWVk7yatY6Pgywa
eL8FFs4XpTJnqBOH1X4zaQf8f/Xwvo9keUl1junIAkgtQ+mwgQXI0P2/dBsyVNfH
Dcg9lzVsw+nuTBJhUcH9rPVLkDDCAHzAjYLUmuPV6yrKYJV9D7R0s03gJRGetDnv
DpZPID6WmMVX/Jq8tEyZpDaUozmbnAaINfb+379EHTAivMc50TmS+FIYen3elR3Q
ouCcDnDFF3FEijQCe4ZT3BwLi12CcxvQqo82fjlKEhLNgcbxeO0ATgFtMh1NEhQq
R/U83h/RNvOdss4BESfujIN3EGJWLPvFi2XrOPJkE7PEaHFyXDfYlmNQb8sLu5za
u7eFwqhQ6RkoK72B01shF1vF5xU1JVARIgQkr5EF1hfrwB1RlJeEbKXZzRMxbTNv
6qzkuYuvtfMgVOf3qA0G4mGcdwDltVnRpEdFaRBZ0neA6bEmFW+cbFrv8KiNyWtl
uzx+Zqn2gveS5nZ2L35k8KAKCOyqypq7LZdnZqJYaI9XXYOoXbNNhkm7z08QT/zR
XbdoE0SSu/PeY4/THQsLKULllqsyX6QKP1+FDBmz9y9moot8GfNrUd8CwQfUhhcq
nMXdNvm0o52PVhXeeDFuEqGCmHQ3Hqhen8BXQIFM+Xnx+7PNPlA6wJvwJurYuuwe
l9vkEs/R7Hm09U3aZSByCVbybxBG97ATlyhJuukV7cQoIp6Wqf7B9/7swQHKw0+O
+EGmz9XeYfIn1hiWdIF6RNZnC/uEeHVHaSsShn/bPROieUZuTpk8nAggiJKt+TQM
HjNlOeVuiNkwMrYxUdKLTyi3ew9iCxq97TkaXh9icJUwSWw4NSgfze9iuChu/H/X
ruRjDaiZ/RfVDvJx4x38xl86jec6S9XCBTWgSryxhe7wOEMlf19bfCcCNXcX4ZsS
Yt9HUwFemNggwWCTtRPQxlNF39nKJTy4hWRD48D0T0PjHkRJBVa5Axa2i0kjbkFE
0cLjziaXL+e3ubag4buqV8XSba8Dts5CBcNodZdQZNUPSAdfAY16Fy7AQY9hYphl
g4Fgn1zLENMSEtQXmc3GE3dm6+jXwTMj2CWRIlyPH9Tz386LUDzOsBeJ9oW85fxD
GglyFH/sJNq+MhF4dsqVi/AlyEH6f+ODVNEgJ95bm+o8xLeV78QNSCrPQPRE5/2I
kVzbtIgI/Nb36fm9ecHqV1ZpRzn+8FCMDdme7hdV3IvNgyGJFsUU6NpiZhR/n/FO
7RmG847JS6KJ+mNIj/xjhkjD0SUczwcwQgTTNIcV5/XhX4QVcT/ZwwBx7zAuNof8
0tnoO/xQvbiAW5U1qC52iXTHFOFGQw1eZG4OuA/aQkzW8VFuaj3nOlqs9WQHiori
DKV0e/KDoZonRPlYe15sifcY5Cn7GoQ6152hPKnfkDgfDhfCPiaO2sIgzbuvS+QC
fTGlitV2YvJdFcWEpZT9OPNL8ruR9DhN1DtIi1uvhWy7WQMASOMMuBW2yZvdZRRd
bTCcIdi0ysmrvaXiLNh81jMksPLF+Nq0Ymh7yYIZfKkuw3vdi+eHSw7WW1OHt9r/
8Cvbsn3/4EpsTZD0EXt/gsNb9k4r6YJIE4MZ0frTnuRj0eEAOpa0b2TVWmqwOSel
JVQP8HljayLt7RsGXjfqQ47a1laqoevS6amrApPU+i5is2aD8RzrmNXh1zwQo3Zz
ehpumSrvpm5+wp5CR/clsXFh5SdJpRa1IU+/w3DaTBfmfSH5vo/Awvv3nmy18YwI
eKvTyEKjj+H1UhFWmr7y4XKNuR7CTmQgfQU9zjC6B0PfI/BnfDOLjZ6dzNjgkWVn
1J6JzkV0T/u1qTR1/UwLwJNYQNlXXZ2AsDi6tTHaeNG7RAHSbYX6xRmhqeqLLTzs
aCvZB1Bw8/Sb7yf/RG9eCV1cgzCUiWO4OYyJLcuESVUCEFEgFtPvraLk7/7whThN
nnM1l+QTVMZF+rjUgrELyAK0zjc4l8r4z0XsVYhfE5icTiqobAnRXY+p0cM1QN2x
BnUffKauQiC422t6kF5eG5NRyB7oipIrvYSsFvrpaR6+0SichXa4/Qu2gjxcvxDI
bAcMz4eSvF7bNtZYynEOX4yJGSq50uaW7IEoKCIZziHW8iyMCrcm3q+2jwgiRuKN
A8YvtLMpWIc9SGbjy2vGBr5PxMjlDGM7Yz7Flp2SusitBSVKsFenXBsI7qztoY2d
xRwcSmgdgomNUHXbYeCKOamq3X2oWbJNGDbMRs4hvKEWBn76dT4aerIswx2lualC
c1KdNRlBd2T9/YjNMkYxLeq3nb8CcFIxQfeenysH9ZnjWeC5txHDLNZbLyfjU6ts
/7LW1Gy8Xxwdzr37MfDAVHWNMLeXfRIIu6xfSQVNjRzARxCrrNNG9IKBisKpO9u7
xPKTOM6/1q2bgl4qpzynQsD7mEVRgldRmTZ/noAPmR5a/6PD+mwW9sSFDDo/f6S0
gxj2t1xFCZxNAhiRheUvBZh3Yiv2JXrQeSyCP7h7S8iuWsqfWDyGB5w3v85AQN+f
nO/PoDsBPjf17cyfzUlEAMj+zXWOSXGL5QvRBnHfy19jd/YbFiBQhgVIE1Sqc7DY
EvFWvDfxtM35rX7Y0KdE1yleldoVyBG5+j0y3lrcmsEz43kG6VzVV7NQvu/9d8Cy
THCrc5maOut8ajdomXpHO7myOeBbaEMtD3+aD2EmFYOe5zzyd9HGxXf+HMkKmDOg
WZa+LuFw/hFNap+VU5JTYSodPQL/Px9sZd55IowkqLBMSYTBZEa6T4Qb5xrahcwe
0r5oJIZII1NppI47JmtDNxj1PI4Nz1y9JJknDSeHAjQKVK1mjBGR1q8KnZpjipvU
mHiXZybrH/1gtdOR2wM9F28IwqddjNTB9QC2j9O6Fh41eghwg4jiDVDlOI8RRAYJ
d8KCLi+LT2htEFT1dOoV7GX4B8+cNl8o+6+DqTS6h0jNzidz4tq+CmeHAB4XA5WW
ZjkAXXRADSKd/VOtaxYroNgrnT1nTYrxwRE0c0oG/PPgyxJL4PYMHgfKD/kj6cHw
+XQeQgIdk1TUM9BAGSvNYIe3NyMnAVf+rv9+UrtZw22YLgpFGSkYz0tLCnWM/812
B+dq33RySmmSIhc/Te7DDbKirZCrrP3H3rZE0Iri+lcAnh+UAY/7ns6RVUHEdiaK
YJ1kgnw/3UKxd5oIR2A4mkiiN4Hk7xsCTHmkLNZtb8QxUr9DVl258KTwIAOmzkcG
P9YA9pDxSrWIqbVMGJw3gC6w8l8DoIm5v3lT+AoVIxC6iXz2Cgqt76Wj3D/X2dpP
g7OvVV+tw0D0PWP7f9LgR5Xo9vztUpOyvWT3klg+BR9ujZnzQQ2qsnG85WDfMn39
T5R7jbl52pY0eyRCbaCj5fb120C3Vdegx4t2DNbxa17qW1JuhlPEeqcZfs2w4S6e
eP1XWVvm104fA5gwiZO7iRBa+gwl4Mj6hWfTi+TL8f4nXb8OHbCwiCV9HoDak0F7
3LEYC0NZUNm32JkeQ60jW0d4ZQGtasV1i8qNtGrT2JXESCxoFMM8mkEzybMoATdI
2E9B8nB8RlwnKPdZ4kkDGAU6DR62u9VuUUI5Z+Sskwq90VxqmeZOhOW/hy9WssrM
ChONzLlmuUh8NkHTiyzFDEF1OD0AodX9X8T3Z4jWcnHQnaQ8LZFBd37xXGHWfBV0
bXrpHkPHN0flpibzMcipU7qQ6XpYZr9iOdoogiLqqoQeo/vxSkb6wWRE7FJB4k7H
YEu8Ilf6lQFtDKWzPdT9KMXD2Vtc6fpwprrpZu5eHm1X7CxLKpR0Wkt4Jfv71bSS
d/SaVLgbwmJMF+XhFuW45RNplAE24OXn7kEr57prtd/tSodH+2eCwxT8CwdIey0+
xdOamsnCyuLlgizu62QSYEtN4E/pCVZPUcapyWMRI95Dmg0fEPolcUZXqTxt1I8D
k+t0vraq9QOsTKbblNc/YCXe8sjcqJP+awR5QOvGtcAYd6/RFQ7manpean0wqUnU
BA1ohpbU75jRXT5+3pZyNP1SFd2JUtzkek1cagzchWVoAr0UdD1qgdAN6oU2fkp+
7un0RVlnGw3RgIZ0Yesv67ZtbpRtMzc0cY8SsYYD2ChNzEx7Y5/AFgWSFBx9omtI
3t03uLj8XHLOdZaPAXHcqd+TI6I6QggrPif+xdBXAEiTdT92AMvnFrLvVBefL1Zt
IscQPRLIfd814ESeguCALQlQAFNtEhWWVGautwcBb2+zXpUuRpYxA/J8egIrdKa+
PA1f+A5uZkIDwU1Qr6hZzFPFN5g7MFkp5cLMXbKc8ui5R8a5sHW987S+1nHf8L8m
sWpzx0aYfuNXuU/JqstOCl/WHWjE30NOoeR+Fo+MgT9pAhJv9pWHC0o8kK+E3dHs
sGnBFXPu1/3oG8eNLZRCmKMPPK6YCiZ32veJx0iuqQle8L9zDdns8Q30FVKx68yF
SfpWY8h2FLWLC3oWz8FAkyFH0M9nThtA7ZrSUPrziY6vVWwb/w4Ex1rq3wQS5KgB
6kIa4qF0ufqx3wM24LH5FtlwhG7FNzOUAskwJPSoVxHoFiYy21T/OULCLFXOUpfe
bgPnFlq2IkwPv9BWQD88cgOICejrN7qGkm1VARLFUSO9PO3tV+Z/K+nLSfhvEJ69
s+syqHzwAD2+Ysdf0K5STkUHO//olLfI5S/uYDK3iH9aCVdu2kJmXfWmR9Y6crA+
tKviBcsgIrt4fanJ79sOByRKaFXfozNHXVX4HnW040AmXzk9FnSpiLFpCism7V/T
ZBscRDL6lbkDOEM8c9tUpt7mZ7wf8iYdkP/XadB4qTFgTWxPLGaruypHgTjJKkv7
K0hnwx8K/A0FkwPW5n2D8U62NLIqB7Ds/jL+Rpjp0sMiyb0ugr83tG2ZpGUA0izR
yaQRuqmIuckmISkZSxinmKNfPjAtlclNYNbtCGtgdG6wFUGqPRHtLvpmi9TtUKLa
2GtNMVLtPPv5TAQKuuzxnEZNe+HT58kr3lFZw2UHsQOn26SkiySn1tACGxdvL5Y8
wfiFwAB94CI5yEPGnh+wRrD4SANEUv/3eRN0z6KUVksxMAGesplmJ88vBU/YfCJ9
dGR43/UcZU8g5KHaPdgIaAvMrdv8oVRZy395v3meiryRf38xRVMtdEEll2r+lDmF
SYEw3naaFZF6r5GCIvm0m7b3xNdaqaMnoqCrjp4bRLLLfWAojdzbsYp6o7u16qg3
zZ17wnp4FcrZq5LUzUhW1xeVCEHfNtZZgrPmCZDFExR2eeRIB7dD56IXW1WXhlRQ
pGnRDHg9j9yZwb1/QdwtWybZaReE5CKk97RODjycgo5VKy902sws0cYSMh2Y2QOX
WkmD1PXONC0JQZUOYDnpF4QTGQBOw3NTRQUS3R0gGmhRv7qFX3g5wrGIFtdnUojN
bT6aZBHWJOgxQXWp1wxBfu2Il+1TchOIlIl7QfMmc1FxhJ0aq9AFluAVLuigJgXg
PibVf3l+QMoS3rMcmVbVmicgFtUk6AWuHmGCDWqKMNW5VP2vXuRx6ShcYnvJCy2/
/IkMb4/u+dOUYUDGBGkTk/JcD0gZ+qMN2X/c65oNHyEZfn6YyCo3yvRKTG0CSu9e
1qLhBUzTm49CUePUBl98BByBKbxxjU9nyA+VbYJpQ8GbDSyOkasViudUoAlpE1By
4NmuibKhR+qB4FBWanMWhAowB3HYyFP9LyS7jhK4/3OYVSkCJhyRx4HOZTTGR2qK
p8AYn7EKVad2kGqP9LgNxwT/oRPK009Q8/vR7VJgcjKofcDFYhwcdetsfTpvxNl9
z+PUz0cnxCP5n1hv1VGd1ehK1yrBOUnYdarhBPA9zjEeFCmamGZVitodAZEzxOtw
uQy8EhkVVNCr5nDV0WICxNbF2Ui00LWdBegty2d/MrgzTC+VYyS1JSfzW3KFTrZ9
yY2tsRGobDmFO2O30qpWTbjhaTkP7RFBomY1DAk3KnK2eMNktFN/ll2avXQWdePf
R234W+Cvp3I7dRUXRXWhGRZPmF8JwJL8xDSNWjcOlbj7y/iZjV3BlfbbFOVTMHNy
z9o8AtWFmkBxpMOUCyG4tlcR6r22piRUg6dsm/LGbm1hz/mHFC+fQu6EYW5cfamg
R+MJ98lWjiW7/OMcbAdIQFVwy0uQfambiI84tgbbEZ+lOljq+XJEVNB2IGC5T99M
ia781yaFsHJ2iQnIHIWLlRXhJRRYm7vnchq7UC2WfUHMoJnmzbLDaPr839Nfr8N/
NnsJFAIyrC2DylN+dwRKF7ZgeKnOaACQJgNdi41yow2Zb90xc8P+6b0dIRJp22JR
hg/DyPg/FFLiqX6+2D+dT2u+qwqo8I6AAlz+JZtUem4nWunDuR5hmxyCdj1/xZIW
oXJRlEmtUfjln2gp4EQeT18/rs/iRogpUOSR1qCdPp0VMNIFOUWijllHzbl+hDAY
oKQTVhktEOz+ISWXFZXXHUFrZyFCKpbQj3r5yUz/wo1RYfxHmVFtxVxz9+qx3kTx
O9paNk6RXA0JIB/yuUX6XIZdO5okNgQtTIyoHRMHBW7R+VSMgLudrQbiAVjWWMkT
a2evIIho3QTyukucgMl7PPVlt5DIF8WTS9fmgIQ2LJmCQpQLwuL352EknlHZrtA9
xrvGEW3DQxLWKxoEj5x5lG6I8kbsTHDS/c8wLoJZZYHaoHhb2xYNrtZosI18iro6
0QzmsZ2L1dvlTC5sfiSWEZ3hcTY2VURMd4KnaxXL3SowtPbXddu5eSGVuwXYWQyV
I+KKx9O8PbObTXYWkjYfoedxZIXaXYNWzLdXwhrAgqk64cFuzrc9JuKfdnLD5KjV
BphHuEJGlVvK2wNWVaUmYMoykl0zFV8lNkIjRf5wnehybSfjoh+zeRz8h+ZHNtOK
bhVmJUlWk+4kSbyakS4x3us9FOsi/f+DwzpI/R8XUagV7X8NQPGZusmXw4G5QfNR
QXRBOjN6X441XahsrMVZ9IEKg6AM21Rzd7mlgtg1p5puLkhLpS66JIJxIw0BV1gL
QLNIOM8L6C9cpdVQA153i6SDVMmeIjBotXmi1ZBIg5ItzoidKr4XII3yDPAafvJ7
+/PWDJg5MW3T91Z1QQTej30AGtUPZZfiG8iPT7eci1NZUiKqL9L/oVEj06Y6z9BF
BpUnfa4k39ac+exeXBVoBk1zzp3VOfY714jVC67M8MK6IH/tFuuRB026MqbHN1Pm
lExFKKOLuzhrI8WzloP66wTE/I8Dis/Idd2FW1vAf8HJ3w09THp2VOt0nfUNND8U
r948FrS+dSR1M1l1kFQLO8A/mFTuHUG5hwWalkok/Z5AbKulqrQRSFl9975r3RQK
RX72MOOX8FWh9/EVC+DG21J38dIQEJ1mBK7Rn6LaJQoF27wJlV2FR+DTWT0mBeP0
eYgTKgulTH61LzVk70e+xHKyBD38hG6M5Lxj+McDQbrpGLOOYSI9rntQVPE4NVVP
BeOyF/bdfF46WogfiUDXUu/XNE2usSQt50Iod471zRDM6HplgMpx//iYxMsI2yZY
7I7tu+k/uYShplELiD9BIhOlccdtFV/Dmy+vDXDLpgbvxoDek9HBUpz8Db9kGE5D
fqaEedaUH34jCTwZv+S5IMCtOqJ97QdTZ8a5TdTD5vnjlnuU+XH8XDQcvi9I3alW
/4HnkEldw6F3VQmzAy2P/bfbW+N7jGS5fUdSzvQPtqjk+7vobqwhhmU30o6zJC3m
GJDTpk+jsubqQMZdJWRcCenE5ySgi3cJpBkI0WIMzZM5u8zl8FZ2XQrJivwxim+3
He4MUlV0u7orCwEMlTMKRjY5UoBB/bnEqYHOrTSkV9tqYcHOB0X1pK8OqXzGnWHX
MtQxyioqMYUf6s3FdHrlH4f6wO6OLkYN+Pbr5n8MBAxM8aTyAqDzUW6KpVBmDlvN
aasEtjFdzwDYueA7cBmWcy04IIXWJcFLz+WBVpPKfZL6193wUzwGkvPY0Bkxs3d9
2RSV0Aw9zqDov+mrNkzL0I64dgJGrXcixqC7Fy7+h+zzZNfhxlpjHhmFYnuf7a+j
VrECISayBX2nwH4jsM8PgNXPOYcM0jrR5odXjF8x0NcUcpvpsyuvZYk+sjs4XDCy
z9CzioSjFx8RXQnJM42Zy056xDNK9Z0ATXuKW3Y/otgOBA4zxS+ykP3DoFTcm33J
XFr0vtnnLxr2wm97RZud6Ta7nb4bcxu7Qi4cPIP1dCxb6dxaEZq1Q1pNs0jzKGuz
SSkDdigsDXQV/tRTzNRDBzveyNwH/ren4K2azY/M+ZihIUNw9nASj5NGIpI4Ejqo
riRJapSLfcXED4/q/qDVJo2C4hMlLe5KY5X70Ro6BlwAQhndO8KbaXWh4CDpnup/
pKzkJ/AcfICry6XmVMHLBhKaCe0VK4kgImbNXYMNZft/9lGgQfOHOk/cJ0IobHuG
9gIA3pt6kscHN0aUi85kCPugEJuyXQl9bilCMaMEfulRyPMm02A58+XPOYsl0j/U
saJk2NJjVtzewK/r3Jq9qyIQ5WWcImSdBSaWKkcLPVFrffu1TI4crkxlSTEtFsbu
+auzWFsx+scgv1lNAW22RtrRwSptGs6KWwPnmNhunPMVlbmGnaWzc0GIfHxse+BB
QT2OSnd3siVnfR40+J3j5cN4RscJknLSmbUweFnKi2wG8yObOsfQsetKLXN/hZju
WFvxCBljj7HYWfNrw3hbQihjhf9yYOZ99Fiqg2Z80r1GdyC2mVC9U+XM7/jA9r8V
Jzhf3SbUmBwTyxXhvji3kwz+ybeiVtDyx5xV3XgdiIkgGMDDdcwEfMOKXhLdnY8L
xQ9WF6ves3cSR9lkc8Yk3MkAD5XS6Z/mSmvDFZu6nL1MT5Fg3FOn3GhynLL3juNy
3H/P4gIvpOA+V4MKftZzbS/lvphK4IuuXkpUHcupo7g1ZS6L+nUUYYxJJK3OkAbP
ooTUlLj/2Pvo3IdAAvXb6FjL5aTpZ4XN/ac0BNSB4Jn6x+TRcgpHQQBdwXnsK/Mo
zYB0R+q+xtu8o5Vmr+E8IZ0VBxK+yfqnf2MZ2hL+fvrdfQam5xghm6C+NaaD70L3
lAsu169lVMdfck3CAf9+h6+7M6me0+sOTVi2xy7ItParNLg3cEVicpP4p9LqkbLE
glXQE3QXrxATkqH9epRWwjCtSyNuKIO+TxEm4rfJjNFQHBZV9tXCpK5QCpIJABvp
2y4T32WHvek9bj3qPiYv0a7KfixzFcX5tZPczbhNi/i/pOlSLHB6M+9/4XhSUPFq
ANbNs/07X/SjBg4y4cOQrb1uqhz3dfkrps17DVpoTc15XqplsaiJqLjcXZFNEDxi
NAIBBCn4cx3fskSoBCuLkzipkOvqIG4bWZGZ9IZxZZetLfodHNsVFD7CDPoTXO0H
46V0Lr1+IhGUzdEZk8Y8tuT50jQt9gT+H7hYldqSV5m3Xvaz39ODADLA+etij833
TdflHQB7RMzem0AXfXR5A63npM7aTaPjHKLbNgFd+MW41/R/qrztcu9cprZqvVmC
t1FPDtGFQQMbZb0TAiPD/k3nffo3bleYq9eVIFMO6VwAs/R7AFNIqOHW1Takw9MV
eukGjMleh6VtK998aF5CSN7188MPzocNC4d+KGVm4NDgLP0lC46lDPM+KoPamFuo
3K28c/i7BavNZJftEGyVpthoCZORiq98LlOOZ6KPAIhNAgkq2qHazAANLkz/HzFe
hUIhitjFC0VTNiCZ2NSKeAKTBrAi68Y+kDAdQCrP37EVHWq4a8LhN2sA9jmFAQhK
Cxr4LYam1TYe4HmwFP8lJRuVBZwnmjO9iN4LIT55XLcJ7elF4LFTbnkm9aCPMICo
YxpvZUSFNBn7VE4AGW8GlJrGQ4a5UKBXrksFjOLtK8CmY3LRDeqIX48gXbtsc2BN
coS0uFloznu2UG96X1R2LrZTDVIymaZs8AtUZDM+cn+Wqi8IRsT7FU0jpiZcUtCC
rTGmmA3YYjLRpcDNWRC5HHvwvgxSoc08xQkLwDNOuWxh2vSjDSMcVnZ9N4T1Ed7Z
2ZYTf288c8YbwpSfC2yh/hZ2RZjBtl1+HxR7QBwX13faP/vFt2DPuVq9OBaicA1q
+7ZH5V4VBnXFTVJ/T4TnufRP0zKPpIMycgXqrP8m3AqTYE5Bim0fcQpsiqzdTBEJ
tMiUE5Pf0fJVLFIIa4F3cqT0ovSG+SsXlcckwWOhG9u+2WYDlTjqIMRZfGXE69L6
wNXJH9/vLxezI95COmKCIrSim0xLjRXp69jPXfzs2RBEMXLIT/CTcBOnAuGSggfq
cQhs/xQs3kiiil/ltmVwcZljCYR24U7dGpfQfnIi6izhGkSMi0WPFxr6NmlEcUGT
xdlwNTnmXBsIpQBmqxhSCO+RwBfxHAbJYIUGk/DnNgaDN80EqVlpJAAnB9FUlfB5
sDoItDobHZkZcbVmud5iDC9sa4E07WPYdP/+xVd8FQvovjeUVlI+UeHspZ+vWs8g
mreUkarj6mzhYRxf6prNxvft1hkHrxEH1bHLjkWNKyRZriiC/oFYNh6QqJn1sej2
LpViatSld2XASCxP2GsHCNO8dS8ssxiNhfmyOu5g4HmYndghgWXS5puUP9Fk+yl+
ZLnTarOM5LOhiiEv/QoCH/0PQr3u9iqAWfAfdmhiLD9aqjDovGBWBpO9RZzHS1Zn
DVHRrbtcLda+2NbtqRDwCb0NQ6kIbz6Zk5e/AwYUdJdEzkHFcuDzMDM+7reoTAJg
ZLeEpL2e16AUs8p8+PVB7RLXOXWNZgKrUCi8Hotwf0HxtVL1RcEoR6W0AbUdGDbm
XQB1HUffp2WPeyfxz4WtBNWNwMzxBaXiweco0e49LKaRfNQc6u8cQrVZeZ2uYM/5
RNSe0nWvolgeNWvpAAC/7mBax1SyXKmOBhKIB7Ghzv4JgaFC5Uae3U/o4PC+eSAP
hktQGqhIb7HhjFIz6GkE3/mEQgU2yFAOTE7dk21GeGhyJBt4wqNGBoX1EdD+KOkU
ceq7L9U194FNdCx35ZmJt1XXPfiiFRSPT2Vo0Hm76ZxOUj5TlMAOh2dYUSed3QH6
Gf/9sgM8Xnepit4IUcnGBJr2Hdy6CDxGXFIKHyArt+9J6n7kDfSN36ESw51Mr9iI
hkGl4bE5ODXKPcEgpzH+pcTxE0WDrQQGQw0gylLY2e3P4GQxYDIg6HuAWFI7Olmc
Ng0FpcHy3hRseVNlF7s0dYz/Zn2abz5W9LAZmnVQfYzMV0oDrLmZH4qWs6cX6/kF
jdmYJOcUXEElH1v41v8HwleKblvwXZ/GGBn58kAstpGCYAXEm/KSOjY7hFU7GBaH
11phcf6Y0inlIpSWrlrjA8DBNsTU3qZDZoDVMi1rWzHWRqpogmg9USuakfYfTenR
CDlO5MiRH5KY0puKdo+qNMCbkhSeGQ1j23rRO8NerOwlBGyZpUjeP2JKuSnqs6QW
/JTEOqiWk79zHAV32KUuOG9S79RD4BrblxEtSlmG3TZLpE953BkUjzd2yln6fkT6
hwT8ZfHwtTiPp2g05YdBTs/4GKHjLFEEIxjzjLUJVjMCFxmZZkTq2utG/5Ka8KEj
0qS37DUWfGxVyS4mwnhlfCD7aAdiEBPwYcTDNeCkDKtuRfFtcL9Ls7lxT5kspPWX
w+3lC4IOcBDFEakv9VwjlIRrxfURfgAKvbv9kaa6zgRT3z1p7sCxNkdVRWuEMjWO
QEbXUmeGs7HscliNxYp26u7gdCuySKop1mFB14gf5lwgIytBAx7hQAYsf1EhjSWj
joSh/lvR37CxRpV0C8ipnle6GCMZO7WZCOjKyJIn9KgN2jAnWJwKCZJXyxosMlMt
JMDhZQL13P24rmtdmI8vm2sblWApWsxb4hdbJ0Q49KZuvJv1B6bWMs3H0X50JHPw
9aP/DHNedHxyzsaDl5A6CtLxrTOxVoYZ1dSKfi7nNaGTNzeSYagegcYfs+AQNfEq
3eVF3sDh7h3xhUgLNRp/F1/omn5pr8oyFa+x+MnmBGWeUavEPNnQycT4/Inv10Fv
gwC45Kki8QmsEVPQIDqqzcd10dFY/rZ3qp7C4B8tipUViqAhJiQZBkOqJX58QUxV
I4+PwkS+ea3B2yt7zRCp1sFYAjq/SRMW07H5hKeeyMNak2+IeteoZ8eQRCz8oVBU
WcwDsZnroExPpMn6yf9sMqHJVHw4yhCiBZ1JYI4q8HuII/7pnb3sksQQF2TJmm1V
XjSsQTqvygxSrzSwpvDr7Wd+BjUpbx+AvmwJldsIftDXO9JX4uJYMGDSTSQGCAYg
wDGODW1dTawDmoXXH6zEdTDUKTxBZjn13vQAmIV9x7f/k1TbBYqeYKW177G1qfKn
oG9s7Mcrfnrn7kxV/m5FMG12BR8MYn6OeZUvWgGJceVsjOJraIdyMo9zBHjfY9la
a+VdhdCHPXi+gHmK2qXF4DqgmjqQwimOT4iA2aBadfCDJ+E3lhrkmovJ85eWO1sI
4/KKzvw+wpZ/GhYWDJ8fJSE12in2zPWJ0RCXnPStS6eOknJpOsb0QFFvgiaEtxaR
y4OC7sk6peo+T9MacP3zwl2WLsPQIdeBg1CFbCwY/wWJiQtFCT8HxYAyWv9lqslq
6++EuiH1YG3waI9Xx2di4XJBfdIEkMIpHiUdVulPXcwNKl5W769RApha3DEetegf
quyobycOTBkd7qzTl3KWf+xuKujEwO6NE/3MfrClDuW7CHpvRFk8XK+5xqsvOAir
G5MDqeCMNfZQLHGdyp4b4lU+oRdEWVpg6ugL3WQoTLIz4ORHtw8avR+8QlUTub9H
cgl6JbIaOMVCHhpXRYuoLn7JmxICjwMEpQq7y5aDsf6F0nza+Cpxhcro6h5VBRcK
qqhqYJbM9hZIZMfecrnMLMh9FaN8j3ri50MmFY/ts7RoCMVGFCWH7cMOTs4CHVtu
+wK/YkpbD8436Xjtk7CCFOffBhaoUnvSB5aT7tvVw9tOpTX3PXcBJE1kcam25hln
wBJTwqWWO85RBLUGZhe8w3RDawcVlRpQZ6BNnKQ7mc4LCg6I1SsP+aT4IqW6t/w/
imZB1tS3mAeHuY2mfc1NQm10IXgsdkoNdZUt8btLERddaRDkxDgdHsf4WlLH0BOx
afdQsqtJN0T05hrfQSGEBoY/1+S017ktvrupWvO5isTmHu0ZQtFbw8LLr8ers0Ku
NGwylspRh1S1slyURVyK7bboD4ApVYbFWgXHAtQDtRY=
`protect END_PROTECTED
