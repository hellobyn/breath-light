`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pG4PdHOWLTRevNpfHQLkyqjecB8ICfSptQ9FSU/71df1aopHqU+Md6aktz1lF15V
W6QKTvgMh4Guecqfc/rtvBfx1p9VxFCrE1N/NFGWqxFf5dSEbmE/8uYiDmDRjIA6
0NHtGDIGxmKuOgGPbClodXaZixrk/KSe2ccBfjS9iY6Lgnoy9l0U6aHTYV/AerMB
rNnuZKRlLB2N4LxKUThwrksG7JgWTl8kZPAdC/zcSo9HjOrqR68NRurfGTcpFamE
rbdY310hcrO/dIWuU06sLkhmzaLP17npw7+YO1dHHl8JVJ6+YuBFt6wur9cTwSA1
exFZpsnCRib6EEHDx6czOSXpgiuripaMAmwTTpq3gyuVDWbOHzZpH0E0jXAUohvJ
cvu/4iFVtkUfgFJ3DheN3hfek3wGOMjL0KVxhxdkH4ZjoFW8MBerZJ/ZwFpdqO2P
xMSSwF6eZFxWPPybKIcJpHTkU9dN2H5jewj7VrgOsSQ3R+3YBHINkKIUC7rd/pJ0
ES5IhgdkVMO71ctt82GvaPimp2Ln6vOs38Qb9FJArRzNyxYyFoTN17PYLQHmpwK4
K8etfI7z5cnKrAZNG6MMQCAqu5YuE4VCXehmyUQqNbqT8NCajwF4lVZnaLwJEV6/
XEymgUOeFMaZY84UrO7VUY0toQ3Td0HQ4KrPbU2gYuRnxsdd4Z9gxZCW8B6pWwtD
4cnuSIjs3yI+RKZzSuEb9wer/mWWAPGH/uzTTXNSUX3Djm3plYgg7sza/LSgtSwS
hahIu3N7pgb2KgnmvdBPrOBJfE31Aw/sGMspgHRBTnUGkiFkXEsmGk+wXboGh09F
UJ/wBrH5pwVBmwCsNQGlU3PBMAZkIh1vlYwgtHGyPqxb+GKKJnFyG/HNHMVuvzZa
wozrDNWQtgNvx7NNOdiGHcf634jjlVRD85VhR1fRMyPoI7Zj6ZQDc/BGZ2N9d1CB
EAqLiZ/28myPyWDtjnENdv4ehycIyK7qVHw2i8QoLj+uEZ20bOTmaKvkS8llfPY7
YH4BUKuhYgd2mLq448EqrLOw3dCnYQ1awFZvKi6ALFeXFGOydZG5rNJ5UiqnYpdF
nyohiHGhYzkCfXP2E1BEcMXMcfhXJdoBnTStM75c12WoYOZgurBJiaP0jeaBEiAH
yq+aeypl+ehu8x+piflkoVbVK7ID/y+ERdfa+5Km8I+EZD6f6tGQOEkOa5x4S30m
/suTz0WAyai2+bLG2HVhSiSScDaE8aPAriVj9ZwWqkvZwuJOp0iJPIHebOmGrBHQ
P83i8sn+wk4lnp0SYQBMRD23CxVLpjy8FF1n55CTJNYdJxQtFf90L/t9gv9Ewbsl
tm7lFJUDuleI2q9OGNwY7PVcqwxBbiP1Dj6hl0dqrsJuXWr0SSbmQdle12P2a8NR
tWIJo2MyFB3/251q/E+T097U7gYPxw9p5n0nk2kA6es8Joy9I13iU22gb809sOZ5
9f4kyaPqTQGq92o8v0jeC0ID3bramuuqwj0teYNbPs23+IWJX0vHGjqJBxhUKU3K
IrGrFx2iKmaFbKSyubshOCTDeXmK0kJmZDrdd/ln4Ka7SyCBd41f2pB6/F6+mAXg
oXxz3jMcXNUiUM0K+jpFIOmsq9lr/yZThqJm8mfBA+kfEv0jLmySbFoRWua4UVNH
wuVt+QJr2wU9tDZAA143DgmyEoUnSrdBngy1Kk7fIawwlUXHnXO900NHGxzyBg/G
9Rv9YnW6xNM+e5/Q+Ib5QQEtx8ZujyZ1QarNvsGKAFB2JcopytFpsAiNLhrWicnY
9jTiuqYcCBnNMo9xv1rl0xF6ZDNYsfQC3fkSKccnKpDGCQzn/c1ZubJiyHWd2+2j
ec/7L9dxsT0AiQQW9mJdzGxVUklCbREjr8LQUoMQIw08pUc34MVAwqw/MerPspNb
MiaYbA7MKrqV+o9GWPzmvBS4kUZjEtXpFy1t/lZa/T3sCZ6sHIOofaud0wMRgwPa
LoeHhLZqrjZsIVJ/GL4N9siq+SDsgpG+BYnBSoXPJOVmiaf8j8W83a3Cn7ugE5nQ
u1jGPc6GLQX+EURJI8Bmv6d7HKj/nL1U6wCKZayK9ZF66xzyL2r0occV2BN1aCWV
7q2g2Fc+6Ur0uFubaqwo+wJPLST5g1NZlLFC4M1A/jshncPGCTSEfZR2FUG0U4kb
wuL0O4BE9ntHLiKmQ6dEt7nddHqKfultc3+oKoZvTtJAE+OhWQ+LpDUS8q9Hdjt+
qafgoRvW3DJihyenq7HUY0X4UAjLQYleXFj14asKo6aVLfJskixM0g/tgp7dpLHR
+56X89fm/BgFWKXAnoWgM0g4AXzHc7qTbk2HI4pTLkmO/UT2KNUjl5EuaYInplLG
MMYzuL4J8/6dWuj/dA/cOrf492w0fLldMJQbdps1evwP9/+bJ954mogPJuLYyKME
PgqN2HrCLrCEcLIKVjucg5MkKhVJ3sJpj/xF/l5+ITvAUkWLM1LTrTQHVV6mdkil
VerU0VnKJwPh/QdUohfPrJeMp1T0bqG/MdVbGWDZNgzhOKJiWzQVVsMSSvQ8EEZu
K0j99FGk7QR72t0GJJqCVJMvK3HK8lyBHSxQPU/bgExLqg2d8f4OJVEUE+zoltku
GZ+FUH0F25lix5iyqpP892y89o90ploYsyFlAjM9oCbsyUOFS5ho3Jm15/boFvEs
RnZN3XF77yi7Zhqd+HY1hkD9Gb5sYniDK+rdoEUsPycwdGW1TQdAgR3LLqdfCl2s
Zty+gJeS3tWjFE+2frQVY6MQE+c7Br+OeBSQSmjZA6E+iCT5rYlwrMqBg9McfGqV
/7CcFT6aNaL+gBhkcPdO7p21wKm7xdKe8A6H8kNKJNTOJ791wZmAJrxSWeQsvq7x
qPy39Dv3tzIWDsdL0BCt5Qxu6x4IAvla52zWgiZzv9B1xv44aGJUhy5Qo8AG/llE
QfRQFYFBmCBHAioZ/q7JLWQYDjXOiriFcD2DQQL0kiTByaEZgwYJye2Zv3RyMR9S
pU9jTKnxmP7CoKm1r7d84CSgffmanhfQ0DGq2jmx2cl5H7kjBy+5R06qm8NiFpqV
A5W5a5N4BXifMfeUKCdR9GcAH5gGzEERnNDX2k9d7dwlwY78YAqvBEtC5GIwRwrZ
zyu1WTRwSS3a495eTYiGbAcBMinkNLrKzXq8PQ2UtPTY4kXAbnsrr/X7CH+sbJj3
VssyiZT+31Rg6JPuvd78xwC+89kaGOiniij2AoQZeLiCBXcVcLxeFq3/5Qk5m/Hr
uq2MLK7kS0J/DBONDRT7p0MVBGT9O4gAegY1NIAa2jG4R/RJAxHK8mCnWF4dFGD3
rHjtCXlTXaVjU5sqEu+42oNgt0o2usMZ1RzCNkoUtTFrCU80dEQXhBkyL0O4vU7/
ZN2Rw9pkgTXp51af4uYxp0mGOWVZN17IbVb8Z7munzdimE5EZNi5S2Q/Wgy88u6O
`protect END_PROTECTED
