`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOkP/XzU3qlZ323SPVRmnpxB4FCqI/DEOzgBXA3FIiaCfmk9p6mqZomyJN/63a13
C1sAQ/ZeE6Dscu7lQILHQjoNwRc0UXLek/jqeA7+1lCQBub4Vd1Di9gO+JfxP1d1
X5yzJMlolbV9WtYs5yfBSIlq0uLfjv2Z5efY/JczHn/uxYmyoVH0h0hOMrfCCdXb
RcFlmyxNmvVHlvLrHFjc53qWzvfWx1/KOmNVxE2Wne/fN9Qa2E890+cjdAlcNgq1
IP/WgNH5WNtK+naJgipmT5LAlyhorX1OgJou/KTRurrFduDUf0AXrE9UL7hdd5Vj
zFLAOo095E7FVKIfscsxDD3BKk3izmYEjrEPKCcPBkpTZX2fcQ82D4LjFsQqd1VW
qMY55yO9QSc2XSNcFsAK+tPQpTip8/DxcAqBMEDlnhNi9ClqraDhDjNyk/JzJubI
kS057DOk9SIiOrNM74sfSoxPpNCtaaVEEgA4P6iPpn7ZC8Eb2e6I7lbSdeUus0Oa
ZFvsQlVRM9aYruROdDlYVLpv1UkhVkyFcGjO4WeoW4S4r02ilN/yxVcXCiY43E9x
uLIhpmPoyazz06Jl/uggIL8J3vjehjNsswzPL2OTtKxwNKiosoH1/sEa/oV87b4C
GPDbR4Lac4Xo1VZor0fUljpZSJXFJol5E+qxOFzNS0lhUXpZcMa+LAc3Hv/cZe9e
hkefYQADlbKD+/wLlgs2Uebvjx1mr1WSCoqL1veXHEcvLfYlsXaDQGvVX5HpyEC3
nm5i/ZKUGOoLc5A+5XBOhsfDImvOg0Db4S7fLJnp6T11Ao0jkjW2vDxRaoryMVj7
zN1RplR9pGRY1vcqWzS2+BWoAuwaxSMBQ7TlTmECw0Ck0vOZ58N/VVUxlbpN+Jjf
Rzdn8MvwY3F77jQkN38NbEsRnRnSPv71ZRt13Pnymil6m3paEn3liNIlCW41CUSI
0SwSaluv4zdWSKcUeKSGGmR4T88ZS1GX/QeLUGkT8ZxR0m4i/+nSmKOPEVp39BcC
K5tOk18vjd52jmHfw5/e4Lr8PMbwk8CSevaKcgXyVeBpcEturdt2VkjEsh2C4Muo
Oc2ZRVfzH5KJWRSs6jC+fqPbIGo9Ehqycd9yqeuVLVfDBBmWmWQcJptIvRe78am3
jb6qEtzMd+IYck+5ahwotgEBmU4i5msadFGAmcjpll3mIWwrdbHqo/fF25GeQw0f
IiXdmkVFNG87/e1OH9uM3J5u7yoOR7pq7VPAGfMgb99F1jWF52AO8X5UapZP3SpY
XZxPPfOUQ94Lz6MoterejW5B5xxHvZ0msv1pf2sdERbD7K08l7qZ2Jo8s2xYV3V5
MQIb+dPNsP/NOM6hzD/WGULCioPBP4Q9SbLMh3J8S/LWVt16i3R3uBUAZTN5EUds
YsHowxuffO+LSBGnjZG34fVcXEcSFzJWCfCF3VmsJKqtPVvNF3TdgBGCf0aZItRK
+IJx/jMWpYKixldzVSCZs1u675DUoSRe7TJTQJ5P49w=
`protect END_PROTECTED
