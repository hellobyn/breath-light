`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWjgUYi9GV5LC2Gt2NrsL+k0fsI5GL22e2uGKYdsKVBcV/tx6t96h1r/vP/L8bB2
6yWitdZD5Ai0XLjO8t9ZNkmNrdjoUtEN0KIyyySJ48sbjUmcYD8Lgga5pJtn/YtE
8T/yceYihax3yRaZzd2a14AxgYg9/V6ji7nwVyKn/kzFp58mcq0gnqB46Nt6wMsf
n6Qyowvc7kqiQaKCPPzeaNBNnryNXjnR1pKa9McZTW61O/yvqIwui9tEbt3s2xUk
NhrfWVGVyAs1T1RX0G/RR1wd/594nCXawaNH7qb82zVy/J7/z7EiVFGWQ7glhIgf
XqdtITtoPXEhxwKLBdIpz1H+Tbqjg7xndSjujWBct7zh2vJ5Bcsuz0qJ5+2xgBlb
2QS9wWaJnJMcYNCN0QMiG0vDjUB//kHCmkMSYQeXnl9b33Wlgi44nhkwWpPCPMxL
9lROZfujPfoKFdrE+4iTP4T6eeXNUnBOJPAkRTvht30K62uZ/KgpKnOP9m/AfV2b
VaTY0yRI7IuVAPQK828uKbAS2CKKp7BIAq+0eQAzM3Jgwf7GMARud9Mlgn6qv4uA
liLcHx/cZcCQPdyb965chZ116SOU4onMa8orkr/wWSSeizrG36Xntelj1TdHbtya
yvaSPQCGxqassb9/Mu1t9HQgIUNv9/AnxN59p1GVHdJHHcwhx6pMRNMX1sP2w5eb
dQCbvGYYFdPpI9/IafTxtmC/vGGYU+e3NK5InxDbFdNgwsVyGiA5JF4JjpE8609n
lJwTOwh4FlmLTtHT4ll/quCnHVsQ4+95hq6B0+kG8Qt6TyTvXBHzoThwj5dhzsep
+q4lr/x0+FqiqMO8y0Q9tQp3h9uPMCppxiaGC+urTZkkM/zRFVkE90LiQ5PRPdJQ
4EhgN2xaVkNOshltP1CtMNhUi/S2eHkEpjDc1kPO9JOkQWw1LqIaqkr4dDtDE4oe
l5yjBE7jMlUMxhghus3NxENtvAKhygh+lwkKy5Kf1NpA2B5R9ujVmqrm1opY3WZC
90TRZ+fCL8xZ1KraF33pcIdYVnLM3trfY5uXnkAOTUJikzTIjRQNT5nlxcmCWqzC
xr5ldcznwDUwJpux41S+hHG+iLGJB390J38Hiz62AXG3Gk95HcjAXLSS8CDpXf1r
bpPYYrLO/H42YfZwlsghkF+xRAuSLnBmRmBhfT1RmHZwK4FWECL0GJ7ktIdTJi3+
CRhOM1oPclJuUMmaF41ZYfDK5bhDRrKCEVk+DPrD53Vg5sgpjj/uSdIi8azlD+i8
Sza8W/V6lXOKX0QxQ9bRoI7cMfCD1jmblp+nDOjyHY4oiCaz/Jh0T2ALG66bPLJb
w6BdPeMRbgZcYhXsigkoOiWxN/yIWywfyXY2Ru+ZssHoUzlSdgRWfasx2qhpfW6X
sFGsuZEfiPvEDv14isdKwkvToJUvPag6oMTXN+D8EPE6yPYQKgDBoHpBcymxYw+Y
7RcxX1/0ZAV6Rm6Daipepo1xk6zDyWvZqa1S7obcEnBl/krh40AFHWLQv3due4as
G+r36L1gfrAu09KVbWD8ft4gv9HnadUn+byk4x6HGQpFiDaERYx6hbcEl6mVX5z+
UdyJI5zBkkCJHy9tDn+sag==
`protect END_PROTECTED
