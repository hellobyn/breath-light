`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pzHSRpkA945KzZL4lEhMVMk7EGxxh4vTWH7RUcarW8pEchpW14IBAtZgWEdboEO
7vnh3RYIPD1MArB2l/kaqznXgQO+g6di7KojcacXAM+d+1rttL+e+VDxI8dY7ard
uQ9ahNQWOurYxzOZ+KRkUMz8B7eqh3dbGBHLXwYSxw3TEiYngm5/E56Cx+Y7Ktqi
8nHkjJDuR8iY8JjNkY1/ZH6B8j52fc5lumKD+ou5XxeCrnw4E6gByhjG4nCunVGA
v1y9rpbneAghdackq5e5lpBk7RbikXUrVVCHbf17XLTiXFGpmSoCFqtboC/1mpkA
ezecYYjNpVf9gMJSNFZ/lhoQRQ5wGlPpmM9T9OCjLzgUvX5cmWsMMUarJzlASy/k
CgF8M7U1bcedYQe1bFFbPFbAPLkSjgQ1hwPV8Pk7GLIu5lu5yJK3tx4OeEA4Yzln
JM5Q3HI8xAbEfnyCkdWp6enyvzUg/194ZBJxqfFf41TSgsy030Z4YNYDLTNrc2bN
3LbWSufF44qlAFQDNJr172zckMPt+LkK7v58B/waBWrDovXABw77i3iJKnc7z90n
zv2gA7MbJSM8V00U2C1utIoFneMLsLHbU+z6jqcjGNATTgJxmts4Gihy6VUDVrvn
fWo6gaY4CRv8v0WmeH3xTsdV9WRUytym5QWowrg30N9aUwxgxOIO7S9M3ybqPv+t
wuuGNEs4IMpDxwnP+PWpp74KV851eP4o6OSgtRacMfi06lafat7oyr1bgqoLkA60
0AROhZBnV/IIDaCpg1pw2camkP/xIfYIvrclu+bWfFCo3/OAJ6EEQhWJwR2kmaGi
+LWsUAMF9K7J+7SgeRMdva859k9+lOiRQiFnHP06ieKFuN81geyb9bTjW+35omN5
DpM2xd9ijn9GoleLCBV7EiWqwGGZ1MlJyK6g7xlsmh6/LsS1ZjtQPvcPMTmN2Izw
r38ZIENcg+hBx52rI9S2OnVBQoyM3/Vy9YZP5dfzd/vdYgPRTmZ+ldFPUB33Xt0o
9gINnesjSG3aJGY+OqXbwpiHgY2r04ctGqv6xRCDpAPF24Hp6DxvPU2h99y3ivWJ
R+du0asiN9JZq/uGK6A0Azg5YxrQIBdSY1kPOFB/vls8qln6M3OmWBjzJMUN7F+E
uTOziOM9K9M7pX4ncviusg/qR6JJjF40laOkv+8rzIScPBcp0nsR6nNFq7JnWujf
VCKAhyMlOvPn3qKMBkQrnMnTaXP3MW83WpbX4023YPZzgbDxOZGAYPU0BcKbL5XN
hBr7U61B+DYk+P66y2pZ9+1n5K3he4nvTwDGG9Nea2c1Pq/YOtdQIhORXQd5TRsa
ydtzVgVY3Xo4xtHmdT/Xl9JES9u0rhqeJ4lCyzOAZS9HnM2dE9GTwHkvTYdf6NOY
Iko7ih0iWxWmKvmVyFJqsihJ3YuAPh67eITttMg5/KjVOchZyMtiNvXa32qgWGvz
3ndWK2dIR9Kot22MrO8jCOoeFH1/qaX+NbFl0wxe8O+0rQIXK/p5JmgDwQeMEOMw
JKM1RUXpVWQ4OeKsJ+5gKCNX2Wkny/jsX0iyPizEiR4KLVovRxE2A6fFLkWRcPOw
44/XPxNDtQ5T/OzuiLcvCNBzcmvq45vZy6zpO90S5Sn4OjuKbe98F2G7NS72VXAV
lpd62kkSnbSyB6n9YdlkgLZdWkr2jsRdkNOdk/XL2wk19ulM9qIQsWWIJ7SoHHxf
wsb/yE2zxr+0QJLPdegWaYsybKpjW8Fiv0xXcE1yFO8GZbtnnRb5dKhR7Zl3e/L4
1j5HN5kMpIm7eTmay/rCfRRhvggaIlI52ofIJINaBMIrW2SvJa9qcNKEvEcyCsXL
+Id4EpM2K6p53bWsC4O1sPTCIDZIszl4p1I3QbSCUuq9GiPVtl2f8ZHo8rzpjEAH
ptECokSsLO8cRdQWV8SGDKNHuyZYCoS5sJKoGsBkt5TOvNPETYq/wjMyL0MAVHOo
H5Q0nvdxDtJCuHs9nm5Od3DwTZV0xSFKY5QS7imQrHkxPgYCQldKuyXr4uA8A2Ep
reGowo9SCOSwC9Rg+Ygqr/gT7IWwpcQcB6F0m5m6MyS6uWcLtzO4F/d3teu1aJEH
EfSmUslzzkMKiw6Rv0csuKE+kEaqenoSXOWsrqIDC3/LpwYwqPsAUs0pchY9bn5p
Z8iPgqMu07vKtL9RMF1jZ/tuxaxBhT0Mr0V9Idbw6d+6MrcJvqwIWs+VsKs74o4o
L7XpSPlRegiM2jLwshHZsDz0CmXJlXUCWCRppFgIZq56nVUc9aa4w/J9z2j+vS/7
55YhDZPTv80JBVXhPfVbnKW1xfIQWsZVcPD+MxuzllzxqNJ3ylI7kJ2EIO1wM2P7
iN1XMhLqrFADy1ON/9jZf58e20D2i+KhCdEv15Votr5jiEtnWB75yaF+xjEZvfWL
YFt+MXTMM/ISjNfc2dcrz1nZW/kSlx8gcY9wCFe2OKABWyMPhV+z1HfYFpehcTBS
yH3r7x+3whL4Cgh4UwGDOu7nnWzhiMDS+K2qNzNAvfyxHeEQdq/78ROonxoekukg
AKNknMrBWYPqD6OuUqNWc/iM9KCq323o2AhDn5xlNzlkOfSffkx2xVmXa1+8LVn4
ijfxOZKb1Uw8IKIvnSlvDzmZgg8Kv4U3vWzyOSxNWrm2ikp1xjxWkPh5WQ7BJlhh
/aWC83UyQudxdZayOTamEt59d6tofAjvQv2gmiHQlCd2zL72+da6Bg0KuOvs1+Uy
g96Hw4VCUnP8iWlPaVB65vFCKj6t0R2Aaq6kUkos1rMbUdZq8g7zJ1MjqxNK8v9B
5WdTr66H31vOviTyZ5U8UUOqEGACzboY5UUmiVifhayxNWkjLWnZMzp/9Y2cI2Eb
+NAjc4pdf99S6jHbHPF0YZsxxCe/kSCARyaQ99kUrn6yBgx2Slz05UOWx1vPLLSo
ezG9VIQ5AAs246Eb5EooGHFMm5Tux6JqgfOKl07a+6FlMxL4133HRUI8aoY7Tzed
b9OMj9BEEs2YodAAB10x4sKGOWtiakt+qCxb2uvllz+JZjWPXXeVBEcjSxH4+stm
ppOUBDTJ/5hiUxGbp4LXCKjjg9yNbrd5zrNtUXe8P8X98kxbWYhiD+8nkMlmlcx5
B31GuYTWmqc5u0esjWM5Zj5dTrP1ddSUIJB8wWs6mmz9AhzWrFNnvHPEev5QRece
eTfMM47CTWi+twkpb4j9ScHleGSPdFCjVbEz8IhIAZWzsVDEiuTVsmBSl/09uSOr
CvsKLgYG4Bl8JtxbhXN+8Jw7vWkp42GjRG+37FW6FKPWiGauBMJWxFty5k2wGQRC
lyCPeInFucAB+bJzQh+oBJQ4o46KxpSvhl1WeYUrUFUxttK5R8vA/01JPJvlHEQo
yhXClZsYCQKWwj6RhBYHmWMakjX08MnND5hxXymIZ5AXwTj8kEp/EqI1trB48328
0J+98wYLgH4NbzfsjRBdkGNXwSNeyj3kYJjDG9ypNsaUAQDxf1hSKLwp7sF5UFlY
kfP/1HF59qVOcO+we2llf2j6eaBHQKpL3ZbxkMxUKRQpDTuHt6YX+EFh44nwVy5e
lI1mjzwRQnAtFwAEyRiEsTVmlaT9ociGhfDHZwiJgnFGUuEzseV4j+AmYkb/su8X
u50O72ic5xCrV9bwgb3k89c1g1SLzvqQM+HdgwTtDPqZEZqcoPid01Lm+Wq1RY4U
w+TNreBAKTwfHpc1popb/BmawDKomkW3xZkuAxgqEvbDIhumk5HfxXeb9cZk1xiK
+2Lr+z50kvlZpdAnIGndbyfDIZrbuTeDSSJgig0BsMMZiGdKyJIv8JaMwzqo4oAS
ST7d3J4/PlL4+RraAlbZewc8d52mfUD3HNRpLoFhmR85/yGBqKPlPQUeN2UmSErM
nY7CXeuY+DysWwzBNrYTXp1++DZnNAMEzaKv2eLlEkH0FR2CTFW0biJzfHdhuGJM
QCPrhy9gQm/hzyoaOwwRsXAjfRxQWJTzYyL6euKdrqLtg13T9tkJPSvUf1mr6DjE
3k5I18NAO5PT9mwXdlPUOfzt8yMOnoTmk5L+q9xN64dBh7kwLk/Xr/xc7aUHAfVV
KNSHEF+LIc4Uq5cA63Pm7A4jKKz+PL1EJJPmnn1pUMq/ca67Plg9Em+gblRLrkmK
c+7uJX7K0XywrVgNvAcutkTVos+gMAbCEL82busY2x2y88k5YHbM+ZyK9gBGSmCw
qdya0zHwzoWcx6fTSlcDZcb4yC2ZBnWR16lAg1lyAz6IiLH5qXUfF4cG2oB6OIvB
t8fbyN8EgK0N2KU3frnflZ9PBYwJAmW4BYuKCcDVkzZ7EPoa/GpbbVKkLrImOdVe
eK945IxjOS6xmQOjs2v5sp/B5r3m72QXL+Lmlf2X66kPFfi46Oj9f6hBdgAucMtV
eijEbi0y2RF7qJHB6UslHtp9yIRUV+Zr4xBdFok+qc1HyPN0yBQuDzo5pAWuZPOp
q0FRvISmZulIuUExdH175EzLK2u+xm9WOBH2GvreJ3UeRjHRZJpaAu8yotsCD8Uk
itZUdlbIr14G7D9HyEBOX9MTl2DkQ0yONZtMP7AkP02eDrLYlAWCLd0ZpBxwq6Zl
GVdLyJ7nN55+R3Evi5gVHn+DnyQPJ+zGdAromtZDEfzXEIEwDUhPR9f0C9ZxAGLV
MDY/WR5cwx/ilpF6jhTGwP1PgvpCYFtfnGkIjaKTH4P5PfsDCo4DhAQZUdFjDflM
kLf2oduC1+XJcqmJg42nE4ircLZ7Ee20sCq0L27YPHR6OhL22C2RY11jxtyK4zKM
yXZ9561Rie0RRcYwGoCSkml09Bg4GDkui2M1w2A9UVhwupYEEyj58anCELlNw6Cg
h5emgbCyjfcFrg/Fk2iEhgTRycoUvZcqcnBK+ykmfPozpKQC4xPR5O5agPaaHbTW
QaiskyQ+DnctZnWGN9BOY77Xjb9sLxd04Tt+XNIoksUDgMdc4eC6C+0mjEuPSWtR
TPaQ1iNDQDGLz98z05+uPXXQj38u5280WjCIte3karmnIjxCD2nzf1WhFLfPfLr1
KOPi33BtXrm2Nm+u+vPjDC4K2MjiKjr0azsA32Gfvs4nDaLvW1jZVb5KJo1lMiBC
SGonFq0410NSejYT/oLG9UZzQwcGjQocnSuRSbb2Z4NjSuCi+W34hqcNB6cVEsZQ
LHXn3dAyKd+5crU3uBjGwEbnjLRlxPHEX26TVKn+RmGtLmzGdsVvJ2o/Sr0o8EGm
YhPva7P4iKhGXuD8MZKSB6Lrdfj7E1L/9TbIuDHsGijlcYfnBODOAAuuhLcSW+IE
+qIT2n7HmhXnqarCbwUzWDcjpc+cPcuhO9elkW2T3ClXW6qYxl0c81UCkJUj2+4y
a6hzunLWNTESx6SuBvSBDhEXGF15UuiWQAune98/SD6eXCiXMSfjKGGoG5c99D0r
d3+AkydMIiLLq8jNEvKw8JCn3+IHMVwkX/JYdi2+A0sJ6ZJ5g/irBc5TbMqelKdh
9akV6joosWAh36DvOuKSyOLeacgNaGgw672Tk0H/zIRzGCZB/jUJX96NW33nQ/cS
9FzOJYt40mre008eVCzHoy5JABLGdQsPcw17eonRFAdH02r75Gevxdrc8ApupDGz
VsialzWqEdSh/a/oku1ditAi70cYvZE4WJr32GC0teR+GFgoCyg7i7GWLi6vCazS
BAIVFq4oPd/YDSRWppLYsY7ikdI5vxMxkyzqh1qSARKM+2p8YBVBzyn4hnwFuw8g
4g5LhaPMDDEsS5B4fCr1vCENKCV/UDqfmtX1clJofbrdn3M3C1SkB3ZbP596cUGy
t8QiJ6QgWC/tNt88rvqr9wQaE1KoWGPWLgpePJwtNhjd0W0Npsm1RtU8RIVLi07d
ER28JExNnfenj0m1+RWGGxArYA3SEJnyoqE+BsPuPG/jJQk1XZSaYAwnWPMeu1VP
aT17hKm1JEiLGMzPEeHp4HCcd2TZDIu7cFBr4C0gcNrUUBoclA/lUJrEckwaey44
rxlRlQig5L80z8MplB5JY+jFLYaIOONdfXmgyMa6DSHlt02MTKt4uJVGFgGdbxGf
9pPhdj1J5PvA17GiSpsK00/nQphBhJ/c+SPYnFn9utD+dRngC/7ujJQLMw8AZrnc
ajofvcyExZgv3PwGz7D1Bb8HiHpUIfMagZ+iPat+1iwkYQnOJ2SlWTQAUK/jHnZM
JaQV07OYL4gvxwTWuuixL6SD3H5gmoLOWvssohMvM6oCDxZ35VXQ7yeHjrJzkztJ
rLPlUQwE/S9BDxZM6Pn/v76JmtOWJ49u/+T6XIQWmcP1Uwmy2ghrbOxYPVFZyxhC
K0kFPT7M05gcCsNpZQKGJ3FxMqeKlr8LTxkUpo894GI=
`protect END_PROTECTED
