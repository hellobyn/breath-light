`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8shNyNe5ynihf9vXDa+MtEuCdACdKMWPT+8UMvYcdQbNlUxzZEAcMfkIV+4UEtX
txU2vpDVsU+bRNAbshcgXUP9/o8oIISbeudLqm8+OvQlGcOw2ZH+KgLV9O5SnK5A
0D9mmxp87sxSXE/6SwpoY5msHz2w1/aO3MGESWyl/m3YDtYmH6UbHIIcnMdD+J0g
LE+4hRJFmzO9aTp31rLnHHbwVUTxfTDXbzQCRcwr1Dy1kKRYFenjusAcGJ0tN8w4
g0hQxlID9ijbdhXgbG3uhl8mFRCPCH22Ri5FwSJGFZBYwT8cSsily0Fkjz1Hq/Op
znoODkX60REdPkVoKNgOTeADWn4MkLyJght7JMR0IdFmu+tNSMXbnQ7xZ3xXyHGF
6OLxL2FGMJm0hf2zZBvL4Mbq/fNP0bWyG2Gp1X4UQVUgpHanhp8isc9fITFJFLbA
ij0K0Xq55B3k59+slictbX5iDxXf/f35e06gnOFjfqHKueCPLV07/woox1ug37e7
eyICi6gIPnlK12ZprOiKvf7UW78Rz0bvr6tLJpLKvVie0SY8lHCOFKQEsxe/+pVs
FHN9uyn1DATa1teRRLlMen+ZF8TY/Q4WuauPzMjCw/1p2ce55+x663pK/D9r5qhU
6/YlrQ/PLKbZ4wcw3K7T4I1Z+Q9ZSnYdkPunEZPTl/oRbGPtbMKrNquhuEuL4q/p
12EBHxQGvEYMzKC7dHvVbVex6HqPwNx8+VgYpWEPpjrOrif1fPK52apqM4n4vJnR
CRxP7fQUfXPau0fPcTl/z7ugGo5pTKjEhljV2OapxpAuJO+rCysLTn4tukzzLPc/
pjm9gnrTTPofEdXhq/FxBSkMEAuEIX2nwO/vWcfK3Ek=
`protect END_PROTECTED
