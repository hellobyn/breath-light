`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9cbilF4+wHf5XSR2O/NLwE0dRSP7E8T2XxNKaaGQ0ahsXSBdPjPAXqLMP8gFhYo
QNMDRsFyvNq/xgQW00OjFpiViyGGHUBozC5Xz+GJYZGguSoJx4fKmXAfRRVK69Oh
87JWRmTDpL+0H2JTepmNTKOIAcwOeQhdlVHX6bfSspyPnkfr4Q5IC6SqOTtmV7d1
B91EfeTqtTLHriKyp5NgG2JekHi40/7dmpovD7bzjwHBGOf62Mp3GyMLL98PnzFt
3nPsh9rpVMXT+ptLB3KJ1MQVOSEdN0RBN3fMe3Um8EzXRlk2VXUzUIy3evI6cwyE
uyC14VDqDnk3mtFmMJy9ZxF58P9aIaqLbbiOkn0MeHlIE+pY9kEnWqtmdGYReLQZ
fPPiU5SdDZYNE0RXUM6xSwV9RrdPBABWl4j1V7RaSNzs0bNOYjitUMpqqlwSBtt2
ata1ogx77VicmEn6iVkevHzqN0KzB8WgeYi0ty9UlGkqOfHEYbMzLptKMaiSup4I
ZdRLWHOuKAgTWoGUa1J1+2mUGhi3krNb7u01XQ5mUBPXYbn0gTlzpHqnvzsysjl7
YXCEExq7cjha1vTngoC7kZQWDYwT1rYprNu6tV0PImkcbuda8koJNyNdLvpgbztU
myjPmTOfKyUG/Qs/Rn7jm8g4cm9IVfsHJrgWYBw35Jr7OOZRU7iHzxRbJm24sODL
KYoXcBJWNp6lfFLYUnh9yUARtnsMGqTTyQVfcGmEG6iCJky6hKGo7H/KgVzkom9C
88TLovyO2hj8GGLlTMwJCNXU/1ttz1dywHOX0ijjycnF3pCDRyZVQk8O0edg8TqO
UCBJdfZpTE35u6RzOo/Pllu/UVWs4ub/D6z0XHd1H3VP3eobUJGCwthh+lcMhRiR
ji/eSybUUynVThbktu38ZS4UoDRpVNvbhALywh49Pvv39dzjkgxbdTl/ng36s4m/
KHpRVJhH14hNnUoDNoTG3i/jlgqBaGiKzPLCbdbwYE6lvLmQoMZAk75pxS/JqGyy
8R23oU72yQTL0Dt07U1cwFIVL1jriQ22SNGbgthqMjIZ0qo0wXRWgW9E+arOCGTh
P0/Tb9kMhERVj2vkmseR+jY4v/ZUFRMHzSjJWzFOq378hP38MvJvdezqzKI+FHD6
z4b8GkvzSF37HKFTZsTuAspxQ3buUEVdZPP0mhjyUy/xDnRrMBoaQbiedBqjDQHP
obM8W/m0wMES+ZYOSbr3Vy+oK1dNtfoAL7s1XuBCChOeRvxY8m4neGdIvXhf+Yi9
Agpe0CKIDHEfs/ish2yjh2WpYz+zibt3uJEuzfYc/WIT7o65lwUm+GVvWjhjJLXG
yYv1FXVTgNZmEs/q0/HZyc3p0SOXXvFtpr4i+1Ox9holE6mCqXM8crA4njA2AOrg
YzlPpYorfYTlIIRP+oPeOx+uN8gCCHsQ6S8YODsMjRfV6oDPx1aBSgSGcPtXThIS
L9h6fZVHPqqyRt0YkPEmZ27LQ6HbRZv3wvjxcqV28sSW8P0omKE7HPE8sm2Gu/Wt
IdOLaITT9RJJ97jSTbHv+AQ+R2pVcosMksJl+/AGt9aVWHpQM2UkmWKQWBx31M24
KET0VLjn5wAXxaBxRPNZQsmWC/vWlH0br/aqOwLziMgbX7pKxCb1kRoGkyX6TgUH
WFtYuE9BduYKPneZXlDS2gsScV3VqymGFAm/NQYwUlvtVn0BrcVo8KqXxK3e3jnc
MBvtuEbmnl1YzDrQLtLPJbj7qMcLKQlqTen7V4cQZqmwoSeUvMLBM8qqTCjelp5f
WTSxrDdDFafmKsV9LYiqAG/qiQCdW826hBhVeuGRe5EzuPQI1YvlG8pP4FH1//Fx
0QVgRklBM/L3GgHMc6X7Jvym3rWLaW+7kLFz0z+0fzwpjeV409d8fkaern1bNTHM
JxSaP7BfwkP2B9JI+DzAvK8SPI6l0ehd5y2vUpJ6GlC0eZhQ82ZvyaMcvFfsbMRw
yEXh9QDSklmRzkK1qiEI5CGm070/M5r1DxwYU+Xvj7qg3EnU9j1L0wxxKdM6FDXF
YeMa+CgsmKmxwGEiu6CtuYbeRT6SHeWmHyvrdBlapbv97HEspUtWjlZg/G8Ruxk8
swOTu+sQ68m+qUy3v1YyKwszuSYs9u+XwQQM8gkU115653XFaZEWMStUbSSmbyty
kKDIy289PSB7Ir0lgmI+I0L11pLBaD+RsNhvv5VVyDe1vTyn64gBOPnGHVEeyO1n
6qPq2jDH5y7P0NoTGx9HicqA2xKgxc+FWVEc5n3RX48bgvX96hRHPiY+Su3dYVPY
x3xiKNzs0iqBJyHnzP8sTK+cAEjvoAlJUkH9mn3l0CT0Ha5AaeZsqkLQClvcTo9t
un+pvDHhFOfyOpo1zCr2tyW7tzdSKV4+G+ZLuR6NJRmYyZKvtI8vp7FM2oHqdZSx
4A9OcvZG2U5YNMREZ+SOR9gRrTQF1kX+e74Mfvrc4t2bPXhdnbBUuCkWM0MhnJrA
uLX/Z0GptPqj2MGXlfGJinksYBNUT0eJ4XY2vfdTOoQ3H5TQTtCHVmQXyK8Y+IvI
+1fLCl6/NGLJogd+ipgOJP8+v6eyiuJagfmJXwqGhZNCr65sodYVpoUKlNhy0sQP
cW34en/gNTAec1RCot9Cnmfc+7f8+j/eFgL5Qp+Uwub+n+zJHBgGQaRYmA4Y/mrn
tZ2qZlwv5QUs0Lrs488520fViXCcA08BmlsOPlNXXOLui8DzecoxpwmOzGPJcqfD
RxghikEXjL7WN3S9zZvg1dRcAI7aERT9Rc6TsulmBH0/LnZqye4wCUPj8FwR1A2b
zL8x89fiiUqFlrH2li0mhXhNWx7hwxwaNBLi0h464M5kgGjJlTpYIrH83n5LOd8x
r252V8Y8OXF75b++VsvQ6ygU7rm/rfP0cNSw9pEzVpxNxxJ4JcD38nooP4SjxDrG
Gm+p8EYYWl9MZhkR3P36zHt9u786HTfANeqXAIlxG34buV3k/l3FNxwzgGIUtxr/
n+L2gSAnLl926tNq88H8Iqtdn+bvnzrDlZ9/bf5z2QAcuBcWGrc4+NdCZvycyN7q
F6wz3cCLkyXCtPCZwXC9hXa4wqN980HEzPb1nZYcLvO/qtcdQcEkfI/HW3N7Lbk6
78rG+cn1it+cdV3lFiEwA1h/g+z2/lZFKfGMLlLwyHon2hf2Pg0VAzjIFNvyBm9Y
DKBihlzMoVTcxS+99WXIlT6Gzf9bQP/7rks5CmGTQyHovrHWBAEOJBhyJWTriRPP
MaH0RFMSpxH5VzI/OS4JJ4Wn4UdnwrHDSFvNo2JG84XZyFxHroK/Ck5J+Wlw+5e6
AmqR2nFdD63po3xLzwg4h/tYBZGeYggHo6/Ak7L0qAIXpRfoGHb2GWN5P2Edfwh9
w1kMHbTtUQLAhA2jGB6C2g3yUD8nfolLVTpa7cChX3DTiR/QEL78w5naWuV+pjHR
8f+NKartQ7xTn+E/f4NLz455UQHaj+7y/34ipXQ9n53SwV6/KyEKB5VMOytyA7bA
mcPduCD3UEw4ZgrRfJVjMUVoUikv4sNt4y3LCvJ6nusm0a8S3jMzCixWrTR33/Xl
u61vtYMjvzQi6loZG300S2ihBbgQvNynAMnz3EVYVA00eiHPlAq9jvDxhAU+3hEE
yx36M83MaDbDNDqkUMzdKry1u3R917HsIU7k3ekACPCElk8Pyht8ZqOJankiv3bB
mAyvFuR5XFWCJVDZYgcPRz5rOHBYyvxgvFFxubfTOtKA+7sd1+T0QpZ8cl274Oi9
ZOECJugS1/0OAW+B6rujKeD6qb9Ckv/UhMozlIteCUAxp3g3sM4wBMfVZMgJVdZ2
XQDv0Fm2q6WEztGxgP+Faaqq5gkxuvw5Uk5YNE2W2q/OK29ScOCUudqqWj+ZGppr
Wp+ft4SICL1M4IExcT6ojLBoFkFAIhaVNduywHSNzlky6kxe3Wqx23q4QXiLL1wt
ESB2EJihe0MRTH/WN0INKqgT+1DSMXoLf4lLVVSpVmMRIojHLq34gDI31JQEBU4v
BvEXNDLmZxD7EY4rTAIrj7Lm7JCidzd9/JIkRPWUP9xxTvzi8gIpwMe+8oip3Eqt
2iRGh+jW5w2foaIH6UIo1pa/vImv8nUwuCEhLrFOG8Ks0tQ5zKMFCe41p8nOdqW4
bC7RxiKo8fCHjN/zNOp4nKxnxyYjQwiZlzv4L5LnDp8i2kd2+I50O0Dozztd1DI7
6UrqGLzGahNgUqau7gGpKL8KXTd1FHGO8uAhMJSOVDVbL5yRI/oCWm/TZIfcYWXJ
OQ7l8PdQ7eYBpt7Uqdz3Lb6vwRoer+NzpNv7BZrBoGOBLuYeS0paJtKqYOgurALu
t4I4Te0RF7pU/V85zCPvRHP1hwCbPllbZWPemQg3HCbI7S20t4xNiaPmmCO5fGEs
yR7tcjHJUSSo9Let+3HkQcfhesgxy1g2aU7mjdviXDHgqfg8Q6rAvD+mqdPXnChi
e7P/Okr2Ktuf5XoWopW/Cm/AbvG594qYdYqGdCZZKIjCJx0rnrtyDFDivzbhlp0u
xSaDeE7hOhcP4RLFC9mDo20jHuuh77+uAzRL5+6VxL9zd2UpJPoGgEnPtW6wq8Ef
/TaUySIWF1JUukpg22AW46bJZQLd+KXKjY7pO93NixmCmfWML18yBrS9UnEwJP5l
EPmRHEVv7U5EqENoQ5NUBKxobmRNCyVhMQIfXvtTpTG8iRluarjl2p9qpPDEwYcq
bzA0dU/ZfvdrKxFPC6AizJlkNl+siWdiOvpvs+K+dJsjbGEAXeYWIk8kV43OEbUx
Rm3TTIliVCdOr7FWQedzSSAvYvVv8POTc9xXJTJcCAKa9hOYioEm2bT/TOnFiSgf
En75enKM4rLgRnJCPpS0qYA7mRZH5jW7qzTHC/7kAofi47k9xeq5Ze97PHSPwIrU
9GwkHS3K2lMRZ5UOqaVHp8LvWaGkO5Yoy0ot4oYHXNuNUgvHQIZeO65qYjgGvGH8
iNon1JLwb2p+/anMeMCbl8O3ZG0qjnNHJI80NAkyPAsJdnXbt2eilrf7HE95V2VB
tjaWj6BdALGyaERXcuFpK5S0OJExrg1mbRH8owzKCEPCgo5KU2NNq0+4Sh0CVs4e
x62T8K1FVl1dAr7Oc0f5o7T7d9xtBkDX7nHxMiljsHondZtq2H46u1z8Wn037kzw
A/x8C703WFUVVdZpJneqTAkXPQrfAOQC1CQUluAYiTk8/ncjNZOq3UyGKmnBNQnK
+kkM7YfRwGFvJIxIr0VaxentEI7nTEPYwev8KWq7O/RFuoNPaXKYujor+Z1wY2cy
EEIrY6DcpGJT9RDzRX3apyPw/REw+61rMsT9MdIaIkNz1QHrq2W8mEBbEoK2CeJp
PDxQcIi9Qy4X6VGKdfoVfqodt9UNbhrW1kc//2Jj/eCkiBvIfijT9djiiwFw7rp3
SommMeCFujfVk5ot2DflWg==
`protect END_PROTECTED
