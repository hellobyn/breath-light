`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bk5d0RTU2nfwSI6DmpGX2tvNy47sn211IqEk1/tbtr+foWZaV9AM3+4av1Io7HU6
9w6pmBHBmSc9zgSQA4xT4eJAdlQKoKg0TAQ7GNhBDpvY6m1UK7Lg2l6bDmdpu298
7dyOva5DkoKT8nDZIeLbAShx2xTPnrIiBsn7VQ6Sp6u02p/z5U4egtGIi7MxdcIU
bskv3OaUGdZ7/LPA3C4nLMrQ8JrWDmgPOCk0IL/LPDUBZrxA7X2aEOqPmp1lp89/
o3iIViTHiRCKfA1TmFsXpkOj52kuSGThr3O+6EwCYeIV7FSARtTvcgWnM0h/hlBf
GdoKm0aVv8zNE7eZxlnUva9Fg3cRRUbuOZpJl9r14Md8LmsH4twxJ50OMf4hl10S
iwzXkWSh9jvkBzLN3QvF3wA8B72INPG3kCKm74z99t+XXvNYiQN6wXTQaxCx9BaQ
ZPeAvc0Gtmmo123y77WDUlhVj9U3akghDpyGMvGEubWL8nkxnvRgf7migiOB1/tC
U/zKbLNf9ib7EFivC21MNvidtaIGr/waBbF4b3yXPAMZ/Zy/2743/TaEUpJ7aZBU
2hgirs/E7B3AxkCLizrqq2D/5zTrDG25Q6AHvZSbp4YoCPiHgxHUp7ePVeSdOd4c
SD94Um/C+svbb7IVUUiuntjwcHBsmmGfGjv+DmOxOHSmwhlLUjGZKLeueE8cKsMH
bEOaMuixYxHrEmgSGxpSo1I/MxACII38mSdTarhZBY0/hdQXVehu6fJtO+jQ8eC5
8453bJrDohgsQMYta5COdqqCwuQ8QEawd9/8p6ZPmbyoDrodV3iXybR+Fyu4cqGw
7oAj06Z/H2FUA1POkTTMPIKLuCf++GLnLT0aYarDZ6PPayviC8ZK0mqJSN6xN6dW
wCjKRmGZoRDV9QGGta62MKRjuv4lcyit21skFewFUNnYH26CnYSIB80iiGLZq4gM
s5KIbo2ZIhb9BnjJmxBdwIXTOlC0xJjf6SDj3BdeYfsJTZSpp8IiBUkru2naoueg
JGh5hMBb1WcRZ5EBDvTlavw0BlG2m+x0HYW7MrGe6oeOAprQNvKBeoLb6P3DAPS6
GA86jRNC/dRzFIZz1UkykayIpHE+bprt14D1g5Ta1t4VA3YgEsap/y7rHQ0hULV3
CPg4k3Ilh3t3CnY+admIP2XM0wGReTVq09dgIVOZTAeinsbiy5ejE+YoQvFRrqiv
BDDVcZI0QPvDpIweGe6WXQhUGyExgNrL6s28I/1jgK2iwJjzcDu8QZv/oXGhEeRP
Er7kGSKOfTZseRz9BTjsLCDwt8hVzbrrkwYBHBA5cAD802zyHJoMm7vDyD8ljcuT
gHrPj4I9ojiCjicPTFGSyrhNLVeM7iZbldpBk1anux84SqXxfJDhOp4gWQdez+Pf
R+LMLpAGoyUX1V5Dw7YJbLKRJPZrE78B6jCK02BPVD/9kv1MFt3qhu18B0iXmT9K
m4H4ElXuhfNONXumBTf4KQ==
`protect END_PROTECTED
