`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0Am5WnaP1kNs2j4JZCIqo/Z4Dcs/JicUTH+Hd4Bx+6ufGUFBTcxO3U9GKwRm+bU
MLvPy/IlDfFwYfsno2WLLEk6fqLBbSK5tcdA+TInVUujTL9xAjX3g4zagwUnZU1/
VQA5XeWIiVPuXwJbN9Xcb6jZC3C+7uW6wUOnaev2tcflwh3fo0kww5vC06+5oDTR
s8nU4mTviWXy3Rms4tE3K3KeH+jWEDyAdmVc9wUHXWYW2dJG2Jqp+PPdJfhApahu
h5OjfhUasRnNw1isTxKjeNwWmj/7VxL8ARA9cf+bc3Ar780AkRAfvmNhqBJAHaMS
/woR1d1ZKiSYLht5Rr80QsLgQgrjQhrSEKb1USCNLyHxPVJtN+kor/Tdm8wYx1qw
6C8dDmbPURrShTMNkKhInNYYnC+6qBXNA27VrfFqY+Vhlf8QZmvurao5cvNB8H41
2ot4To8uRn32uT+Kq4deLjHoGkJhJ74B0yz8h5+/ml3hfgdFIPRXJqdZb1kP8+Oh
xLx+ZbBRXZOLbHhF9RX0/lanpkVEHMmz06PUSJX/25OZSkd2gIRJp7HLq+TWQPD6
Mj9+jfH6qDO1NYa1HHSyClZOb9q+Bj6mPwiGUzomFJAF7Z8MbwDt5Ouhyq1c0hA7
GoXRrb5M1N78j2pyX5xYvZmZsu8ITNnLkt3vWeuYB0cUcdYmWsCMrtS/Hlil4MZ8
kFRmr9DVJ+yvUIElqXkKrMfM7hDWZx5dU/BjNzWMWQalWup54WWTzCt/BfK/TI+Q
SOJfu9+48jw/bA2Nwqj+mC6IA2gjOr16xjV4v6dPzl3YPAOy4matYLDhhfQ/O45S
12c/gnXFw0GguFPGftw595OeOl17y639U5R6uiun98b/Uceky4ITjQVHIZyLqApg
SQHUk+KroSmyhJNeAVDe3ztzNsOeBId8wew5OfbKj2mFFmm+wwZwIsQWEEeQsT2U
mo3EIlkWys379VmZeuMC8lHebN/6pkNDCOQXxPziCLWk1NQknky5l1FAL/439bMo
qikci52bdmOKMRoZwWjGrNRAGTNVPNjt8E9VSDtKuYmWwVlhds/nOwR1WInGuoLX
kitxgKklpGEy/7KWaJrjTnTD0ed3iLPaPTOX2dcSrh4w9x2i4hWVFVtvvjzLBENz
wMgOzjHNzZeus+ypueCnscWDH2/VGN1zLrmV0lgNVhh7/XH8e7qyGXPMRrOL91jD
ZubRa6rMITT4QMEaCwlvPufPGBrUigbCrENvAsSf8QSA46HvXxiHefpSgJTy+2+d
HK9+6Dgpe2KtL3JIq+eZi5x/SCiQr1ptJBhb0FqFuNc0c88owgnb4loruIutzWxW
qsxuCQxKfE1KCIvQbIZOmzNP6kXP1llcJrXqJlDjEes2JHt30Sasl0QKT9JVEoBF
YuthHpwW3BiAAnegUqLv7daCjXyEICkyBKXJPtmDmIvq9XL7K2q9Ov/Y/6skN25K
tI3lLn/Kojr8TfziaHgSfEwE2xd+dLGno6ceVZHrMfa0Q89VUpHFodHCU29CXu4A
/i7xb8cJvMkE5Od+AeJ0tO04awz+/sm47u9/fYX/hc4vb1buhEfxp+/dVo6pXyym
9NcnURFsdAKUHj97kYSIstKZjLO4NLKkpB9iP0nKI7imXCJ1bFLuaK+EtfYAvEoP
DHVcVWx+iT/cPMYNOsohi8dhXZDrHcuaEGD5ScbdoQRNgjcYILH+81i+v5855Cng
KogOdRSjcKNdcdLqOGZA3iX0zKiibxu7Toxg9DnKvWt4gD4C7CySALPyNPLmpdtQ
vx1DU6pppfU9M5nVx0Iq2xslmbtLpJplI3jse+btzC1L/Ao/XZkmpqAkQZ8dfF3B
pzJbi9a3NYYaKs6W+2fAqIM7xfMwBviOlbxyvAspLPeABjpgAPuNpe9I4ymTUiBR
Ajf/Q8OncotzL8ucij0+kjbO9jKY4YJ4pj0zdB0/wCZry5p2i4M4pdfKnhjfKvwz
nMK45WBxI1FwNjl+Pxu+s+T+YHaqCwLyWkUSFw6aC4c7z+E1yZkiaYdAhLu8JtLX
gBKoeefC+3ojFjgqXNTqYRKwoMkfIECowAQBP05vXiWWtfJ4wx+gH5VmzBxexqkk
ONq7Tio4EmPdb3Se4gQF4zFoEYdbUClro22gsCVWq/yWmAGE59fpA2w3iS330GNv
jYhNEpmpn3+5jiynkq6dy/2IQAISWLd+Vx0hbb5W0+85/XvSV+I9UrC1HCTdCN3g
KJsuLsaVQB2X1iDnBblxFzo8i9Yr6AYCBwNhsqkWy8c7TBC+pBbW4Va6spTpuGeo
Pgil0+QtMjtN7vB5+8qg4au6Jlwz3NDKdFn+UiDO+ZlrXsxQK8xCklZvbBu6J3uK
`protect END_PROTECTED
