`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TymdR/lWwH11fnigyNX5FkOSd3HglS/77OKC9DBKfjlEa14J4u0uIe1M/BG3R5GA
YpNJRiTpfPeT7wMz4+OHK+FVapPk3IMhhezU55g02XwG5kuzNWjCq0C2jBCc1OC/
ulaqln9v8lJ5rGIco9c5uRgGp1Ylx7jg8b3HOoD+sQTkj++/yG9/ktqkEMqvv15O
iFBwk6JFh6GTbdrMMZvxNs0GZu8JFUjBZuiLvn7YsycURlCrI8ek1Bqx1ergpyZN
afFkOXxkWG8SafRUdq3iMwBKBqdsKfUX63I22hkn03Z0Liky2O2it4M9FV9/zY4a
fGKl1MYAeQ9JTGorag6fyo6/4hoodhNjoQHEX6pu9x2t1tJths80DFiDT7V9Kmud
fPg/Wf0ULdh1Jy8lHT0oQxod4yz6YBk1c5qKBJhXsjb74Oo9V40mL7zM/UAFx3w/
OAkaDUvbPIJuZPwJPtrWfuf9rwCKD4X4lIsUG12eWMxz2BLyaK4uvmsbkdQdrA0w
8w4uOc3iaMypQvauTnOCqmak1QO1S97ywHqCGBerdFwkXe2Sa551w4VU6CPKGOCS
8dYXkOo1G5+LCOVVjeDTg4KS0QnhXarPTFSV7Z+yj8/cNFEZRTpff9QSepc5O1Rg
2lcDNhZM8XhVlc0c3X3ZRIfO+qAmF3KmhsvF4gwO4Axuv9eE+yjtsB6x1/RaYBJc
bEvZFdaqWxcEHjyXI1TioSnqnpcLrzMFiyjuXWP6CKzPDb/XcdUP5T4yZ7M51baJ
5j/lnFVhfaAJNJvRV9oFMu6EYxmFc9qFFPtsvbbu6rkUSxapA75tYo90CNlxMR8A
Dj46+SVPr+piiUhNE7E6OzBL8WbdAqhN7tAG7sS0niwLaWXvOQPuyob9KCzmrms4
A2g9/nCO+/8lAwO+tbFKb4pAAKHhsrIIUomfeVfv/qWr6LPMxAqEibRkP/+Ys33L
yVYHLVFxPZWIT3YAIe/fBgVo7XCl7zQVfUybbBNvH2UQPQ+uZ5sV4n3QfAdTW/Ax
4wNOSVmobWaMVr9lH9cU3xg9+kNP9RKL6QE55g3BjbU=
`protect END_PROTECTED
