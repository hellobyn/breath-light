`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97ZKmbf4aO0CLlwXAkjQunL5F+mU4MNyoXa/IxNpee2qewawcpKTfd6fcCB4JQ1a
Qxu3M7MrDcbLflIhIEDublGL9rCYtnt8mWDYKMP0PMlt3RUNycmkbWlq99oC6vdW
FEZGiw/XKgO7y1htLm9PmwpBayKZRdYjtUo/LSe07FQCD0hLKOvbHTum7QROYgJe
kWTy9LV1vevld4pUmHLo1DXSNjB2ka4T5G07dgh3b9ajiIMz/KRArPgQWtu7bOqJ
mhRjcJ53nZYhIgSFBY2qZRgOiLFuYAKHUP0ZGj1gfa281P27tKcQbPYtfcgwiJZh
aN1hQBRYlBrYvXdi2MVsVlkhEq8g05ey/2N0z8Ojkx7sc8DyNRvD1k7Kvih2sdfh
AUtaULPvqU2TFEOQRQeUQ8ln57qAobXb5qFnLYbdF2uK/kEK5rNsEf7je24TgZXb
NWcamJTOP2Fm+PFHoO1UMTqmGqHXRKPgjmYdN+Vck/UHtuQQSze4719bGUiNQTu6
7jWa+RdO6aRogJb+IdCKeRfi81MfXqqMXV1YztIAzure5XxFJ8lVVfcsZ5zFBkQ/
TsjlHcNSXlxMxNxrl5j/99EqZQFSS/YydFlKtoKtvvsMRc0xrvPgwjend8oUcSKQ
HgFtrYIEuJ2ERYY0SNhNoZKLiVjtu7GrXSos16tUpMA2C9I0xFOU6JIyFMcPgnZ4
s/COygFCLzhQqzaK5ujE4qBGUSHTOiOsKLxG5BuL5KSrK4piLcWa0mdSzNPISMvW
xGDqFtpBEvq0J6mhPQDHjKQJDP3/mR+xezMBVLQJskrg4PpCGr4HlPa00GXvAF4b
RQGPGh4G2Gaqrg+8HXrfRSoUttk0tZiY4+dtGpono8HgIkot0szx3SShyFSILcJY
VcYf/BHnLLqbdy1YM1F0GjeRrg5gd4kzu0OC+nv9Ttk4pNZ1jnP2K+U8AaGAtZtI
FmeYH7k2+BYEnlp2RG7nmIlBdptAv6T/cOIKebs9jaZ2vqf8XOWGbE9PjmzAFNSd
P7/jxqv7YprJ+hsCVA8YsfuEqSM9d5C0v9kM0T8ZIg4BIXz2KGDJ9yiIf31K4grv
fmcluyF3/7JT9/uMcsLanxEFCADyn9XYu278yc4AX3zIitPqcdjwgZ/XkW4mG985
6NWtg+iXhSNP8Frk2Tg82pa/a0H/tj2oFaBN4mbzRViCW+4Xre+WS1EhqLx/zWM7
NAYXMU129mC1lsp7C8v5LQqNyHYt+ku1VqPy5hC5R9CvpXPzmafnU+zK0s7g8BfR
eXfo8TCeymDxl6PhtrKkZVpPPT3vB0yD8qZkUFarOF9X225IR/ogGtrYdzM7OZ8i
i2v4Br60rTRXXc7/kukiUHK0HI+XjHR37jMz88jhz8L7PXvx9gIXTQgnbqFEsGpe
6erlji2kw1Yl0KDlNxIlWosGMHoP9C71zXYmGImCSfm+7yIS3eBqIl3C8T5VE3xm
/H6Zw8qW7AO1P3e8B+vQQwoFo00IoK7fb3CtXIS47PEzepE0IYsDlIDPyuvXW42X
ai7InGgYktR+6u/IGVUmM5P7/A+hT0W0VM7C6YON+jzZ9nNjGFMEEjBcKunYhuQP
nQ3NP5f9Ilb0tUqqbbJNoxepo1s/I00UQiCAhI3rQ6ua5wamW9QWZCViikWwMNKg
3OxjfKjiCQAs6q+j2p3iANmOGXk+wA7r50AbuxOgahJ6k+tY7s3hNy5guTUFUaXM
T+RzRR3+pcW3EHCjDJ1DWCsqhHcpx5vNSb6+uWLrWVb6X2FTklZ7oWIAZtDINmk3
mjOJKAYj1y7v5YgoBMF870XfDYmWKQsTo6Bz+BMhlfU+oUKw3jhMtVgNyDgpi4BJ
W1Od6Ju0iOpf+cTr7URGE9U3LI1IJTjly+JLzbAzglln2woCYXsBYqdY/O95q5yG
iU6PwAXonOlcDAs8gC4dazkBlFQFNcwvqyhJkG+SmEx5Uvy7pyXvjZUKL8p3mAUQ
KjEla0dwIrS0kKYxl5g58gt0C9B+4rgG8IRqEHGUgRsGc9T5nv26ErJgXk+poz9E
7L5gs1U8WWIzTS3KtN6V2VXaUEL41IxJCK5CX2bVjmbKOL776EwpR3fRRGgcuXUo
6Am494mpch778G6v4IvgdaSvLojVxU5Nvs0Q/zXRmS0igQ242VvQtn/5Yj5mtOS0
U2e8aP6+il0iiAi4UdU3+2AGJqppARbGTjffpM8oVd6P92xGRjgxU/WwuDKQBc0a
vPjzeckzpp3DfNexZIpqBdbEQ/gGSEKa7q5u9Z97AfBjT4jY2PXnbZ07eSLXY1Xl
FREe8dBl4gvKH404sE/z19OoMVhHUGRBxEThFpQA1FgFH6JLPeqZelevUDW1u2U6
uQy2mHtWUaztpr9fNTDDothPPqiquEsFILCAdMEDsCI7d34X9HF8J9BSwcoNbtLi
cIoLna000VfJj4yeld++zQ1SA4um6PZ5/kMEDiOWPiNcp/J7Hu4Pd0YJREQgH8wd
YJ3yKetHy+REUfgDnCaVICBFtha3QyzBxymF3uemKIMR3Zyy7sHP0LKV4D1o7VKL
E7RPlmDmy5RebKOKMGCm5HSf6K/4lzof2ZNaTXR1u86XaN55RwjnRM0zoGC+uo1b
oHR7DFgkPWjO/qrrjOqtpqWLtIhB593w2fdSSpyVltpd1P5WCMLV4rft0vrO9FaC
ZFea/AP+ctDVncsu7VJ38ULmB1k9ucJIPSo40uzmOzFTk8itIfcGMG6qw93B6koM
nRe0p6T3AgGPLNHIycCUFusU83WWBZmHKhKRzhxWXnDnXe87wneQT6Obslm9LaQX
4UtN0DcVrqMqwzNSEaVrAJoKtuyBNZvd42ePKPNjCBQZppZditNB8YpKzbEiV2ZA
3t1HWriXgDXBruin2wYEJE2HtGqB14AQ8eO18cnRNGdnJqI7Yc+mdKepqpCFukdX
L7mrHNRsJfvS1rkAnVB0eaKb7QwPZtBwSx3IOSiUiDLTFj4oCgvPcATgh41HywAb
5XB24xbLV7h63Rhbuy3qd5S8kPhKmeovDhHozevaryRwWbGxzz4/KC9x6sOaZIFl
ELShi/56H+3R2s600WOZ44obDgbWtHBgf4mKw3v4MA0HMoiZSpXBIJan8Z7QIaDG
AeR2lVHIf2Uh1Qz/crZhvZ95A7M5DPzMCII2XVySeFKuTAO2EIW0O/2wis+cLi8K
u7kMqMik5jjcPShZYaHd/GsshDWFgEK5zvF5XpG1T678JntcjlFGfbXuXlMPdGVV
u6CPFojaVcWlxk0P9P11Mm+mn2mKDeSpEoir5g/lg20/ojh3cM6zDhjrFgNxG4zN
n8MSOAv9FI1dQxWEiszfsIWWZpt7TzHb3ldlITysXgKDgXV+CgF8xmH3KO/ToLcC
wJTRF4L6vsXJJmBzxSYvfs8weDgvGDMYfVOPyC459QlQKU/5QIszhtgdEbc/S8LG
QKdGihrLrR2GzZ9d6RbKXkkMMotdcWTR1h1+8uThJQm8x6Yy0azst15aAGzrimwP
BDeOTFVtyP3600sxVb1MBIzeDZyBJAq+ZCXKWaVuT2c4tcE3en3qolcgW0Tr4Xix
1F2eZ05WxPT2cjoJQgsuccY8I9JhuByo6jR+LMzBI6Tc8XaMcQ2Q0KbEMzKZaMJu
hZI2rZHZv879MAgU1tkepdsVXk3W9KamQ7Vxn4ryKk1J6O2oBFq5zA3xEWJMpo+z
4lYtvSNrRLMl3Ao8Uu6/nof4kMhSpj5yHK72XMuDeNps4MGcrJKkf9YV8cwDLu/x
Lx7A6YMTG7XGbd0bJPp1Nd2KOU+EgM7pkEMO2ffNLf+zKOjnrJviZy4a5MIaTSiw
BzhNrKI51PiVaSDZTL2Ak5XWdzGuflAlLSYRYMUijXPN51iALfWG7RggRr27lw8c
UJ7nXFetUOhyq9rF6pzXrg80UaJLYRpFTHgr0jgfrJLuiRb490yFlaQEfXaIk3aU
r1x3PuGSvMSXDi1enCyHN6Bdafnj8Y5DGI5tPr+BMpA7b4D43ssffYA0Okj7j5yd
2mgJH5TW5+O7TTdURzpSa4Gewwo7B2ffQVPOgbf5QFANqIPXKKz1QI5xLw3TY9pP
tDWbdE63lHytITyq6V9qWT4oOQEf6gYwJODAfImK9i7qGNtPqyXGvXKyQcI1wDa2
cM0sXkOXVQfgYmobEKX3FJ9TYRsklHYFgyXt3O/+HIHuvVbG0gUeg8qm2YqEI1O7
uK9ivckb3iylgEoEm8xtR7AK/PHty9jBPQjaEE3GbAtB21erA7FtwrH4foFMmxXX
aq7Rz7ysSyCA4BYk4vhjL35jce38ElrU6/rFtwD4YeFEhn+u+FGy3OX6QpgIV2ki
qepaaagEgCgUaEWT77c5gG/XAecBl6dEzbAE85XMaVclLbb5TciYO5wBCZgLqs7n
EsJUNilWgwTkUl27Wf3Hl++guPGwoLhsEf+h0ciUcLEKfYkW6P3qdgHukM7YPjAy
zmdTr9rNj2aJqhGc/TfH2EWKfd9fQKvItUw6Q2IH0XfZvdUidXO2MCY3RM2pAfGt
oQHf+ltzelJmZxgcxzRZztH4eIG8zMirfBeCwB5qEs4sTDWdPSMDxAMUsJjy6Ohm
7ftd9av2zSwnK61z3JbkRiAWiHjn7gwrlZ6kwE/utm9k6vT2zyNal+EJgJf40SFf
dM3B2CdlwP51pi8GcTzZ1o/RAKG4vh9FWNDMVbuK1FmM50bHkSPW6+ll+l7wfFLK
4Ys2j2loN/vkF5bwPmRZXPfjuou/WommYeyyLOqG9FZ9ci+AMndI+1rmaM2CYTQ4
U+cNrgyju9lLBQWXrwwXfS17RTLyWdQ+z/NhR7/nEaDm1+0WVo2FpnV8uEQm/KoC
Bmz4bdngCdVawBwXmyMnxlRWckeJ0ivGzXIu+i1qnH6AV3SuZRWDDQ0vK1leTwIf
03XYhiTbbMo0/y2UuI7IgkjWasXj13R3voPWvAMu13Ub9K+gB96wybKXg1ckiwpY
0e4qJS8+mQeXy0PMiI8YI17LpBaPndJ7KLPr7XmQZ42u8J+i31KeH96HYmZEttXf
CTzBY+pxhhGZwJPAOI7Su1Olv9AfH+sKkEWOIpdRErM1l6N0LkZ+lxP52VNh8zwC
IvM3oBtinXWSJGEN4eAWykKHOWQ68HRWp/fE+IW8x1MLGN0nYH2LcUHYvoCxMVgn
2tHApZrIQQbEbogLDQPGAguRO50soW8uO6uebJdbkoKQbGnncmTL1jpMAqR+tmF1
81V/jbnTjHpQAGRt+iQwpASUqx3bNrCPQDf7emFxqD2WN+huS/sOUNJCasZXO9Lv
dixOOPNzYmRQE9xtVs2MFyApjby3yP3Ar863W5ORJ6OGAxH8hEkUM9BuqrXwa1VS
OTGm14ZhNdUBacUuBv/8fweZ26uUTS1MhCMSAlsbdgslUjJhilptOlBfRNRN1P+u
Vjefvcvw220QzwwD7Fzgf8ydoYPIue4YgDF6rD7HgJaavmYgc9uG8qYiJBpgGZuE
wwq77A0FOdFd0ef+Yo8plfaVWJsLi348PlEMKC+CImvwSp4dgxDGR5c63dT9Ap9D
OkeDaW5JECgnQYN0KhmFK6Y7pGvl9Fy0FjNlstMk9R4bWxEFnvhXO4EeNqkDqWT3
beZynTxe3QAGRnvEsb5kS7s5QY/D1xcaMm0SiCLuXrm5R5n9HfkpIDd7AJxy1PDx
uzKXJ0a3pGc0JBYlebS2vILUjw6bzfWEZ+2n8g7xhOUuCKXNd0FabcD1ksntC65Y
n0ujB+ezLQizeZAyzjWZPkpr1bZ2N0X1fga+Vq/vNf/l0eAP+C9yRx9m5eyzLkhB
fOkg41yjVR7rz2aRMQeh6kDykyNJtSEgtRiYlb6rrrEACq+Ge5eRK1meeCI5zqHt
s4N48PIvG8nKczv4tjBi+IquXxkT6hA2r7SJbY4wZvFQ4BDkQwpDumtb9xmE5XeY
varbleNUCDDyZIJbRp6gQ0YZhin6na07x9KmrZUdPLICeoCvLuUcjHnMvxGHjVOX
1auCLZpZYN+JgR00osijm1pNjcNHmRpWsiwjCiAbaWecTmiA9UQl47UTmN4Bi7QP
zSlt1cblSk3hTJAsY6rv7LkVKSuCov3udQHejefyG13TjgJyZJzGsITDrv1qjBGb
s6OhklCr/OAm7CR3UDwBXm3M+7YE283SfVml+4YmR+owo+3m3YIVzrxGxeVwLnzc
p4G3RZpPrP2SMznkDCx6JCA6DbceRS3OBAabuc9xc70Zd//Ev7/zvKZ6uT8dROk+
4D7ijy/D3KqHJUisoKyFYOMWfUCPkfOu9jQmKmKLjNYe5YdeYXucV/SLK+DNkwXQ
TGXrGZjcE+egcqlFb4ck5H028VbOGVYJBU11Y03/UJkbcaxWEQFL2vbtEpDUTicR
PxxeccoHZa46T7CE714Zj/5AfoH5xLKL1zkFwWuwFr5h8D8iceZ+Wr2UF43/iBhi
lCTvzSNzZ/0sBBEF87t7jcoefmfBwOsPGL+cmuqqsyQr8+S1+rKL05IuKuHsE7Tt
1lwU37Nx85w4EvqOoC4yLQvYr+tXpTnRZuN23WSaVL2GX9xBE9rSwyIF78fcqLP/
c83TEqURZvsaNFVWUGFNdbv3OlSbHzLt588tgBgUeP3DM9NlExHcv4ol+NEH5wk8
5ws4e7vuz7RrRfFyZRTG0wmdgAYz5XClvWxxM0mF/tbdBnCb/8nzAZ5sHIupxim7
evPCRPFmnkTW4jTC7eW9KrDrZQxlU5bBRXzNBGndzxkyyn/no9eSd3CmYh485H+U
bRUV8CULQcAgaEPFaNjUHLE+z5tBeJ+Uroilv5tJAfLptGvyfI9DO9HK+Sa7nbxx
QkcZjGtmPe7upGsYZ4Eq+8IuGbywcgDiUXt0cLg3W4VvG/bmQaq3EeqKqlrYczqd
jiiguwUhk44lrS4ya3/FSEUzNxAFC3pLEm+HBfFNT57Eno5sXTdB2npHcrqxtYD0
halIfLVCURPP0Np5i0UcpnA91GRqf+y0SwD4XQEVvaZJPgNnC6bQ2cRH2Cqvzp8k
JOqODPkDmrJ3MeGYVwl3ZR2kOQ5UiAfFTtkZj6O0/+JyDYWo7i/8xRpttFm7TdJM
U1TKssLQ2SSDF1gAyK+cJNPCeEbcjSUDWQz36IkkoYuxzAMtxLnd0/yoEPuczaBP
YP9sgbtLmlKTIiLTyh2yF11MezJ6hHUNROMK1recxUibM/wa/oxmWqjnN3Dhzcaj
otJMFsBcxX8y5YAcTKmpoK+XGjUGcXui0qJMf+aMU2cadCHiyt/MzDWuKPzFP0OU
glw3BU4UsKmGXK0s5HkClkXIL3RS8e5afQi/+y/X/ifwD3Ftv2FHIXJ9+HgYmsbp
Q+3Z8WXz0jHWIxq58AbLNzIhpcKYgnFKhJlPVGJVBbntbtaNcB57Ov2G9pcI0MAx
FqGk6gF3cHOVBsoyynHAWt23ozYzb2aRQAcgymiICJvqQAEEtAJhOxISknUg4ZAj
/dmzb0TqW3BrurG/OH6iYxbw3tpxLw9MCtA8i6CrY3h5R0dQfSikVbrAXXPi4SlL
I+f1ASzVOflRCjt2wgrvPrcyi54+NCp74cIvq3i0HgrH8PRK9Vnd69fgeQchIwHK
nwEtF5UUkqbv6HRTeNtI9qxyM8Z7pZ+b/6WIz8U2OIYOKbMPYQmsm6/MD4DEvpr9
71XvzUHgRHxmggLdIOm+YLNnP8xQumeCeJ6IUT41FYYQCT9M8r8UAW71DDeOjoOu
68mTRM8btK6DvteWoceKeYv+qExYt9NxdOlaHxCG0hGksg/zbihbJDaXDvIEiCnU
MdH6HTzhDhZN3q/ikDr4tWDA60PeN3NAv1PpIR9U5Ln0EtC+Q5Atkq6BLr9MLOpP
+eRtZh4GOpYS6VkG24x4IFIu9Oua6OLMKPU1OXKtn5zWpBs+Std/E4E6NsD0rtHc
70IERD/ou69XPC/FLxpjmQZlaVY6KhX/zXxvYIC50//FYZ8BbQl8nz6VWOa0E/Ni
oc3VVThO4loR8svKglAHYuDaIPpG2Cyy4neuYoDWDuL7BUzVhZ17g6rlV1djErL9
IimU2wkoLdDkJYVYcuQu1r7cuMLl1vvIThHmeoOWYuxVp5Sf136F4VZYpeheDhqS
EWXX7HRCutfxs3cvx/TMgeiLLkf3Zv5SbRrNMjG+e2dlP1eRk5KeI6dPRB71oaGs
b5PiWJ5C16r612FEVpMWdi2wR4iD8NPdnFnSwUptcAFTQ7TTOgLKRJv3ecE91OSh
aewwzznctDcgiocxj4GKeCgS1oFsRjufgaCgeOVF4R3G2IfrGDqbc1lfoXet9o14
9cYwusTAx9Clyd4/QXoRS9T7+GVIHlSh0L5AjU58b638wBvHCkQwiggkzzfMtpXQ
CmHjyk2xztRxHWeYnQccBTfp2eKHLqCa8XAFfatnqze/0UeiMvQxLn0AxU37f1UZ
hCVvrz9bbztWj/6hAFpuFEqIWxpXvuiAWM/uShTkfFXXpnyQeVGdG25GcPraV0ew
P8GYl80/cJQOBfwciZ5kMeXRrb4paSez6ENiCtEK46BR6X34vRURPWY045TSlO1Y
kCgfwN+IttcASIlXspdbWrzcwmXKf1vlnk0dMZ7XqHUXjIGeZxfWjXkXHOMKI8sJ
7LOET8IbMcQdl8yDvQIiydap+QutnfMXqR/aoWXU1vXKAQXep6IRjqtc4+OY4F4g
LMboe0flfEVUTOXjoqdq7GlteIIYnvmFGKdBZmU8Dpnpe4T0hIv8SwMpg+yjZto7
L0bwo8cVKi6aFw3Tb5gCHy9JVW5Dve4Ip2P7eKXned0d3hIX63qJvLUCk8dQbpQR
Gj6Rl0R4gi76ClZ7u0ZrQENTkOQfLRk3mrSKWAtYQan3tv6H0mdKtV5sZcjaBMKc
P9j6ycAFjq6v0CI6Xp5rlvkMkVAMEfWxrIepiuVAp1SkXY45trqzSYHT2aIONx46
HM0PlYY0MbiALREs5n2VsMyQtcr0fHGtTt5VSGDOCrC2e164ffJPlqcHJ6tLQ/py
Vt7Fafhurlo23gumGjRNaoovM3KSKhWieu3uh8z5iHDXX4/CIFu/BKgDmzOYHG29
VNKwdzZriX61WFUR9oJoGIrMLCqYIKgyaJQpfE04sSnQoLc/gyzv8SS/Yn9UCxDi
9zMnqnqJEcMEFmM+mVvmD5MIV5H4tLDTncCI6VQ8Rjficko5IPeKjRfIKlMCRSca
cdh2Ejo3WofHn4YGx1Jue2SthobNYQO6nV/brJ5hx615A4wHPi7qnra5oMAH/k4z
j0o0pwdhRyAeNQ+/EffAJGLeolIQWj+0SVsxjxAvfMKIqtJK2kSMMZedhXnWrj0A
iMhhNQw6xPFFmrqisO8OFff8RxWUDbmoXxZ+N9COl23ODZR6kk9CDvPl4Q3U3yzD
grE/LNWDZD5lER1wLU7Fnq/pbChhJ0RLIkb5TtGpTPRGrdtpSFF/RqX1vyaQ0TtQ
D52BP7nd3bg9opNnCI6JbbhhJ/px8BWXnCZaS5jqZc5uPWgQZDPfkeo+qYjtTVk1
4PQI/bO5NDwcxubU0gMtWeYZ3n9WrybEf5ysZn5L6MDoBnyqc5l0fGL/FCAEcDJt
Nme8gyJcV5CmPHXJY1U5PkbiM/KX4IAJG+RExxgYH66/8yLf3V7h1nn4Qe0bXY4L
ko2cZCqsMi7c8SCYG2fy7KiZwgr+LGMwEfMt/uEMF5CoUY7pWnPT1//VKAvEVBqd
ygB7mXK9zXpebiSJgRUJ2+WlWHk/Yhk5DN4pAah71rQLY3uUFpktp+hqHCJ1BkeE
bTvlhY82YarBFxcDMGWT1rzavTI2To6AdIZmGOZ2K57yyr4t4lKYWt39MXG9FYb4
JgpofCITPNE5CK4ZqrzuaLvfJg0LFR7mjGlDXEmeBNJXtE0Ija3r6c7zyvESUi1l
dfeMv+EeBpnk9fUVRUsiRkPIO3pHcAUeJdMeIIy7sn/vVz8PHoObr+ccS/O9mube
ySeswM1tPqctUH+TMbrJdHFPhNkco2cIL25sVA9edVuT5q0INHcgiGppADRlFthJ
jgykBDBkHynRdcNlXqPGWD/wgTv6JcpMItJUZA1oUaD2nbdFdhkAZLoUQGn10SFi
BULHBi2B5Q2EJ586aeoSyOeA4w1RRhMnh5FFFf9WecFf4J44t8I2u4o1i0X+AfN6
Adf23JqulpP08uWN9qI8rV/FPtuIASBGJIHqglfPn/pt20wjdJ+aORI/qSAfn79M
2VgTFgXtj4ZfeP/1CpD7c4f7tUdlyQNk9Jp91Xy42pLzvSsk/VjRGTMfa1T/CTcw
7BR+Zy6uaGK6l+3VNWhDySLFOd2RB49EAMEGXgUFmybXkpg55QuwqSoXEED13eDk
MPgAZO7w+3JkjNr/rSYmLptpNc+sX781q+akT5AtOx1GlhYTt1TxASodu+ZZlwww
44VOBYS/BFKORNDp/4EWkj+Bt5UZdDiuhkXRp49lvUtJJhcNxEIBu/GhVGh7uhxN
gXbhLnS4jZh8cVFg8l/ZwX0zu8uXdKUGwl5folJCyqrF4qXP/D1tei5vUeSGQhVJ
46Sbg4saaPNt9cL45KLopP9pNh6HMr9JpusRMXuovQnV494WrdrD2rVlwbPWE+1b
CzClsPTbh5i5GQ8WvM6t8VKnw3Kk3g3KOgzEb9jJfrFHIUCqStCztcH6B4PqxA00
yX6UBHHaTUat7610j1uMbQAH9J7Fs5Al5zIMjk5MtHWPxzb07EB1HmC7AR9pCmEZ
2HKwuv6R43jR07+s1wGMlCYpzyt2g/E1p8OV8Wz2P2PrzTZ7PAtjdRZf5U9w0kBk
ffmwxZh84s5DtXLBSvvdvQ0r/L5F8jj0ryG4P/PgK31Eqy+FAAsXtsewQkQs+48u
BURMncT0VjjX4V1/WBG5a59II20fBuCMioAmoz32fqg79wsPJzcsO2vg+wRpEZ1n
UN27XxjKalBHpRm7adxBOpePg/kBUKOQWDX4yfxj/PkPihXt5467SZMGgn7j5yDG
tTppj0W7Oczckch78234xRXFDC56eJZjHsS4ekBBTyv7WmeNhkPpSUMMpD50gCNQ
tqnN+PVHa2Ro5hMdLv2eAoIWWL3wIvph/BiZPpVXUroxklb5qtiUQ62JpBkNmadM
PgYlPJf9yWpzSld8KazGj8KoPUupcuKwNA/E8Rv7A3c1qWTUK2fLLeHc+pgs0lf+
nvXTFRh/wTqjucbok/SEgfTYIyiQoETvPBgsQpFVuoHn2tBtxrQ23f8Ts7edptV/
qq3KPGRNV59jLqOR0RLAM1+BsTCgzei8Tf/PAS4ITeNaPTVGcTNSCmAbLCDTCDrH
aMA9Yzoze97v6N7X53kQXRSGi/V7lR9KwdRcOv4GuEEzHKkS/WufXjufLab9HqMZ
WXGv+cZDZJ207ALrNz0K1rvmf+vlRsaLXffe++1KTYxBQN9TRzXJADwoxIGcdrsh
oLJ04mkNHrTeIvb1FO5tmZjvC2mcFLluCbu+fdCuCEVttwGtF8joVNj6yJQBhlOb
DLl3Z+FuAFbKpJRcnXqduzxX8F2GpriONozy+P4SwtJ3oR3fJD0V61wr2Sbvp8GF
fjuGhBTU+kJgDDu3PTFURAKQHENjfQdZn+pkbPxmh2CiZuOjstMo5Botm5sxLhga
hSA3FfwgHic2dwDZZoGs3ut27JoXgmbIbv47Gd58fVfwSkOuUpOvuZOBIjhCkadT
r/dA27IOUHW0USbLDqclgS8Jkg5Vsw63vqpMPwve+SoLgb/0fG92WzYsPP4qYTG4
d2ZNwYADd47PWYEEms/eHYYRiq9IcRAz7sQLDArWLxkAlTvvLIz/Ia1jCN9dBMIg
JSAw+LXlQKZy/TjrtIz5sCfPu19mE5ryHn0aNiOm+S3aeb44+j5n6Xk8xDZDlIaR
w2UTOo+bHpWEbkRb3zkuY4ebLvkzt1wYq18zuvSgRYnqw5jC4UDT5hkjQtJYsL9/
aV0yUbvd4lrQmYvbamtjKxBRYIl7o/vcgrcTEMabPMPSIwVmBpmdcDX2QkU//48X
GlfJQnfCmw0Wf/2iEz79w14BUqG/+dk+aDBL7ixgLdKZYJzBooKTL57KsjZjE0wr
SPQHLa7GYYRP4d1lT8p78yk4Lzl6l1pj5XlbBb1mX/rVTPottcZ4LQLyeqpbhvnJ
HShas5sDWS1XiQ3+rXA0DY/ekrXoRTY89wojuCaElelWfyt6nulsUZ7onKlIho/P
xU8DzBmAmcW5eMgez2/F0yAViUoA0P9yswDzjiFjBFd+gOtzn6+OgABg0JuA/5jJ
SxvoOzBiZ7+RaPGPCXYCdjxZjDATTt2bWiyQ1Cph9a6d3a61XUna270JXc3hJ7Q/
x7UVuWGzkKvRH3PkmoOfZZ/UFtDp/6L2f+PPVN3hgXwSBFnrRGxw9d06bjZQIzOz
CuZGF018nl9KKskVnXrank8uQtxSQ6YD/geir4RYJ3Gvb4wEhbDFhwTGkyEmmkEq
YuTsxVNRpArpeiPZhiQxpkj0a73klYZmzVXMT7Ih/oQEOPz4xzSrDRFZ26cbseJ0
Wk4ReEj1f417QNi2vPPdpajRPikkBP26NcZ9dcnaO5zeXVDWmz9kzMUakN13wzma
xkMIT6R480phKh7rSxD0iy4h2hr+whmgABxBcBqsQdOWouzmnaSymN2OkEBIGB9t
sMTP1pz98yUC2fdwoZPxi3IVWG4iGRMR/HzfkFsmHBm9X1bXIvF/rIKSvoHO7xas
d5+0wBiZu0mhYmCd3xKbY947txg124QQ9GflnftQ5rinQlG1Ww3OZKC0t1LzbBI9
zT/c/TZNfkFydQ6SPorr1SRkcLCPFQ3bB5qLxmFKU8NFOF+dv5U5VqmtptjlDcNR
lz3UQcBCix528tl9+gbqBIaq0ilkv0e3t0lebIE6r4idiOunFKrepZIXhsPzr1G3
MtBrnkWhML24tQkRZUP6XHARmaa1UNRoOyfzmGuY7oGmjDx66cfpwzb4FlHVqc+D
FZXEQHpx7LO3H+zhWURa10Mxk6Zsua0DNKeRQCBdB5G+2dAkeReqKGiZRAB+Hvsn
av0Mm5u+ys9OYPAfugGb9cX6zGU/WlFFikqDZREuTyDr+XTYOfEEQlq4DMehvD5w
oN0hr0dlb9pUgRH/khZq6WBmc0KKABOAPMqOJLOxklCx+Eya+Y16nZ05eDzVC7VI
LcZtKeEttT0emZHUcqkLO/Vwcc4oEf3lujAdaoUCWZP0KAXwmABvTaZlstN+rt64
MMXOvCwoOy1GhH3Rq4yx2+IwbOjcOOZF22BIxq6uWGM=
`protect END_PROTECTED
