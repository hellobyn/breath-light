`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WfyFZsMv13fynKQv5fOWF6p9ySsawdOIqO7GmkTtJkP9hDrNqJAHfyB563sq01He
gLZuvcO/gC5HDNzv3FFJx0zc6HxS4ecPMBdeUed3qdm/LcSGbvVAwp0waoTz2THQ
7NMfD/Eei/fyCSLbdIQ8aY8xmTuBoOMVKt1VqBR7zCxYtr3HrUnclWXXIseUJQWo
yughK3H0BEDz1kCKfrlaSAMyRdmSNvgvY+68Z8MHbzWWKLutl/JRCdDHnDvjv5sQ
FqmT8aLqCdnmyZaI0Ot3CZmLTnYSoGABn2/GBp1Ww6UR6K8O6ozsRP8kGc1e8vBX
IvKOd7uM3RRNKork/qWzHWvi0Muquiq5ONmTpQDDc6wJJVxyU23Vnf7+yHjYIGOC
Tf37K9g5r2+qAXzz0fQ6VFD+8rIwSFRaCzD17mIBOS7h96YVzdPEMM19TMfR1RtQ
kcmHJxc9pTrsPfte53lUN7PXTrbMe4VHBlNGiri9Q4vgznCPRoqV8ncay25GD/dy
vaJzu6oW8+5sE6BqlLTioJBWmbRNyWZz7n9mAUAmljyuOLkdK//pEGKchSvyyvvY
8LYqTXIMDwESsZ4VSybYujhnrr/0NqMBM19d3rCVQXd6/bKEaSruBrfhqVAgBKG1
ycvQMckOR1CpHFrOV/ZUzlW6NRb6VqF2Xm4Ka7/vvhADhSyE9omsLj76oxdPBuq/
mIhMFwvPkbyxAUYxaLT5tLTEXuruw00nfUzYlpHU1FnSVuHF8m9XTpBmHvTeQhRO
51jhsO3mU8IaxKeDOYlG0j3NmkTOV8zxm9WeUp2EX5Dqd2Z1Sl69yzhQOJqV8C+Y
mOkgMQ0jMmkWOTSf2cfRDdjBZ1Ywp+OdVfEWPbBD+9FdNRTXoP7e4vsb/VthKjt9
x3IQ+OujHk9r3/n/8ILuejG4DcFTq+JK3oAwQClIPQDkvcS8xWI8twlEj4EX8EgC
4lgZ1aD14NWJr6mZmASwpujRP41SQaX5YNydEFtGFlrsqVLEIaEyFT42yRBvinYu
eNxRzS3QUAVxGhPZ0ueYEoXPM4elqi0OLNMnaKIvDzDKU23XcX3eYRvJGRqfXpns
mnkjVGHDWIizFVoRtpxGcdsyOiLRKi7GUQrJeVkoiKTtwgZbW7o+tgjklOh21v/4
crnO+R6AFZ0W0ahAgsw8rI4q4pt0qPwKBHoJJbkYRUBE2ei2O8AFlPoiE70p+WFD
0r4/yMDdm+RpEL3J6V0YasFuackTNefNmpokEqmHzyv/35AFuyFI+5/kIP10pIMJ
dGHJBIbpHiL/sS12ziXvpGzH0+CDrqjgWmNvTW2fPnj/fgRzvR8XmNx1nZVAfapV
rNjwDUbWfEDd86OpRtuHXmC2WJO3M5OG8/JfNQiFBoVE/HWR0fuoSp9DzaaR1xQ7
rLkmv8tmSWRovHkKWfkbVa2oEkH5A19z8EiPUcR48g7CTPsvKKJ3QgOXOcDhfFgi
YRd8/YUCrV8ziNJUTDdKEYS1AP2Uwr0BRM51saX1rw2SEyDnk+H0ouU/bsKj5FPr
59OOOXE9VrQmD5kox8R/JOqB5tKYZjlgESqHsTY2KF/d8ojYQMRd/+6Vb+eXM/Ry
TvO4LKkeZ+RMR1Y46Y3DqyrWpRdTe7ocSbZApwTNLWMvakD9TLZcKHY2MaEYPuar
d7CnqKZjrFaRsVNncobv0VBi/19TgNdSSic+JLZ1Y+Dd9IPsjzEZZyJRYx6APFYP
hasrNMPCBdY9Yam9mhZbvyyD5Jvzc0RpBHxozSRuyZS7dr0uG0D64MCy0hhp9gbv
4f0vIAc+w9XSlnjHQNrsb7b9hnEuAptWkofdR87/DK1u8VAiTrH/OZh93M94Ify0
FCxhANfIn4UGBS4vu6cJXbQfiA/bSTeQXgg/jO8b1wo6Df5pLGk12L9IbCFJq47u
RpIbEvJoNoBwb4vs2N8YjjZDQZQVELj4/JAK1Ztc5Xa3D4+0gq9XHW9ctBPaLgDN
g+lDj5u3Qs0v15XB5/NV+o2xhV2A6JgS2+gjMLL6WQTKhrY2DmfiWUHzpst7cmB/
pLz9SwZDECNLBQpL97zroEBgibENQ4uAiKhpSYmTMbocZO/L+vZxHZsmyBzi2mEE
rOvLjW/iHFnFVKeEZDNLkOUFy6AaOzs2v3ii2ekLPd2KZN26H1+ZXKqvxjuLYESo
iB2hEsy9txrccfbIdT3XyZO56c5Ko8jvVLwb08AFIuS18srHb4OlrGE2oDflt3bw
U7ixvwTmybsmGSSL8Vrq76WJq1vAMYoyw6WG2hqtVdUANu9hb0hGD8H+8542frvO
A8Ybed06S15jlm/wJByzfzaiicu02/vWC1AHDSE1c+j47i+y5LPuLcXA54CNooRn
yOHVZ6PnmIXRu0XN5X2O/easxTD48l9s0q1qHelEFdRzDpJ2dUJ8uHRh7Wniu9oQ
u555r/78U8moqRtPN8yOKiGgffZ8SrX9ZW1ZSoHS4tz78WEkTOMPh6L8+ecNsykm
ZZwD9O+AsNP1kn8zRI82r9pmgJK44o+JAUmO2WE/a3Ak2JvPitReX1QuuNQLrwH+
da5rvCHebTR75SwMGx+6oGD49Lj34nh1EKiDi5UjshRguVID5FjST6i2GHcrP4R2
Q/Vd2XRab86X8yRNj31ApyLucTVJAdFdxspcWcGZYqgfNFtkcvN5oe01rZSAHiuh
tZsYaN0k+Eut3XGEMRL47az8frB3+Laagk2rud702gMxIWa++5VJqcraw6Q8qkCB
o77nojfQt4XNv7t3WJnZBFRAcRBGfc5E4AXiJaj6tIcOjgJocrrX74QL++nlU//T
xyw6ng7OQYt3mcAN9rZbMUY2ekU43ywDGXYhYVM3WWzqZYEeLaeEMluf3eftV/MM
sqLWfrDp2J8mQ26FH8hCqsyS0971YuKMhsSYC17HaKYJorc4RtMV41RW3deNlW+D
G6NG7zUwwao64fDzXz/b39/PyBLY36dIABvdm7x3FpwA3iW6Pm7336VLA5+VnH0H
z6Ynh1f45Muiz/+5A1zhMwGs0qEnbU5O74/FjCCDUuxMmnHl/cGVf3aitIWtt5Nn
6yoqE9+/PkjepmQWjg8zT4pxQ+orc4WQ18bxa3MF2BIPi4rDGdIxoGREMBJORAkA
UcIkZv4KzqRtcpqZ/otwbh9VlBL9AFq9uqZuLNIlDwxkvFIrdZEcE1gIqWL7wwDW
u5W5oepd9zsmTp2/8tqOe5lW2ocn1i9nY/vRxr7EOJ3Tcn8BaMv4Sk40hDWo72rM
Lp9CM50haschNa+tJT9521pYFYbCrNuqkBQMiC4TbCb+5qd3dCtAaKWIpRib5uHZ
wGjQYg9zuZUIowtG5BFu4ss1kkgG3fGWTZEM0Qd7T+NceLCL3L0BGaMQ+OeksCN1
Jmvpz/b4HtUYIjuUxinBD38xv2N6zVeyoDJHuDZEdmLuG5PAffG5gqWQMVt3iKy8
lGVb2N80ODgUGbxGgKx4fKQikNkHeiniPpO4Rm58N5OoGOacSTzWeiiqtxGikmgT
iBbye4t0iWPLzlwnfcx0HC6mWO2xCx/5a2AUUIdez3whYvKATzBIbApXF/FMhU23
5Xd/Gc6l8wmxs12tTeBmF2L4fgX7M8ldDH3F9vc/FAyhAM+rOEOZGncSGSyT1maQ
u72lEvnAcGkYp4Vid7M3dD4AojGV0GRuZVxsORNiO8oynKcyitaXUk0F0m4H6N+L
o3wFnJvOL6NaLxe5S92oF+YfMWPCWrGsRMbq6GA1a99GPekL/vEKNPHMVCnvP9E9
fG5PD9cqPdxaIqkJHTy5qln9zp74cZfqjlkDOjZ3S02BWziYXDWv/bAtTxBNqYiD
VFLr+C/X6vzBf/pFuJSwNQ9ZZgsvHUUGzU1yf2glyDMS3uLD/n9NUNxWvfjVE0KV
h8KYb40E0tVpj3nE1ZeBB+2eZkrmTYVVHtyqj4lHK3DJU/6LjRWLJix4bDB/GPbq
2m7YowLvECapwEPvs8896xjgVwBMIzpyKah0eFj3den0ZHaBUhrikuaAlOcCu6OJ
IZwxzSQzn1woEGZiKuN//BepvXy/KkLLwuEg5u4/VSXheRK0PhjW3FXETjdopJuJ
Kodr0S4Y3L0qm7QfZgl1dyVRLUH5LJYxEIPxo3bzzUMATjL3MjKsQAFKx81lwCUL
RXOiiK97+44GUi/8p4sMnxfukrLQMbc9ynhPoHysaNygJFGMDLP0UThJeL05snpi
2MrtvxFlvZBMOm7/YxKPR1wDDcfTySMRFw0yHgaB6F8yrQBhxt9P6d3gDoarV2lL
/0kAC20qeAce40nzxPpliYr2P0Bts4nuwwOOhbR/7m+rpNudYAlHIWw0FQ48MbK7
5ZkWIiW1rneBSZ1L6TE6TKgjresTi1KZGDsRH8ZejxZEW+8+ns8ACjPUPvJa41X6
hn8zdA8KpenW1DK0ij9QJ/YnwujdANzcsrpSiNRBb7UmMuX7eX5JdZwoitFOxxu9
b0YhwHng0/tINYDVtH+EXNReEWVzi1hQcqTHmjwcsVT8kchvuVOa77RxoHLHmnLH
m6aW9+tUUiv2SUAi426QzNF7ATtzycxeUYlcMXccKLLFG5BFiOodVqV3/wfysGY/
g605YaOLH/FqB97b9d/v77p2BvrmcFuvPl0Lmgrtw9ZdoR/4VtaibRUf8Y9NVBkZ
kKpHDVopUdnDGahXavaEoHiGKgNcZQPvVxtKMPTz4AEmD0wikpymAkYbM5MhGPcz
NyNxVNZt23FlcXLoGV6noXFTkOE+uUN1qYlTx9CN1vSkagefdmYc+iIYUPKPOitm
8MD4MtllTKXcv/04AU6cKZN5pMMdLSF8Eip2wxLOm/kQYFip28mMfVKddE+J4hTY
MKA63g6j2OXv0qBttB1P5eS/rVQbbsVPx6exatu3fB+WsZnJOWPNMSzdZONoB7TT
bYfbV59/watZFJKMLER6rlZtJ/4sCSGZdL7PzzPoORDKzHVi6RcEhKLkaxDv2XOR
ZZhSmdxR8S+nqkliDGzVNk4Ls/R85IdIhhuBSwa2NypB7qtyThZwzzj1J0ZqpR6u
jRXm9lScm1E+b+M190oa0PrQIOBETPgFyLc1LZ++8m7Fzcqw/j7CiTxeOjtejjhw
QaXQLPA4PqUU4TUzvK9MqEFM0WNYuBfLBwJ/TjS56bs3jT8exjl/wppL6XhXAo+n
flVQSTfI/TKDltkHKtMIBMbc+G0F8vXHBvOj8z+RIeo9IY872abcHy7ESf9p+CWL
cg1doiEmGc6n4v7knCSIsyE7BiudIKinWsIB6Ct8coO2pXYH0zW7nt9Rf1PtH+Uw
TBA6ueX9PK9R4WbJXGr5XJZeLtybO8WBoaMApveU5FJiI+EgBpe6LKTbzszzmJ/Y
vaO9GJtPUHqL+3d9MNymRl47lQbC2i4cA+ipA6jK5B2v2SAUV0cP2UmSZuqg/2RF
0vbw3xXo2CyIlUWzY6vCS/Dhf0+d2z34acbxg2N+8rz2yDYzYvca3RBL36R0DVP0
LVbK8/KfeSeTgeZWKQLn11G4sYEqYPgVSB14LLYCu8GxOjY5WG3cN/CKxL1K1QFg
cfgttO4Xye/uZhvsUJRS7Zr/rjMOc3IPzKoI0a8eCrgu6O3+b8AhB1vgksfX4UfH
hqT1zOO08nMPdBHUctuXEx179+Ql9opP55KzfOdRXw8JB6aEmR6p1nNMW6mOq3hx
8Yckx0XXxmNdxU/qKc/4r/qGJS8O94WinO3hv21HrlJrLSbUbTlvd/IRlP3vD76o
A8GWFn8YL3j3dvlBFxWT8hp3AZp9rJ03WqJaCoPRo2Hk+W4Lo1r7SzUwuOG+ODbZ
iDvDlUDnDFgDPAazQ3iu4KZ++85vP7/u8ZgdsVa/HHWDn94oyiQANFs9Iqo6QMN3
sBVvSeN59FURPdgl3yicMwFfo9Rnsz5NJaqUl/zjcAmPTYXJIuKZP70INTSNI6Cf
1HvuA/htxw/Ok+JVmv0NvH+btaf2DNhwP0NYJjUtEAmY6AiYLCfa0P7FEK5Bow9t
ut8Sx0D3wBe+gYwy0YzvgHPx7rVaCezbCKdT30NtZ5Yu54U0T3LibSeZj5RRdKRU
R58JNBs+jJeuI5U/FFVmh/6z/ou2cLcugXwJ+E9VCAvp4Wmsw1alHga2fyAsQu5c
sIRdHYsbYwoUe5M+2Xqs7imQHwHfsmOQwBsWd+ucY0H/azv4wTQ+zu+ir+tP0Nnx
gEvTOsbaQJP0LQdFoxTij9/U4vSMeUv4pkoEdR+NtcxboDZ6YTzw7j5leN9ZYS0X
LbOcAsYijxWu7Z4c+fI3SlZCB1iPDniblB+w8R/04CRqf2AiALsxvNn2tIG+hSaY
XC5DBMVxbljHIgFk9tNsyuK3zc2s9G1ZcX2plkYKca+8EKWX9E6WTkA6+L22wMBO
/+bXE0BTUxEPbHvLjtAnr53lkBBjamGiq7XS+MtqRN02qBMb7Qirf6fwPTvzWzAj
3rtzn7y+2BKQoriMz0SpbzcNVsT4EHvW1CA4xs1Y+SaZRmdXfQoPyiPPNrmujLQ6
Iv4uIRiBgNaqyb9wTgSRaX0B0m1h/Tq16fBXyQlHTfFEdYeuyeRtFDSnZKsj1INZ
M0AUDCbfASEtZvBrkIlxMF65HJdQybXN49XLznMu/xbR3M4cE5TiVL/mIzhEy91n
T1vm7XiSP7ahRarvdjysLhM7KmI5HdJmo2JREBVdVTzTFaFRVrdBU+mQpVEA7wMb
NxtJeyc4YpjxGeXkGtLOI4IE6aOBNKgsELUceaKzk0vT0yba3iQQ87+V74rypf6F
SkNnSCxKSvvOn8rOlnSAtuglHD7eB/CLgiUj+SoaDCCDgZXWJKPIoEaZv73u6wZv
mfcOxq7e1BvrTpX0j1sPWtLOGOKOZ/jnKn3nyVdvRA+iFR2dYc5N3B54Ztbzut+q
gHuaWg95XhCcG4b0lT6V6HqR9bvH40s4jPZ6AE5QBzjbnfPa2EtrVIJoLNrlbMsl
s/80APrS71hugL3WyA+Fqxxu/hB6TH3jo/nV68i3WkAVnYPnVS4z3x5/IrcFQH5n
WrnCLE7uTUNPZzkfOf0WzB/xEWOEJnOYw403uFem87+a2ZRyka7WXODUYXbV/Vz8
Bhu+CHjg6k6tb2vvy8xai/gSjQPJNTZ8AuyotY+/vy865nfeFdWnMpNqCqbG8rkV
xtMg7Svp+3nsmmKShsQlF2HRMWBdKw+ueBx2CR5oOoIYQU3v9Bsvevovi0+Vx1fS
RdtmRwPp1kegX9Y7iy5qg8wa0qfparkxgwGK5Q4AR6wZMhlYDazA6t8WTbksbgQN
KXOmZsmQ/EEk05sUjO2Ppb889mnFxg3eiTbihgWhB7pNh408YytT+RaMCozwwenI
Ti92jvfqn1Ly6MuXTKcvjY74enP44kvOKwIs28djCpeRMHaJZwzjRRqpKyShcNYK
QiInvI2tGff0t7Bm01ZmFF28kXzMun8Ts6evqh9skneJnYm0qRKiNQADGYhnBux+
C/2Z7U81pWVhb60roku+OeMm5hPzfiJURQHwlh/zkq5g2kYrRWwkQUQCIlhcA/NH
DtcTcNIZZoz2Yibm/vbp9WJBER/QFrFey9iyaSPtSohleocE278tcWnzveB6wgCN
TmMYcFVdBIelncHjHSmY+J+qBfYN6zxGsU2eIxyBlfgnlZz8cXAVkwvmXEtbs22c
qYxie6nTJrHJKNngz62a/TAFuQPuCGM4mL1yZMEmZ79C0m8b/NNkk5ne/v00jpx0
lT5xUmYJTz/Qlfp9FkAJmnpHAVKSzuKy7U33n1k/pmrZjD7/LGX7O236ulGEy0ty
DMaSBcJY9B/DYA1PwsdMsowwODrbYNQFPGGwVmQATqnntW+twp9Z46z6zJcEEW3F
+PMsN5rGYt7T7h+MDB/KvndRRdyzCCKsZW5x8vtrnEZXg2+vMyuTg37qT+phZyaV
oNu9XoJRS3iZw/h2CP1rGgNATIQER4KzhnfnQm8qfWYv1HyR7FBuskZeTeE22rnw
dlcsbpZm9xwVhNON4yKlgUcq4YkID6uZ4nSoIIFZUcDOsmbZ3hXQBlpMFSS0oowi
yafbZvUil/Z5P818KNkLgGdT/QmUQZXktrXzASCuIKNEkKs/Y6kNMiHlFl999GHF
Jzd/Z6bV+qRcwQ3Z6U+aBFM9tqCbbjiKH8BjYbLd21I=
`protect END_PROTECTED
