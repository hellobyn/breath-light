`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZSNmDKQOw+fP4ZPAy/sVz7zaaT3OTW9FFWUjOC21BYd6aCgTemJwNPQDedV5Uxa
N5NUGxxYmoJLJaX/f4z00QxTEjIDTygDG2Laeqblaqkg1GYS9qFxYSWmBdlYK6M+
BN43CtddUFdj1k6/GyjSoFkNJZDb36a8JpLgY4xch3RxKD9PX8w1eGFgDYQPKala
xP2LaRHQfPRM0sw816S5M2E0yfuZPxez54dK4uAlQJJP+P3lN+nncyc4GOnRg1M0
EpyMiSyQTDkX+aoXuQ+jW2zC5IB+lkVUG2f0yXn14iCkSeND5bJ+Q2HD77OTpurx
yDamCB6EmAQCCljHZ9zfasj8vi4JBE9O1AtoqpLPUy8lanVFrLB6/l8ctSLGs/f5
JjG9COJSwey+hGtWM92URdss7th9sIAdHyt6OBcp/PcpJ6Mm7mjVdbRuVocx4RGY
+K1fPevwkMmseGKehc6jYbeHKhR9ztOEy0Z41K6XUb0rLoJ4lU7BRZc22bs8ul/v
gnroq53QFyCZNIbEpHOpOwD0c62ynn5oiNbpiEtMOAcTwsTnODw2Ap3JBmOJ2+b5
AmsIiY6PDJoi8rIUcCgGOUEd+w1gYpI87oy3JIkOhfF+9gOvRLrlFnqCjle1JmQc
0doaLnOzVxvL0eRSodIB98XP8jF3gvH/hTQk4DZp8BTgnnXfDfQBQnM5zrw5FVdu
IDy19237FgNBK7KDOe2chjVo5a0pt8FcIn7LGaOwJnYdS+MPlW2bod2p4Wv7N/nr
f6050cEavb66skohwKV+VNwIWUoBqYxvhjbVfKkiei9Qj1YFPIbyLlEZ5c9d+J9j
`protect END_PROTECTED
