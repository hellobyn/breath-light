`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uy6o+LuMGvITFvRqhv3Dkn8UCFS/c56rMYY4rulZ7qYNhFeAh+HThdOhcPspaMZf
Nqv5R6yxBPJHZ6iXI7X0czuV2skN2yVDiIGN2wNFqYyRwRGWIwf3SCn0sykBMqAG
mG25KYXIFG33QU78la+37OPj891hWiHBn9Jj4IfuvPAdG9Dt+8ye8FjphwnrUtRB
YjUKvl40VHaeVqUsvt69cjNuvsjtAJ/iOVAkZ3vl7fRtjThOLv5SyvYkVB7xQb+h
emsxOQ92OXP8j0X3ZNT1kzA/ULXKIPeTfcmYB/v1K+EgSyqKpE7jd1buepm8vtEO
4/obGwdLXWkBgbQc/CF2mqkOTLNuq6Jd413rRiUXEff0pxdZ6XZUDEJjL2ypjOjJ
aZucuHOsky2JJu1Ld/UrcL78X+YdoWaU3R+kz/+kI6SU+uaZbCQMjesY7l0iK0DP
fU45CcY7wcYz8cbQBn128HIS2Ze2lAsyGZtT7UWE3nzxC9vlmf2bJjMq5SBG3MY9
eA+1xZBGPuho9b6DisTJqs+EdADCCXAfEM6An+5QmP4hmH3aAWLNqpdZjceRAqXH
OVKFbt+HSqAUv6pCNnpKnpXpl3WLphnZEXqQejsIZHcol+tdwRrAVv+kkZmn4sB+
tF82b9XOFyHG2PJFes9vm3SIGJTtr/dDHroYlZUFPgEEaOR5CP9rvH/AqM/yJo5O
Q//wsdCAUR61ZVMjPtz+2ufTMYjeu5614XAt/wZuX52cwGo/o/nzefWKVdmeAmhh
RgZtq6YpLQdtYITBhfWImwYNgI4JXnWGJ8jvuqMnGZbNbM8BXJm9zYu3yvbDmp4f
Niw3/xcw4eBurd6YwMaJdj65jrEbRwkxBb0xdpv2Cyegj6i9RBUN8CGUHGg5hvS6
myf44oGjH53mHjq8dk0ZrWg3FRl2Az38XPF7VbbzJp2eCUWBVTPmaIcPNyXhyRdX
BjTaF6NCVroxcUKdPAEz2M0RzL5VFl6mYDcFY1qgqb/zf5gTIGrUGBqJcZPJMaGc
h30+C+WJ0dn/itb/KcTaulzdNdFi9tkS2yJ7c2yZAvEuzVwY13FiLDhlTbezDmsG
KGldHy3Z0qv5wBzYASm7e0hruxSIjt0Dj9gpSPtMmvY5dOChGjpQYNw0WnTS71mZ
L7VqYslgkLF0v4BsPw+z2qAD+ZoQt3AOPAFQTcZp8HjcBHDBUO6kDLA62SQR7s3u
lilyT0mQlEKTdDvVMhxdgtZGtSG92z+Et0kMPU5PN//h5tB1I82+JKWm5Fv9rREV
NDCFEHpKwoE/YwIq5ccu5K0+HM7MhKgCndoagwDssDm9EA5tZgfNN3G2XkdTV/Kr
NZ/1KQshRF/zbx2TYtzAZHwZtNB0VmclUr80+PSLrudhmnNkqtIFiEUKuRIv65pC
H+9QYOWLaPIGu6/bhBGR9iHGfx6k8idc5G4wTksdUyetlglZnOu310Wz536+npMT
iM8mp6bHQ2uDY++3eU7o6lcAWkd8fh8+TDJCzrSN7SlLCFSXcpbwko47vc2HReA8
u8PfaY3Gg0eBP1ZiKy3fyyT1u8U7j8EgAkaI4hgoyJmLpAVpCGMhmKTU5DfLAfkX
WPMOM83ZIhIr9YgEk3yDN9Irj9FFIWHWu5wcxQ9HucXX0zgOFklRdfvQnyx3ea+u
TPJAkYwqpXxHhfikPP+blVeE7J/OErIcdRjoycrL1BbjxikRVtOoJpzZi7gWdqTS
XtlBeAEOg/OXFlpysVzJ5I7cGTBuruUxp+YY2skDzTC3z9E3Kn8XRZaUxdci4rob
lHCwxS7X9mKTW8mTs88UmRD1CeX65M/7kapWsgukWKi5t9pnLDr4SZqNU/bMx3sF
fS1nfVDRugVfRSsR+Jt1ad7FXCk1jLcdmfPcMhqFMdfRNZXv5gypfcRCKFl3PLJv
g1eTL+a2GNlrqBtinLp/isDxBXnowCN2XK6nQbj+cYlRBRKNxpIJnZ8GWRa5Qw1r
inw2Q3cFhZgh7zkf/AYGQxwyH+5WUVEpwJO1RyeL90mJ2ve08q13GbD9mdwcEiFS
bynfw/4GhHgfAukQXBnUYUioL38IHYeeLk9K1QmW8F2kdJEe7Y9CKmFyTConEYJq
HRmZ86x2Wsu/q8LEV/XULEa4nYC9L6ISpJKCTGQPJh5GoCLc2dmVB++EPpQ3i07o
5KxH7h2xYaN90euTyNBw0UNp4gPXQZa32l0UoNv0BrqhMDo+z3XfkUubtnkRhhNM
Xu2CznN81JOg8mfkmUFxrgXVUijmch5OCfwoOj5KSV337pz2WmmO//aLqHSSSuVq
KmCQGSMW9yn+UpOYxh/LHtGTPA7qFn/g5CthVMD9XdwgO2CsUK49vdXJl6AKZzhE
bqP1QDtKyHWhbMUIZULYqyUJry7bfw8Dasb7OY0b2oIow1sZe2Dj+8Rf7OWXxveY
YAExAam+yjfx1NUm3AGnmjZau4zIAF3dfgEdm6KKEBzygHZ/Ju2QpI0kdV8mYstM
Yp+uevINq/uZ6L0frE1tTgCpZhm8AK5ti+/QrjJKJhtLVEMkzDBO77V8osS+dTQy
sWYnMA5fmtkEMAwQO4ZbOaABib2rC8ZN93SQ33MHx5zUjB03Fk+LC9Tzabu0L+AC
fpq08zE0LcXX+uiEDrvUeBaeDG3kvZdwm/cLNo7u2Osz2r0QN+nZxTgEoSegBCl2
PWpEvwBOoj341/BXZwjCn6zmhT/ZoM5BAVtJnyJAJQOpwWtYhdrSQ1YV6MihLfKJ
GGGTH5vZDb9zZcfLnLq7rqDUppYARjyJ67WEdWCQNT/NB8zpZULweo3XCjH/Vt+/
CuAelBOa42iuWxosjx6gO2v9IUhcpiDDcRzJq/caEGBDkTIMW1vtSuBFRiFRY3NU
p4tr7n4uoNiZPEhEoHRisk+q1JXXVqkAVIxoX0xpZ7tjuqJUwa4NPWlV/BlFY5tr
FKIqAb2VgSj9uYX523J34Ovx21ATrNqCKbRZzQQG4qRS8wuTgAYa21Ym6dVoBXd5
pTNZqSp3GdzT2qOlfn0s+xCd/lKHyHvDXi+Ni7qtfre6TwLsIw6NEK+R41xwVYuo
fQXfeMUr62HTtiQ+OHh3iuDNK+JbMPAnpbA9efbXfT1p7D6znrgFZI6BjXMi5ukv
+G+VIHj/8oEGbvDpW/KxZJ52yHig8GZGoOVmtAxD/Z9ImCQLYyAlXJLjz/H5n8FP
PX0yxPIb7X/LtVCc42bIk+IGKpBEx2g5hXWttRc6IUrA4C9U2gLYOx+uIF3CyA8n
MTypyRKc1IE1gWUvA6Jiwierq73L/cVppL9cOVe9X/bk+rYvLpxWNCg9+ovS48Wb
SFayikUatoRzeduV9JdAzQDItVV40ktAch0lmZqRyqf9ZEKDizb5plQLFwyqKuCS
d4ODavteCSC+CnSieKoN8KgdrvLcFD8FqZXM679VxGcCxdZAQELpOuGPXFiiNJ6N
W5Fktr12FTS5yEVsxpohp9mOkAndqN1NkmRtYAX197jzX/BGXIdwsCsA+J9JDR4f
q1I12Q0qG1IOrWXkdfEZ0plVGX6vHT94e831qWum169nIkM1+pbyWZ4P43pWqVBa
ikFDVnXLjNH79c+EUyhv7Vl1IqTFAJV0pdFX4+7619C6c8PI45ETY/SfK2vmR6QH
BiQCPxBhXkvN/hfsYbY9HGpMbylyrbKwh6bYNqF2Aot5zLhijT5eVimV54F83d8r
gXv3IKfMlE9DVW9nbwWTjG74gRS0w0xO+FVoHz11UrieoQDtrZBWd4G5ewepr0jF
XzfibPTv+7OaW/cbGoFbXXkmC483iBDYXvTENjxGHwOBzfl3IK9UzvbpYn1FbF+k
IVRTU991xs/oo3TDu92zBpmfvwyeFphwteMR8pWNbetcz8xbsx/lc0Z61OcF39p1
rYnXeVPlruF0euGNzwERBlG4yntmDJM62OMhaLT1Lsvtu8TxS0mkjoy+hyT9cHLN
F1cWmhaCQiGO5oX3/9U9vnPQplNC+c/NAaIA8X9jAOOrbMZUOLUCSEv5K1rduf0u
rwSJmnQ70RxB1E0RoDyRjWkZGLH3Hu+aF9OylAJJTtibmduPhkZGA8i0IT+IR6xU
ag0oRtHOpaBYM4yOq7QAk6cRMcIUhmGjvAqc+H+NkVqknk9VN1fk9PwLNXp7XLsO
Lwqx/PftNjUVAeqP4Cw3yS8tNLTPvPnQdkdYbR5KJa0eEe3J9PxMzIHqAS2sop0a
bG73BmM/GpvsS3LBpMKqpowDonqSZ2lGnFZHzngEGI008RQuBX+q6PB86dP0JTrf
05CPFpHitJnsweedCelWzvnyTydT/sdUo3rcSRNRbKkC9Q25U0LLeSdtHmOuTct9
v6MW47BDRkHXLZYz/7hTbBDIcLv2Q2OApbdew9jvg2+JqQ9wfS5dcodKnTylVsoA
6fVT9gXS3s8C5CL4daiD76o6kQNkPOx87cIH43QnPhJnwA/Q0H7opiGNhjfVCzhF
`protect END_PROTECTED
