`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghqqORKtn6pHaDFvgKqn+Ler70T16eqyK9+7PyWd4DiOc2CpendMTxXHJKmZCIZ+
1K/LdburocbS3IcET2M9AfRx5HxPwKLtlNDVZJRBWAC66qKaNWMoLwrEigwivuch
VouXl2MsF+BtyYq+A9au+6H3hPHkwIuN4JrthOUjgE5M15SB8fjpUlxD9Jfbqiqr
RYRom6wMEMMQBplXfoV5Y1bVDgivs9cdUh53PV3FYO6mF2JV6YWwEU8eoqrEpmSc
eks6qDDfS2RqYPg9BqMFZqcReFW0Z5QIWsdCimrznvh2RAtiw9arBy79BzfviLnm
Ap2zP/0K09Xp039EhGHbh05+r/drAF1V2MNuRQJ0S5eigwTW5B/RnfDDEdcXop/P
HGQgn3YQd/KtqJdlgeUR1sSGuL2klSchYTGT9G/XxFhBs2SsuJTZa6+eVHMsiP2n
Bz2d2yBHVXeQ9BkAZqvmgPvCNs/tTFTr5rJJZy45un4IU+H2+2OHYKRGB6/g4QW5
kZs2HyHM6O/W7QNV4I2nUDziz3erWP1an6ZxpX4Ww7B3Gg7DrrjFDJbF60ev30q2
nTeHw9P0dypZgBNGNOFRh6sbQI/GBWmhlwhzj5QEXXD2+vDB5deptLVed4EHZIfg
Z/iM7f/mWimDjTBRuFGZnhdrOQA5czAbBpCTe/x8ZP/bcKkEhRjbZ8PGj1sN+EFN
k8Vs7itePMJoTuUizZAUSUV/RrI7Cv3UTTyQ+CvjJbrpaNprrweQMtulRzzd9OG4
TUGIwz5adVzImUtWi4uzDxoHpdLReR0TZ5dylx9YSZdSiOcJ2jm0GoWL74d5sMos
yPv95XhwuJ26iigDYLqtGW2f6zBB+FYRP6OSm5gBTIYyciyJbs+g7NOJwttO8m30
t3FL+wOdyZk9UMfCMjG4Hl13tXxFrjrgGpAlhSq2i6jltZ5n/tIcvfB5j1EF2i5E
7QYLqblC6Z7J7FFPsrqN5ge4t0kv9njg/7liZW3e3tVSNZt6gw0bDMYcwXu8snZB
bCfZWHoFQbRYzcEQ4awvtkgsOv5QFM4du85lbf56bzY4wRG8O/IWX8gJBhHJBSQE
qVEgGXsxQSI5xFM81Rpo7mrpiOpTS5Dr5uoqLV/O2fQx8ayZ3HgQS3IMPL0e+c6B
JD1JhuYXCIYg9a29JfZLIfN7K+EN1jczEtFRSftkrKH6kHXmOV0yDNxdKS39BkDL
+hvex5BjleGUe3pgsJuniwRsvhmmioC8ISMi1jhPDcIIuhLcfh0el141SiAkvw+g
T2INLytJnR+VMcR2LYfltCz8jnekGeDtRwgmIX0xqP6wTWIgD1fVIieTQW0x/uSW
EE6IgPr2ErM3IiWP+zoVSVq6kKHzrMrmVDjW2dyEhM/WCzwbqOJi30Cd3p1B8iES
8q9IVyHtnTZxxGViuciZrDOTceRljk4ozTLBCR79/o8L5X7mUL8WQqp2ujhBfF/c
O/h/tYo3PNLaivpTmzX4C+YnG3dMbZGI+TsIpnE/PhaRVylHh0O3/CNSeOyc3yzj
mp4f6qqqnP1O9i45RePhtih5a9pTnpWEhk75RDZk2islJC86jvVJ9wlBcfjCF7+b
+Xq/kDth59mzI4+g1fuNOg7hApHpZI8Pi2IoPkKiGNyd61FAqOe9oVgFudrvfkwd
X1Zy1qC63VQlGaJk9YMeZLE2PWSDIoZbgYcn2qPvcMKXHqhc1LqxwN5NTfmX3un0
QW9KI7BJt7CQOZpavX61Nl4tnYvKK+Jy5cUXXFzOvMZ4O/Zx/dRdoPgyOaSsq1Xt
e1j0l6SXYuM/taS/00/8Vs9hdf9HkvQ8Ktb0i32rc9htq0aEmFJrTVA+xCkcZmvD
3X4DHMKeICdRabEhqmtRyoZd5Oxqf+4s+LcySGTJKwV5+4nLtPf6lwy0Ksz8w+Y2
U6H08ac/l+G2+pbvB2+9RleRvCCxRGSq3LxHWz9a5TwNQtbLk+G0NdiWhvN1grtc
xL+Jztkx8MTy0nEiDi9uj2r6JjxyXtAVpryU7tt1pxD6Zx/eQPrHVh3A4DTz2ZRW
7oAZRDIyVdZDGG+fi2cwf43ZwyHYldCva2CVTB2ob+OMqeAc890PYZNv7h5zgXHf
bxOoJfG7opQdg2/7xye9FjED+jjLGCvXPeV0dB0neE2Y2tIcRdvg8zcZg8T1II7j
Wg4ltdmKH0Ykh+33Sm4POdAwHkCsu4WP0xC3wEx7mNSQP6777uS9xjKCPv6qPWMT
t6Zs12iT9g7E2uGx32Tjn9ZyMC46jwgkVD8h9G2FgZkOG9FXnNI92RAA8tZd4iNE
D+gHTV8vaqpM1mNNJ7pSONMFRDa4XtCjD//W4XMlHerX7vPEC1pFDpySf3cGiXaj
tL0jMPwqoRerPvykkV5vYuGUKI1O5zZuvgu96sJ1lNQJOZdqA7njyjoemJqMRqAa
ed9oLbaoe39s6ZkIZGo8XPR0bK7CoXnN1Ps4CJwXGzKqh2kACAPG5aGqWLHX8Lkg
4ncQBqeKW8npVq98ppJw1L9q1F5PY3Zl3m0HjcqhMv9vReawjsbszoZE800LvCzk
PVgu4hpZgekHtPShLAEJQNd6JZ5trqUBSPdRGbwnyjeysrgra4zcKRqqCSGTwjxd
hSaIa4M6elXKR44QeC+5EuJjKctYLbdOhmVN6JQ9klDXKTTZdCsIxkqeZYHS29bP
Rs30BJ4o32WZRezrhnMMbsZDFWNbul+KRC1r9FUb11oznvdNBGq26rH89BZWwAqC
3UsRS2CweBTDPNK2VrrIylPgafzrKAGu1xJvgRr5qe1wDmaYy2jGpkUKgAoEMjas
W3AFRx1hWIFABepP6UFR8BVWhEgsVRhO2hX0VG/LhMG9zbEWJp92pxq0+6rzf9iP
VixHU7/GXCtf9epVsOKLxvUrU97OePZbRPe8r+pG2NTlgA0Dzj52eWNPjHzcxEcW
DWNuu/aIEGHNvfAcSSTmUCOkMsSNdlqQZ/AkAejj0PNl4VPKCNwiKmAqqa3teZV9
gfb9tFu3zV55DqqIjyTHcxB+23wdXp2YEeRV2yBetRclIh1shlQafEQdiimiESGf
EFNRBaWRJe4Z0FlXnrhsg0ouZMw3o2/XVqoIkLtzH3bSBI/C7Q75KkY0oKpjgX5m
ZzCFm3rMqhPMk3jUQUYEn5+jx6KZmDx6586axVce0GDzRwVrdHW/lZ+7SUQiVNre
+14S8B6lFI07ZxAPjOkect+q2knWifpvzUL/dQF8IJ9+4cUFxBWKNTjnVIL4RApW
YG7y8SXUADkfyuy6ykYrII1ZnYJQElD4HdzEHpTQMk7zUbjqpJsfclGYUMIhAw7V
tfhxcdjyRExvgdQiKbokcihlohD2xaMthWs1CQoppeTcJTOlkYk4tEbB/UOGpGno
uSUDtfliGFVsmSfNXU4EEMiOwglWkeZsnbPIGU5mYV0LhZMg38J0ZglUx8RssYR9
HlR0jT3Ok3AZbJzLaS9DO25epvgX93CkI0vEDTQBqXIcDsVELFiMUvTWfgI1uqmQ
xX01ht8W6wvZj5Qr1J9s4tCA1OCokTxY5YwmJ3XoGm8DI98+9j3bokAAcHXlNVSn
hGtu4CNSKeRkiRkhGWUkNTckp3EYeUBoszCTcyvcUqR7lKOMmenpTaS+AjV30a4x
bvnvoIavd7H9foMmt6PDmNfYVcvHM6Gvz6JAJdHbjvv4YYuaZbOYOJpWFmvlI5Nb
f62SBzZGDECZ+pi1zqc6HZSdwFvMHHJgIQrYAKDMKpstXzM+LvXrQfiMNr7LNIG1
us7h1IYyzAVG/5EwjTSINdhfDyUUQAPH6Kv8DigKQn3I7TE+VBoaZgorFkyLkX5M
UISJxfZp2uubcOoPwzvxLZMgeXFy7xtbjcF/MSuL+X6JWtwVve+Jy+SIicgouOpm
DaKT6ZQnNac7tNtsJ+9VbYN5+jasZA5u+PqKN3eHcGDeUDTJs9Bq01hopOsG2Rvx
solECbNiFvyA7RVWNFG+pKBucQ0XkeAfH2Y53INaM90VdxQXljIOPQC1j6nM4gpa
kKVm/iyihbm2VP0Cvg/3PDEXw1lc/x1j0fygNOvxXpBTUgoJktuQPQi7+wA77nnM
h0SEU5p5RNZt5GsnpFWYh2gfTPU9QQinxAj6S+85uMmE2yLxo6U9h+rzsAB+Iwmt
VfM4saV0Y0+meQ2Czt6oSOcaRbNqfZGJ2U1cXccidEEqgg52lUMNoi5I8YKwCWSf
A7VaMsuZRebP4RRbyYKg46x4TqYTeWySfiVDDw/MjxSOjblfDXA8OD3SD19rk+wE
ZYsTtV5mulfxvI+qcGBLZkteAo9U//unGsLdBVBiFryoc42j6MyM+XW8FtQ5s0By
SADwu2ENnCdc3ONyCoqZdrW1HikxU9bR7ad36o1jiW1u6x6hCpiHz3wuHwUARHVm
FjUjtxPWLIQ3kIWVmypIAjb6OQlEmKGyq7q6Jpwq6Nlk9Jw8n6ve71WpiLW4kYyW
EJRBNdqd7XFnOjzvTQmpKcHGi0DQAH7mrGB8Zr8OTqSH4ALoDfxL8TpUPf6IvhHb
PXw6NVLc+mTCNSkPcEohfR4S8hO0V1qU1cQ5R3jZfJe3i6YcDe95ZlXwOAAojeAS
+1PQXw8Z+aeQeH36sl1dl4irF6+5rAFRGCHMgQkonC44Aqn40UAybdtYEOxd06GN
GAYr/Tjls2v7rT5CY3JubXyWz5cDf1SEKzQSehYIfeq/+vgzVe+KOsyF1Ay2Wbz0
vrMu7UZu7hicWgXFMN8phER6GvexR2RjI+IsP5dB7JbixusBoxFBREjT57Md71h+
IhVfe2daOS1RD9Gw6a+c/hlPL/+LoaP4s3oiLOIt4Aqv/URg37BpfVwRXA/huNOl
nyRL6Hf1NbZlwWwC4vgPvVbdghftnADKkv4+th6kLF30vFIT5WPkdq+4gIxckwl/
WUTm8wDv9PS9NF4LiD0Spq8wn4c+B5r/BFesnWsvaq0hizwEbuhBIxHEOnXYfz3x
A8xfEoK/A69Vd7taISkp7iT5gDXq/27ULA2naB2dX7i+PveRxdlFg6SVmeOGb/gS
hxeGKZ2ZSYljWhLSGxAynQ7qh0PE1bGSHqL64CjK0UD4eo1aKp4rsbmXL24IaA8t
llQBJIMfQc8K8FqIufWCjRMnGYUtznr7agsn3OQYajc+1IVr00RmeW9dG5N5sW3w
qEFiM35wM51Dcmr+oT8v2N6bhkll/+NgTZ7keAvoyI4yV0Ckmk5RJH1rZHNVfl4r
AS2lxrF/dUOxY/LygZ2Fd5veeyQvsImPMxee3TF+wfIQHbZgfgZ/tvZbFBBzs/jd
ydlb/1kU8Y4U1yQuX4c24NVaxCYC5wPlZR48LeKV4cB+6+rvWr57kQz57CxBnyxo
EvjGh5n1YafW+dncbNSgg1JmnOpaX3uY/muQTAHwGkP3wWDkGKmGkr88E1HYwGs5
KrRiNOO6WfVcb0RvEyZ9Nr7nq3kcB9rbolT5WGH6d6YmKp0+Ic3jYkqDkEVnbvCI
FTMTBmQCdmrNfLiC4RAaXH1OVAboVyJQWXZHj/L6r4r8xIrmQoP9zjmYkrbIaYxR
ZJ+JmCVgNTDBNnC6Dkl7TXJRHZSIu2dFcY2w34gch/R4ZGC5swy8Hfst4upEF1hM
Ux/oeCGCs4ArSyXVmtQ1WfeuiAx8m4XU/mZsEi9fKW3OPsNPBGKz/BOCvNjWdW5Q
lyS9t47u0r3/1jW1qA/lq0lunO8hlpcmcnyu9DT6jPy9+zUM+DUypcqsYq6LwMwK
t3Z99kinFutH+wEscxrNootuMRgv2v+RH1oBbfdAhPsicb3IVkGcTcGTePNR1jaO
m2oR9q52NHDLcxh1+Is7fiNdtrJvENl76SBwRCbAfjhhARRIzp6q6lIKigD9NMrM
7jaV/Di7c/vPRib5s7GtbpcI7FlJNiuGzsPXgIuehAf+NOAA19qT6cHfnxxvnGuw
Cywc3of3xeEXetmBlazlW1B7bRGsiNN+Hi+CNeqBpMXnTxw8dnmUmMeouUA5aYGH
lfA8lNlmiiCeO73vHZB/vJ+qq7Hc8rzrOUtpx67/ksBS4VGk6GsPWGwkqJeX5/4w
MJN7PYmab3S/UB62FxNgAfaYcowectVDIHW59M4cvt1iKMjTMK2SgAZ7VMlTJQbe
WMUzPBX1IbSJomLJtquMFO3U7wogmlW7oO+l4G9d8GJzN9U9S9azUk0xq2LkADUx
QVGZe1GVvFVOrAijjpmc1XL0HOfMXyM364Mh0Ljz6VHtoCdrbaKUZLcmsqfb51mw
6Ea0v8uC1zbbm6EGOJxEKR9RYbLodpmNSYRn0smjnW4MYo54xHYsCDD4asuk1XUH
r1PMGO7zWmq870gHsAWw0nGcCq9iaELPG+t762FZ4eXx3QDzncnZ6jTEAkUrQPnW
h+rkHL8iFAGHmTMFW2CSSoQty6BZyvgZxcZLANKBhttumItm0eWjOR8DQJ1CGwC/
Fo6iQMGALx8YTxnrihxXczKFleFnvuopJ3e179hA7w3LXhxDHci56XBZJ9Asfs17
X9dOJ6XbfZpIP0BawrRYLrp2MCExK7ggG0etP1oeevtpKoQq2lAcIEeT11W8Am8p
nfN8huHs9m+dQJG3aQ74sXOgYRwLJr1Emlqn24tV9G441lnFCGvIcci7uowjRkY8
nIQnJo36Z2HsLql7DmK6crPOX3SQR2okrwZBMstBZxWz3A/QpvbDhsLWTO0S2FM6
gdb5oDCOl8QGDLjfBAAfoNrXEbIhMH4oWlKHEoNKLZ3mrD9G+t+QruKjd/tePJWz
BbBlG1p4m8+NZTg7jknkXjVlcHPal28vO0p58QmQluAjnS1Qn0eQWdf/mACzCutE
905BDAXgPCIf6A/Pq0uIgFtBTgrIVnYjaJFPiLSGHPlhkKMt6Vx/NX09WSdNeoHh
q7wudmqbJuuchnnEX6lv0LRHwWB8uvM4manz5kyjm33dkm2F77zoRHJbxcPGC4PP
XknhXgIuAHlBXpNei/MbC3H5PoQ3fveDlQ0BZKi5OgMN1fIJKq8v7O+MSkvY7J8Z
oA5Fh7+ICC4RxEu4oYQXSjpITjihrituZI29OnCkVxeNcM10oo+rUSKHLRWZX7O2
fTaqDuqZoM/Vnc5KmUddxjs5Ym//IQzannf1DH8X1a4yH/Bad+wW0o/6hFZMYnB9
y+HJabIA1HRC8GRrEinxWwUYErdOW89LjjdRAF4f6CpxNQMq8FPgVz+nfJMA3JaX
uxk6DVZTKW3MWnNLzOcEx4FNkrw8oAVoqaw17uv0UQD0WpYQH7z2AsQaygw9HAia
kTr7KIk9sdTV1sNkoqbDNlRnbpyYGbJ8mkzeXRh6++s1hf02mdCzPW78pQlwaf+C
eRV0csR54Bkte8VQsk20OBqcEOlpPyr3Tb62yfjbuSbFcbj2PA45rfMja1NrcY4r
QtjjVeIerkcVvibs99+meXxDrsXee7Uh4dsKl9U6D3WD4F71ex7Knk+PWonT4iuS
E9rsVF5lVEoNe4V1Xxm/Menjnfh2DI9jQjQ/veWrkOne3IC63s6CN5k7uy8/Obuz
qaLMGKxqt2FKrcpEIOd4m4XZfQnVHdyf8xMqjfuuIEQExcxrm7TZQDzH3Z2MEmCt
KeKUlQ0JUd8yfjgF2sVQkyBN+Ia68NjKinfohakR5U3zx+cVYA2Baj/5f8PIN8oB
EH74JGa4SUyGyqzTSXfIWMyv4wN9U7W2AtwD5i3xjfxHsYmI+aVpIOsU7expebhP
AD6R/MUw3yav+MJSsWTe5D9pptwWa/8SjwF8R9MYOA5kDkkyFQyKbg0TbXXaqh1I
Yi65Q10cHSsAKXY3HmxxIAz4lVf2VJQ2CMpg/oXp4NRfk//+sL9QMno+FM09SOF0
G/iTXisKjvq57VemN4Bu68UT6aDI3jr5MebTZ9p913lDUOcHCKAzCkeSoRJMN242
Uh5EEFsY2DM0CU+xRR/wpGJSwxk/882hc1jQVpp+WvrD4IHieJJNy7Yo0ESHwWHQ
P2LO7nmgEo+wdKqen7SGOLRCYiio4uKvBZDwU1rlTKXCgc2a9h/CGuU63IEEIKlW
HLm3ruYu+G0BbG3B9s8MEJrrDRRY0+aiOwAt6veUQrLac08j/jrXjHv0eTS27uN5
Y5Jkn6Op6tulh5f6jrz22/VWaYHYzJBx6qcuLjw86QuQHAQNdH2FE1E4N9uxKuAw
r9BfHL9zdTXuftyHU1vR1zxv+8+yEUhAIkvnNF85l2cF4AGnPFpsBSsP7uK/sH6u
gTSs6xaA7jiWILk8PQZ5b+FkKiNNdpg4/N44FRq/qjQni65JlGAh2Lr/5LLp+gy4
NbIuVFP2zxKQvprajlKDB7L1Mwr0HEsk1ASvQvCJZDDv0vNV1lBKtlCWTmfjyAr3
eq/yomp1GUdH4wpS/8dFTsuVgYZP9bi2jB780k0xwh7fZ4WDzaFoJJH28qvp3iI6
h6iupEsJ+m5P8sd4b8FStmoQy7kYPLytvUVk2izzzPKBMZsnf0cPrOjsGs2z3M1n
nOSyHR5CamQ2+0MIfl5OrORyREuuwyvlsuqGukk/l/nw4/MwYPkCNR5Zsn6+D76C
CxLt2eucqwKG/RZ1uL0LJ9EwqtQHcmJYLyo9QlmWzbD4m+horfmHwwadek65LgCc
atJSDvIEJTndQqIMVVA7CU2A9C0KWyBkVzR7ZukzELs0uz7PnMLoc0gSN/6nu4fP
fBWizTOVYUOKdUyhWri+J7sz/f2ss8LuOfTKoJ5nJ3qFNoaRFKIOF2goSwHUcy00
uJJcYrAx5g7DrggvTE1hCy15gamB9ltPnqMZvEJsIz6LjQk8SOzTPZ5CsbA9OkfQ
xlFu+y3e2O5Xf9qBA83VhUr/pO++8BE+/Eg/ITaOh1ByssqZnV7TrcTzYI+4j9bF
PjNKG2QE/nC7WzKAb5uBwZpQ89fZUv9zZS++62OvoKVIg3JCWHhTiwhQ1/GLUKX1
Vt5VzCqrj067XEFNjGf0c+ju2xWSRKNHeVpKxaWHOnp1LUk/zT8snUagBfBBrly9
5yXMiPJwkilB1Dw02NZ9AWiyq+nPKvAgNCjh+k3FkiGxPncrfE/QA1564thIeb4o
QTvXPJYLBfmExXlW6A6TVgnNOjctooEqY0poGv12UgA+kzDZaI2A0flfI7oCz8ox
FiNqZ1LLRwPKssftKWzLmQZQ9czzS6pNEP2bnmP8q1Ghj4RPFLQ8Msd9mbhI1Cao
JqAj040YYQgck6Cz6rTSEops/zKYQWn8FN0MURl4/bIRsVDX46sMgOqTycfi/n3K
uVhib5pwSo3f9YA+P5B/TdKNqp4QR6cLmbH4w1noeuVy0YjxoeqhxdnOj/8alxeA
KDLNfAPp/btfFYci5GtdNVI1XbX5tC09/B9vCuqTDhL2jcYl2WWAeRMfzdfHmEcg
62qyvXlZ9qFCtDXpzSPqVvEPisMZXPBRZMIi3dZ6l+Lt/88bKJZopAgqBewSJe7B
SSIgFh0PaDDjdRj3vUKqYvGCcWxoPrsigeGGAja9oXUVteg2W3NN9PbTqp87ZEym
E7553BzTxOUlzFziTgruevPO0Aw2SuWjQZTxAJ5d5XoaBwlTSZ8ePr/emiMpMEBL
Sx+xNFfuRBoT/HPEe3iY/puxCh3vcnABbDHzb7t510D5+XD++oDgeWDpkIRSZ/II
DQUCVLzShlm0ULS3CdiEOr590V0NMbBbeaAnzfnOO19Cdh8pCWj4I2m0VFvd8w7V
GWZDMN/WkpgwLKGWdaDJnlq8ucZcWIyiKiXLasVkNt9ZKyUL+xWJbxgvI7Iqv8Uy
X+WaCsH+5UutfDzewNqzkW5ydIYCo0uIe3BWYvPIdrrvAOOEH2lXP9OwW03NL6Bk
mRd1Qo/OxSXZ1IflBPAi/Qy/fbIspW/qjE08FiO1SjqxDT7zhaqlQCGEjC+L3HPu
fJpEhj31XcdbIl5BrAaDrAXTq7EcVXUGDE5VpqWqcxPJbt4aMqDRrSmS9MyEQBuS
aACbSnnWR0M74HRlpecmgw20weEnHH/YLZNetOy3zgTNZeOebiSy7cr1VIEvJayx
A1f/cq8kmAOu5cPjc0S7/EbxsgcuGzIH75zCquMNIbe2V9BzWQOaEb8aNtNMKbwG
C3WXQKjkSjQtC03D3duvHLcwEjeNtn3Aco0zkaUhf2pK/2vpB/Y7GpJGDM1zUqLC
/56iciiYtyfV7NZqsW9L+HZR7h8bO7W6VOwnaEJSZMr3n0D63+TpABsLuXJzqTEm
p/3PPOCiWnSJGWwEAVMkOobh0VxFcd95F6YT0Jf1/K4sbsaeN8fImbJGZ/SV4P1c
ItVNWk5HcS42Zj3HwrYptGWjyvwArnDpR0YQd1D+f6ZG8GJc/eIcSvXw4oGyv//g
HZPuDCqqXsnHY5YPRonULI/jdyG04+sW38zCt44MD8u8nOLgXYsPDeihFvtZf1wa
nML/2BMhaHfA1MuLwWRWMXqJlTLDeN6dMG7bfjyC9ZkjKx8YqIZC6J90PiH4hYJH
I5igSYkx1bHlWsBivEVMJMxwAab/BQtrxPxTQgSAtETaEQdnHLcp6wvR+w+ibNov
0vfeCGljgDVvQxr4hMC0dImsYLyXAiiU/3tth9y9wGjAbFFDIOepV+pKpgBn3Vn7
GDk+4A6kLZNxYH2nfRZ/G+82GWQUms+FEHLhdK0VSOkw5FRcIhlx0tAz3KlWiUg1
bFu8cdzCc5TOa2Wz8frE7YRNRjFT1Hn/3LWNSssw6V4aLQT/Iv0xEI0h44vQ2wJJ
Epq0bdoTHRhHWW2aO/OpnaHiV196UeEH5lQsNOO18gpYmT1VkacwJN2vd6ZBGVnt
xM5DTeNG1j9mP5lbvhELCV+FHvwxk6jfAJtZvaITV+BUsLyyQ4cnnAVTn0d/EtHO
DIstgn/Tad9nUWMq/xsoY6ZQho9aicoeTWTK9+cN7Mqut43iMVKbqg7qzWcj/rOP
/eM2wpGGgxH78LUy9Mq+2bD4GD/otA+RitijOktL8Rt6XBtSOYJzLaJVQGhCvkVk
QOxDGmPx1HyU1/fWFxqOp5Ydmpi58lnKulqK9LUpZNGAxBwHa7B8mOix1tZeAuXS
muP+Qz2GPrHlhMOQdnfyyee6fuPebGS9O7HkxYScPO2eUbP8ufZmcqBTd1JSBXQa
4PV9VM9lQ5GkpJ3mBZhBwysfBEpTfcUp2UPcZmFj+8j2rnRWnOn29pl79tGcm7HT
Wk/c1M+qQDmueGqZHO8estQMNs86JBSYmZe+WLr1AeSr6ztNvtKJG6/gwGytz9oK
tk5h7PMWx87B1jJF1zNBOw==
`protect END_PROTECTED
