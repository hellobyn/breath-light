`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2QQhe+q3g2DidCrjeiGcXvYWSD8qgKXrJz0lG4geIsLRLdp15EHLVjOTYRJTXhL
+FMQX1r+ghFaqHHG7hnanj8oyOjz79G1Sw+XhJeSprkYrV5AWJcqkv69shRNYu+W
bhl5Oskyr8lRGTr223whWiHx4e2SgJiao/L13w3cMuTc7ecHWiFUWtAY4rvSXH/y
5aozxRe2Vu/zQAleGxHY8PKh8iapHVtvMR0AY7u4Pb12nl74Se5IKyYJRm8NG5CF
ndioogwPiwKyO8iDe1G5Vw==
`protect END_PROTECTED
