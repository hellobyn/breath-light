`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUT987pY4hMHuuSldOXHBil4nb71kmOmlYtRheDF7JdeJdJrfyD/WFMuhDCOvN0k
TVJ9CB6kAW+1i/sneCAh2vGR0qiwBQ3697yGwOGoldh/KMttLEOEI7QHc5nDcaZv
oQdhufnes6ZBbkIs9A7bXmwgcXGcGEjZZ5QKmMWmqjfIa3TeJK3CRKPPiIM/9nIb
4mhNZZqNfkwbhvKC8BKR2DKg2lioGCfWsAPloeAcu4UebMMhA/WqLj0iD1Isg2jp
QJnB1bLEJU4mSefGuUhWbLbenW54if81rI1eWIqy7YWS6I4RI4GOTz54Egn6pcBo
JzqGemQsXbmQuIuz/jP5T3AAQOYeDVwht6J+Aoo66qyhLHsSzeIBj5iS8PKxk3bL
h2ci+n1+ZKoanGg3zZ0W+/s/+9+/M5xcCkr87Wrt6svqxPhFU5z/TUr9/5OgwObD
ApjyxmYlCwppKZRoGDFnXCc/K4H3oQ4fEEsqfNMM5oCjHEypM/Y3IWvbkKQmnIRN
9gCJLtoixWNXEmLIeU+UBBzAx1NxnPkceqBl6XHE93j0Wz7t3FyLXd4n6yV/faYq
t1VyrGF3OayDC//Pu/PhfYCffLZk9jfTlJV9BjnK1y19zPFe2ohls9abocDUgTYR
F2lSPMY2IeEYK3B23W6gjpaTVfT5hJNWJ2Cdh13wrKE2ryTlnOh+djQjhdVIkre5
fYiYDPr9xH6iK1p5vUrVwv6nUyo55QKcMVluXg/Sm8dN/lJ59977fNE0aLGij51Y
zQewj2Uie8Cr2+pYcRL1aZ/sQjFsQY1WozGOrjjn0NB55G2e9DwL6Uus+3fRyMko
8vijVq4jR6iBBOW22gWaEobl0eLMTTr/tx9crRcpHCATkarXegmHZO2vckdHM/jt
uyi1Gsn1PSLgmoIh+jLUZXsEUWJdt11fVv+B3evI2TMEybggVi43NLgKncKEAc42
Yz+J+E4QSreD58jjGJvzo5vBz1KpZblX3njahaTvFDNy9ADoEZU92D6Cv23RrHAI
DN3Q9FM4BdczR47G9TYlx2XopYCDp4dmYCvG9D6happS5BVl6lnlSulP72lFpVob
MjZUyql/MKVuwgVQLSP1BG7PJS24QWmT8/M4cYN8M/66Zg1NvDgtPn73SExC+94f
L2/G/m9LiFmOAAuUmnSecwImaI7cPpMBbBmQUo039QGPRm1wGZ/xwtWLeatgOwbc
3sET/kejXmaPefCMJLJl1S6n1yDzyxQu2ll3wfBwvhLDYgjkdMYNDb+E9qe851s1
lvrMr9aCIELYcq3K3iIi79p52ARV83XB3+M1FjMRehvZ6oFQ6umqSOPhR42UhJ1p
QGIoGdA2CleBxiOkgR6vXgi+f3lw/HsYoaw8JW0xECd6reAqtp0mQ3tZCK1UDhk8
ms7nNVQqjNIwwfypHupwql79Qx0IguG3gdMqNS76UEO1L8eXpF9UgduC62jdq7it
sWebHnH+t251NoGGpQ4TgZltU8z85pdNWI81UtG/dRa+3S2MHA1Rk9KodEPpGz5/
2I11m3lBnDR9hs0FRHO15ACRD9KEl9tWAi9vhO8JGhaFmP3z9PbQd23pb8uoML56
VpWsgHerc+DDQIVhNlkj0h4PDfUn2PyybNHxnGKd7Km16A+G3l9dKd7+YhHnm0nD
aiTC0fthhoVEDQKL+2UWjuGGCfmOkAp+hrsvlmbjyBXJnCaQT4qFQHdW9nkupprF
gPdGawPA9VzI5juOMCR861oEiKYSqSP1FruwwXoh9DhRIqXTaaKrFbB02QAlpmXx
jL+hj4/ounVqvO3gzoJWxUmETYG2A4Qtka7LlfarjLhsmZyFe/ldI/y7PsK18pY3
K6NaOakHAWY0yUyg+Jt8FJC4fGVoFDcfhmjjnnQUtFc3fyt++6eD7oenX/Nhmotl
ettj26lMlDyXAqzTCIBtf24d9wnjDyu05MonWmqIpC2j52N/7xkTDSrJbEcanKfU
D5M1/XKwyGEE8a1I39fQofIs8slKYNELolsERtFDjKiZ9Qu0GPJU/ZFHsUbBG9rz
Rf87a7aYsJ3Ze6QBepvkV2LsLGqs8KPv16cttGFJHC6FF5iMX9FROFqr5mPULtIO
BmN5Son/PiYyqVxGPwKa/uzCFU0zQd+oocpCkJ8lUmLZZXFbOmRFv7uDm/WgZ+bP
vzGKtSwj5CFB4ghZXjR6Ay/m7gi9YKtz0IMBNCrja5pEt3t0G1Z8Pym57RXXp4jl
qP/D/RpA1oW9Flwn8Qr5n/yS8z14df2SgN16UCFTfquicnc8isfJteMN7UiHwmhj
UbSkSq6MCMFF7lZO/QGFxbdWBl+9qy8B4K0s1HBSzMnA66ZSVn5z9j9TovvGwf6g
fjCT07c6cBSCkUmKd/OXatjIYpMDXNRK1JTia9Zg+2Ta00qb2qLsYQD8dlCf5Drf
XJZNkChW1Rhkr9eS1MwdUvfKXRqKqrzB0dbgmbJRLg5aEDSWtxN1y+4RAyy6Szfd
JM/1hIHUfMWNBaPAz9E61apFwI5b0Uxx6BnPiQkj1b1wBRrZcdzWQ9fgoFW7wZbB
e8tN+KoJsSkCrfg4Ozv0xskmlwJ1+CHWXh4uEUxRCQU80bdA98u0x6M1vzszB+Y2
Q7HygIbR7HsXWTg69mXFCASZ9+7LmVj1PFuBrKPdeWOvRoAIpNxmCCgfJTWkZDTG
KMyr1+Wjf6UNK7Z7QGZHru+dt6hekBCwLOM+a+yj76V8SwbZ1rRsXtirGjXt3wKS
/mSW06COVxkRPwjXEr8881xkeaPZkkYBXngQETIlPe3KhWhyrY3lrPyJ9vWc75ok
1EmL1ApXtsnBTIFrj8wFcqCMCb8ILdpQqiI9Mnrt7/JAIDosQQcybV+74h09bcK3
1ev+gV+xU3+d9XKMtNHl2wbjMcW8v6tg67HY+oDYVDd9afwzL8e+pssMorPJXKKq
jLTicH4QqBswxwG19pleSWU88OUDZRhKlFaz6O286qZz7BkWKBtLRJN5yQ6Ub2Do
rbriCWJ/hOL/ER5Bt/M8a+dwhi1Nv+27/KCK57O1iDZbqedq9EkZWJX8oYQPwPYK
pS3cpePZz2d+L6MSfjVHSwR7EJkgPOE6rG9qaJTdpIjpH0pJWYr8xFzytfTL0b7U
EflHIqpoG7KsOkjouOrv9NAhsbd5VxGweVkDtrKycNc+Sr8ra/nn8cK2s2Ikl+T6
k20AaqpVhrm4qXdCH2P+04FWZDxvx/x1M71ACSQc/YkduViLGU92Jg5WoTdifvdg
/HZoxxgrSukpJU/6SH2ssWhXvTmnezj8ZO1iO4jG5oSCsyc77ZyQSmHKLcTMeoaQ
8qBH7eSsETMZ0zLTzp4ZWWZk4hxtFSRflxi9HxcRFdC6xFP/MeeIjUIkmNTKT7uy
yKBpW49IC+//SjmiJof9/LjAKFMgtzKXx85HAdcD/m0YKTRCUbFDd+NxqkEUYl2p
LhKAmiy6/1+rZr5V17EaVmusDrkEJq6APfvpkjoTZCdV9yVrC2w4c8Te+Zttx/1K
eNAabJ1yGXQOmmVsPM1U0anv0hLkpWxsi0uTuiHih9ZzY2vWh1auqEW79sc00T0H
luLbdVKAw1cQwa8o35+sNrk+jzSxPxYWifJi/Jx38FKfI2LbQs0f6NiQ6mJgdOUK
+BS4+hxEZFUrRSAhSajs/xscLitG8cNmCsSZH7Ih72vdX+QN9JZxnNGNnCoSnAID
w5/jLgtl3OVkijXCYEz3DN5rGBvPVbXWa34urKDUmTaEINRtxUni++PYg1hbfPDo
oAuQDCfyawyLdowaDkXuOec1aHxYSoyFO2a60vKrf3Cjrl9TAWxH8mlg1G3Qq/4N
W1y8SAbIQN52jV53wr5DE3YVJOnyCZQ8Q4Il+itRstgn0LGqojt/bJT00MrSIqn2
j16FZYHhmNLTDmEmIxQFJaGdf/gYT+O9LbRyzHvzMwVR1Nec+WyoJwKtiTJpAZpt
dGO65U4TNZRmA579Ar1AygSBqt0pNm6CT69W1wwliNqPaKLQyZJHotSi2ue8YKlS
QlV2P+KRh82v2/8RPwDEXQoIFq2RkEOCD0M3IOsJCiHcothWFNwR5onlxJP6O/HJ
Ajvi+9MWFGUWUrOKE/ueNTg+zADSBe0fSuXjedmMMyVZ46jkHW2ItuoNRJIbsu6x
ud8o8j27KzDDAc8PSxlZ0CrNLCS4RjiHF965v7oh0E4g3br+NhljqqIacTFrI+CK
JRkK3ou4LfXZCe2DfYI3qfDWyr1RYoifdNZ0fk/wRcYJuWOsZMr8JqGh5YEoyUCt
RiYVAqr6+JGTlm/XBWZLCm/WODvMd7ufDr6KtCjbxb2Z3B/YQv8YPrSC547sOUSI
6nGdT4xAPOJnX0dKnwQ7P+/tysYGRiD/pO8pHYv0ElXIeqmjJsNjLqJZB7SyrtYO
ym0hayiTCOwtPOcHOKuqXI+XKm2j/OS0VGYVXHIDzF20h/3tNJGzlsh2g1jNsrGD
yq2tLiPKCsFloYX47IjSwRHOHNRYLkckUHyisD1GdWrjn10BnDN8hgmpI4Ka2el9
M9CTDfkFqVRYid4OrUMROTy5ZoYvy/sgFzBGHmq6vIL29Xi9yJ8LUlkrUnYgHD3D
5m0GFr+wDO5DTXNNEzEBcBQmHa/nFkvX45+nFdCeesz3gCTQOYNQzsDuRsw0rlp6
kFeDkx8mFXH8OkKsCrYDKLkziwLmgV+9aPsig5vXzXk=
`protect END_PROTECTED
