`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kQbIOUYGJCMNyu8upeiRACx1U5LFVJmyCetF6o/SP0dOdH10JYDzcnX8s6lDzkXp
C8BvEh1ptzjkGPGR+BglskjjTZVn9pvYPbPptuvFpI+0O3ox/OGxIvnA+BNLIpTi
eUbnOy9XdI7HgzrseXTqiwxkjMJBVKyQrxClNGBvozfv9rlAMBS9fKu4IzY76Vfn
eMX0FODyseQQ5uLKJtK0rGSMEsEp6tV5VrqMpK05/ew1PI4vivMvWW9JfqN0lGj4
Tdw0nAfBg/+oufugTwifjdiaDnq2oFgocReiQboNgHSQ8y9k8taUupj3I0v9xOPa
vxkDPI7A8IawCttX0A5KYMa8pB9nTZqAHdPscDq72gs4cZ4Q943eBL8AzC333T7q
LXmwNsSHAz0MzZ4p6oDG9FPhFyaPH0NG1MVJefJjGeUsowWClZChK6Vpb5RWyCQ1
COjfESAE/StwzSCM88yhMDFsjglrams1bZs6WHhyeAPVZ6YcjbR9H6eOGEp2D/b4
Qg6PC4UKwdSfUxkqbCRoKG02T6rFuLcengujIwzapZ0HyVmw6ieoHrQGxWePRYEj
PKcbhE0k+NY9452xvAHanZpAW6E9MULDnuU97LXobxP4p+t72V9fJgHu2LJnrlgs
50kN6Te0QHZvxaaeZATBdcaU74MyRwW0YnVEgk74FMZwRVuN+BS1MktfjRjUig6S
w7grb14l9lKjtF7qv1+vPcqEoCD2jJg8aKLSY2AlAfg3wPuH73wziHQv2XC1GIog
r3nbTqcNDdzwwC0mSOQCaw==
`protect END_PROTECTED
