`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdqaaQXzmi/JKygijxjJu2zwKFb8O5aw5NJIQRs1wk2cVnC0p63w8adFpYHnmCD6
E3PUYmrZt5vMXWJX1otZh9XvEfqx1vglnhantDk6X9tP8Nnk8zgNf+1xrNVwu8pW
YddkxO64bWdcOcPNBu63iis1/7nHDSaEs+R34x/b0L49ONP1dK+iiKj8xW8HG7A5
44cLn7rNPhAki19fCPNJqJ/kePbWEaZFVVRvFsn75X3h4zMZiDjTgogAgd5YjgIe
Dx5n1F+OaAXyVOrVUTxBjzytzBO2xaptyjAW5iKbMI8NEF2Ga0hSp2L5Dh90wiN6
5+Wo+oTGdTDurGjxAgm4JUXw71MIjqiQhQJq969g1QZ3SNw1KcbGeLdgfd4VEVCL
zTWBixJ97+5O8V7drzOpag==
`protect END_PROTECTED
