`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmcVyxQ6xzmQ5nGEIGb02lQ7dfvsSEo/l0FSbUSdOr8Cke2bCKOWLrFXjen8N2Tq
FAcU7Td0UCp5VDAMuJo5OJIJ5j5QKQOMxefMdnvgmno2qxh+XSBS0yA4heim0DXR
3Ew+08fVxG0wFESj7EUwFKCBFknQfbzelI9ZMqjwLnosI0BOpAwh9jkTvF+YeBVZ
+Fs7K8tXpMmwlJGMWfTRUJuwFsx8y1l5qZSCSJdRWGOdv8OD24rBcL+D0f9FBbHZ
vN4N298Ywn18wmslbuXpcNl/cJgVF7uX0LsUNWcYweI97F+1Pf1lAR+l8pR2BUbp
kbiTnLqoTQXmyx9+95oadMCIHLyGB92KKk7hDOv2dkfOE2WoFx9D9kKVr47BW7NB
eSny+oAGP95HL/ohaYGdzddb0urwYYoDLl3m8OPzBjG3eGyVc82fh2vqKXNH5q/f
Wj6uxWtoOtiHS63QST6aYeeYoCV2/1uL/y0exLcIUTrlFBGo6mElVXNXzxtNVTwm
3L7SXpjdBTSMp3yOFQ7KPIJ7mDoVh8e9ke4c4ltf7ELk1RjhpyBbjciB6Qpg0FUE
yGUffp6V4sRmtL4xrnNg6fW6EVLMXOb7Of2PnS0miVipmI8wyI5Ix4MTmOLbQe3k
`protect END_PROTECTED
