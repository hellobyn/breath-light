`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CueO2iL/Rq2B7PtRA4I1t3r2BOGLsTn0FJrOMn+AhKF5ZBabrkElGppJFI0tyeAD
4cG521ScZ8exuh/cT55O027VQA2z0UEF7DEFA6/FRvWXtr+NwhnW1OhXRV/6oN0C
lfQ/9vqPlT457wWcssd+Dm6i0PkfINhrdpzAI2ThpxcU8pC+Z95GzRJOSqjF7Kjj
VschbKC1Q53I0ENk2Fsj9SjLapAU0+WCIpZL6RYKHYmNWHLV/hWnCMujuXboTNoi
1vcnSYt3MtGQCwn9B/VAhfvgXaelPnGqzL6O1zQ+sJVxUaTjtzFkMFaB1tRpKrJy
7JRhuUO4+la2Ao5f7rW8zeAnPox6kRPTdkgxzYa8XXwls0vEcTH6alWHwuVfBrGC
zuXm38umLWZC+eUUL1nbQE1ku5foLrpZph7yYYc50TUyJIKg3E0GTAjXhz4t79vR
PaszjYDCBGRshdV7XSpYRGgNlHh7/V1MDTqHNLLa2RQ6zQfBMqHkkxoA5FdeUtvc
4WaQrORC+iTC6mmpzha1To8A5mjvobInBQFngemR4UrxGBmg/xFIts6T2Gb0Ky8B
88Bc+HE5X5cbgOo8zYxUMXTqOuuWVYBXkMdSx7St32Llcldmvc14Fk1smRXLSQpq
GRjQg0HsZvR0Pc0zAmo2sUEElcVGeKP51CXJoHP5mhhZ5/xxmokGObvphwT/DEeG
+aLwOdB+HKEl11bVWoPjbiVRgYcDQ25aMzaCUqFdoH3CLLKN/s+OdzeyvUIQLm5+
8ucUp/6qqxf+M0nM0pxWWxbOL8KNvrrLp7LycAUB2qN4Q3IUqBqEmmCNjNf+bIUo
Nk2aTFnY2fjmO6E7ndjoKDpVsiNBz2ETL5rpEEg2GrIWsRNTrn9FAQrQ4eJK1I2h
WTdeeHEFuy5BHWruyNiJoqKhcw1/WF9oc/1s6C/JqkPMvNZvd+LfI+DZJdn01wX+
clgg9rbS3Tcspzb7XK+YdQB1uwaIHzg+c1j5SeR3fJEWBWTNhEfp3jkMKm+1BCVb
3+8Z8jc4hbY+UxChqRsvZG8v7v8djKqVMIM+U6VlJm8RL29iHeVyRARPkJ+LBakU
p47qoAJaHgPrrHcoSJCHyP8OqZnxFR9snsBiR+mTrUWUl4NAQNbKhOkCof1M1fcg
dQcIqP0D95nt/Ctb3Utm+sYNn1+5ZvPcfLcu7VQYpG7wqkyKK5/mGrZLc25GBJJH
CqPRemUJRQzRd5Pe3sLqB3AO3NxnU2PReIymiMyUNN09YcCCLQgHGVRChOYfjZYa
a9i47uy1TA1oYi5PFksKJWTzBo8DCmd3NPoXg/L4YElHtV6wS6eY9KomLayYu/7n
EsBBvTZ6D2h43qCNC4564WxYKOpfYG3Euda02Xh7biHDGNZtigqZ23aD0RJZEOo+
wwdZIMNDuQnDGmLM14uUk/qEW9AdTYU6o2y3UVGaIIWh5Ao2HrRRf/+70kSPgkHQ
fcKkevouvPnPUHNkM90IhiuJxhXpa89oC3pxFZL4Bz39B19kg9TLTYc1RPLm1h1A
/8qznjtHoCWvLRNlA5EfCVrlhkKKw7amgTvuPI/pI6Mvpcf9pXx9DboFuBOhcRVY
WSROuTq8t9Z8XomjvyN9CLNHVcMPPfeEAVuWSw6hUT8lX/ibEdEtZ7xpNnFjHszO
G2B4m5mzLBcMeOXUu2zrtssCKaQ6VeIcMDQnLAaX5SsWgu8kkLJo62APiPDio+/E
1gNKelfMHCyDhb6saxWgTKS0Nrq6YNdPmvZKbkgf4iuKaosz6OdAlEgJgg+s2+VK
hP9WmM3usVryKL29LWcBClB7NfBjWMuVF1aw6SnHzS0B5X8kPhgg2Y9kOpCH2uzt
86Ie5XXHC19fn/26jK4ZIgUL+min6broj9V/Ox2h8PmH+BVC7tE56OG+wvtBNXHG
Md86fVSuMPnreOtoS6waJ1inmyJMvTgiDRbWWttHzpup7NZYEFnX+hglK49BgTy6
TO7KEkpNVjf57IcOVnlWM/jDE2UccoZBDiFHV1wUyWq8JWzdxqEASqVVrBUz90nt
3Y1sWwBo721gaWmVMX98xcbIwS0MvUbimzMqTmHIPiw6VVn/TloPFcjMN2AJSpJ3
YXuy0t28jtQGq4iB2bcH+JPhVo02iF3/A6xSspXdHrJu4v2GiY9fWaWJGFc/lu3b
qZQt1A61Pc7P0rFpRrhG3jA4F+QcdHiDFBpYIXSWfKgoWvo0QPmHpAAmFtoLPf5w
B+z7i/u6rWgSczbuaYg36xEVQUcoatoWvMW+nQZftFq9lf5acIR4yzFy6uHK/YPQ
kJ6AVTODx0PKfpqtSwPTodjkP/JcLvliqEaNMgx263Yz+U0MdRR7OArm+VntQR9t
hjuZ8AoMwct0JiyVHOfMl+ffQ+bfdf2aG8TIN3JBKsPCznFaLGwipajhOJDCZcca
oNG2rhl3fDUrA9zGZ1O64XpBfoiCHJrWuJf6wPtiNZH8F4BVNjWvA99ARuwmMowk
+hwjB1l3y1LRwt1o0S64fl8eFoAJ9sOi7jq/ockulp1+UAa+eaSOXOw9r6yJb8cj
wfpqwCxpccBOzBrCsQZf+f+Q3H9/zMxBswdsSbcZgBaHiPFQ7cbhncPkV5Y5CMmE
9dcGV0lhBIrkfe6uR1ZfQ9+IejImq0rcBz3tCPitBaWs8vkoF6F4t2nHcB4Gtdrh
QrT8m0wPIGwbY9AmW+SJB3c6giVFD/wzczjmwLNdjTbKerJumFwuKHIvrcoTX7aF
+l1VNQnuQrwU1oa3wO7xIS/hLceQMoMylXjW7gCtefPhd6Yf+SJzptpbNpBjS5kv
q1j71UgoYgYzrMjWJe3n3EKmx8R+vE0Oa0XBgGKYa6QHzGC3GZyGHEQzuvLMW+zL
eNsYlmbZ0u6hIDtsNy7qGBc9YQOJx5UbdS6UUxIaSBSiCkj8r5DAmWmKU4SK0f4S
Guv47FPmSgiAVGirdfMn/4AyHM0M5qpR4wVoWxQBr5L4VcydeMc5ko+TwijSjOMi
ViKIESlln/qalZf24QAlUmAtUT49h1Gl3Knf8Mq3ng1924ryOgxByQxLhmN13+HE
mEy2bRqBbsR6FLBMj3I2mRI82wnD5d8qRxCviBvxr32wrd67GeopF/3AgL3c0A14
2Pbzllp3kl0gKI0mVV8Y657mnYFAMQoMJluXaNNeXL2CiRqZnF6aYU8VzaKMS/sB
7iUOJ3cRntVWqsemzNLNM7VD/G/EP0oGEpDHVqR0f7kYnbGo/lHixDKS6DXScV5V
RWFCq+o2aB1MaGKATuIBJdwlcxSMUA0yDna7nW8XwwJr0TxeMDRz+Aq2PGQI9G+X
Ga/FsQbsxJL0zaXt4AbAurPWMM52x+1Liis/ltzasg7gIMfisSKyVjKm1fyyPM0w
zAB9DO/0kEbiO6Qnq+0lBtuK7x3yL1fMMo00S3VgKxbrKBqtKN7K490mNS3cqBR8
Eh39zno0KRqMaXYLTHgkZpRwN31HGARetMAMq8tGKmXBYHl4GUxnJRfgXABcjdTA
w7PI/RtMppuvjQNyn5WFvH0N7IdwnKOryD9DYAHGzNvkVqBx9fq1BB/xIDL8nNVt
BrKx9+ISXoxhsIlBCMOlpKp5iXH/1bgx/6u+W/RUDbYOV1gzSmVEzGeHk3q4x2wO
M5XMx+dNRD4x/AIYDVZ3vdeVAzXv5cE9rkQONq9GFdecuDRZh4DxtODPp2k+zQXx
7xxrqo4lwzyJswYdsbvxxoSIsVftFXKq94+08LMh7wS4FcKy/Em0TGHtIEocH4tK
yf0XVON8xM7ZpreSFRfPTl8xr/Xo5UUGyzsDQnF01NOMGK8IDuO0s6zucUIzIYEg
3Fj5nEahEBLU7uTYrkSVlg9aLduz0IxkWmeLMrqA8Y+yZBOt9cYxekE+zn54hqGU
kGum9aIGeP4XyQRTCqMdpZzDGOIuz6P9SXAT7BDWLkiDd9SbW9uEKO5S7KXPSUgJ
IAGPQDkKMfs5t93w3XHodTvNoWBSsinbM69BRkmcklrX19EJnUPXI077MUuxaIfK
y64Z0a/iV41U8YxzDplZHlrrQ5qGy5749gxyYYjOAwI40S5eqFooffn9oaNlCvtT
fCpPo4k/EL03TcVNbMvBn4h4D7i3Dhpd3XGN5POeDtxjku0Mzs48TqAF+tlmSWJC
1TxW41E8N0djvfarScpGiaIcenMtEX5EUbdDNcDZxJ6GRJoeVsaWctr5im8O+oFd
tNWVzOVyqK2udQKeJB1821WwGos2MVzg7Bz5Kmrkxi9vH8MQnA2EWzqFy3eJ3esh
z8SWyDDURTNF9Ya7AxPUpkVLiY5Vm5Xg328mAfjek6IYVhIiWiHmHDZFoHDPJM1Z
+I4Tr/lPvF/0FXEU1nXtCukOfrNZ0u0h+za0IaU9KOoblidu+loxzAaxFTZNgmmN
9a5qG0BKQ+rudERfk2iEkWCiLar+x21y896YGEgQlE5dwM42SPosA8s+pRN2ooD9
yTY+Gd6+BoyGI06Fx2a/IugDwbevADAPyP5PNm+pPlNyjfPQTzAFXbPGOFx7rZ8x
7qOUYOq6iDFf2JNjKdDPgLJErlZouc8Tqd49y0pE8Ra8RRfbD6vO0iFl9cOZkJRA
0jWf+i9yPqKTP2u9bNa8gFlSo+XyaEx4JIZUng26lf0Dulc2OGmw/BTFgxGs/epB
jfPkSY5niTSBr1he7Eoi7Zd4kJPdmlXrhtfHtrLBziT/BdLcTM38VLdAd7Vei/Aj
DQMbqmVLq9PPPruoE/eP/bjgPfhUz1cVr7U8mYlHTf3xC2O0NYKgcMNeYhizXnF2
JWN1vl7/2OYvl+IKIaM0aR0pDWp1Jq4m4lyTZxrGrjjh3kdNWffglBf/fd1k0Z6P
vTJ9g4Zl4skqd1TBphARPRAoYgPjsrT6q8Q5zyg2aZL2clYPOUcuiijdbkpOv7TQ
o2iML49L5G6lg75uNumsyxnqTnPTwTzS5qlFr++4CzHTaZp/HMoP5ZKZpwZRAUCQ
+79XRNlGM8aFUCJf8/maSG0TkeL2PY/s04RSv273k8BzjCEESO5NfkJNc25BZGOn
AoiIv8Oap2ZXnIgHgQB6e2ZBgMX23f9CwMJD2GOKqVOj0RJuB0wiKGuxarYn0WMZ
43Hy/ECBlFE1XNLqimx/JbaH8gH2+1BVI9wzdqFx4jHNwSBG9INJq4/1YMa7ddlT
cyvnjRq7to9pNTTRJno1MVwJykL6yM2jok7tZYhApUsKTBl35IpeLligFbjXG3W9
SqRGOeyW++OZ+mU7OXIT1tWIUjkSYm+QysETPcnfTC19vYCf6iD8RSCLRwTUe5lX
bMKUv/UrgYX+bId3eO9uXv/Jmw0eoGXucWQecREe4xz8aupAyBRLRnrydFPszdhF
yapZZgJCvwYI8EM+C3H9P4QSch/me6GrZdicMmtBcosXjBg7T70ZjzV1F1G7T0K1
Ea80xDQK6Ehwyvj1Alyd+hv5yBL5f1sGC9RJtai2wdpzP8qKLnkFks/ujLBKoJv1
kpc8fP4HO3d/EFieqb6SeytljlpuaHx5jwlVTqKvbVNWXw1UTaTblI8PC2mTxvDx
/0M9wJPtE6HOcx1xxHUE3LW+NlwaOerEe0PgMnqwXH5plbagE8367jy8NO5JmQPA
CRvOaLMkmAF22wp84JtsYLMwLDt5NkHNzdoEBkCKFzh7fkAYGrOASCzfXgpndkZY
+mOB634BlnngYVXpovnzKQsk/Spdbny5rU4r/TLowDnW6NHUWKSRZfqs2Ty4spBf
PyjTDLoMnupSvW3YBgOwNdrgecf76cbvuLVHxWN81H1xDXZ5sbTKXJUIZu8ypzjj
sSBt4Vy3kV/c0SlEHifRAw9cjJzeJYBXVHdNHDo+TziRm89jzVyILl5g5sXrvwOu
XWmEcpLPpnvr0Hc9aUon7jCkttHOwlar/HUunmXU5i+bhbk+YTlQJSlec2ue9Yye
YU6GW6vpn5aAhC880xR3cgFtZjJrkPDhmFNgj63gdqJ0ZcL6QTVy+o9+PgWqrcV6
zMssE0oGbsx9SGXGzMyURjhJTPsTvuwXEDbLbHbEAR1fqB8tJYFeaBRAwJ0mAvzv
77njJpHFxBN8lr1BhpzxmjcnrGyqWK7lhTjlVoUZcJoz2H/MlYXFeOQbWHDq0T0r
vBU9NxJT8CeWUxlKmjAsfktSrU5xcWXbc0XRG6OLE7C+WF6k5UxK0eHLMa3nxYL0
sWmYUFiI93Kn8trgkTWBlWCQxlaqaiekGQV7J3UFqLZw6MYL1s5VInECWEp0/jaH
jrjDMQD9C8HeWYTqC8qS9QzdBCRAz4NNlhW9VDbeoAHs5CKE6Mm2NZzupaRa9Wpd
2d3f4y8BGG6bIAj0siiKIF166GxzbKb0is47n8D+cIb6rYiqwtTz9GdkcegLig4q
tXSrYEHe1ztBmg0ie2tO93HcejUW2uuHCsQSL3XUNzYcozUR/uDvOR043AE8Ky+q
KHcRD8ROjoYvR/cgfUCXER8a8QGx4cF2MET+OcyMreCSdUHPG3vaK7Lb2ACCIeJY
XFWUOS+nLikjjwcN0XsEBoeDECA8iWtFc/hNn11pUXFMs55xEq6Y7MH5JpS11tRu
T8ipOZNXHQLrP82uMxjyWtgpWjuCtx0tkyOJrlj54x6G74RpUpEWaE3R/btlXCRm
sIfMCb3g+DEFWpYOhVCKfFLjfkDzNPjgTVtdp3dpAyfmz7b9je9mUuPHUI5Nl44A
z5jxluFSn/A4uB2aufX5gdZ2ZJGODW3WrbheYXdEXfquz5p98tMqDxs8tPI8Ggwz
Ez/wgzwc/5PhlEKSdCPeD5tfusUfKOb5pmydhUOlpw9RrbZIQkRrpcp3ZzDLpusW
1T+M93uiv/NoRXmAnUu/3uN/f4lxIzQBFWjpMAcEAiJlB74bEqjECa3XtuZOKmfg
j5jLmZRE5/KzfHnA2BsYoYKtoH+MPM+cSgOlapy4RQjSf2OCfWHznKdJo9O0E/fh
TMjJqqjIxvvHrJGKVOUL0wUjRa8OcjkExCW8qNaIkrBj10pXpNi1LlP8jvz2jw1N
PRtaE8cmM3z1iCWT2yosUErIIkmenOaE6F4CVLZVXpEpmmVLP4z3YsT/j0WuJD4m
IvFrQiL1nemahJptcpw4K8v6I6W2fT9sOGSJ1urYGXV6f4qOls/6BXRejkmi+XJB
pS2SzT6uXx1kmV9Rs82Vhz+hhJ69w5iD4pjAqWGf+8HytjSaN7ZKtaAFjs7D5gZY
g2D3/Jk6Xz+PSSTyoOGNHKknPq7VeV4RGkSD3j5imsXV9hlqH12wROV1O8ZZBLL6
Zd7qhrLE8/cYbHvhwxqv2IbqBRB4rUdt9w3sjWt4rwxmqViBzaHNZqH9ArObvzeh
y4ZQXzONFyc0aU7EnERyXrj5EzKR2aOgYEqe8qZLCgxy+UNwikVupbECmFeeKanJ
0V7hAQmIJ4VDnwoY1hxeJVSb3xf2uCGffKwPtNukH++3YD4xwp41IRAV4icz7wNt
6ll3bLQ4iWtPhm3acG//NRHzk/KOFdXBDsFwmYwPkO1Wsp65JaDQcRX5ULk4q5R2
bffHI4wZvb77xxoyk/pkb2qMzL/s/FUk6uvSbbE4R6J2UeXdsysPwByb7J02m45Q
1qyC8WOJmNrfJYS1qKhbkdigd9Ydowxe1WAsLR2xZUpSJui4xzzlnqgd/4fwPTJO
3INODMSzF3wIAac4b5bGMQ27VD5PL0J7wrBVQf5jeR26NTbFEoMD640+IGAQ1to3
iLPdNlfHqd3Zk4SV3d0Uj2aJlWvUKt5yDhaehWLIpmm/dEKngaTx6ibCpqlIJWSo
mv6SwtjCEi/npciCtX56CmqI1Uq1EioGFLuOY6uVhNwGMeS5QWki15GEuy3rLDxN
b2PGgV2FG1uMVjRaomSJ4ArqxrV29rkWIdgVg0U0a4Bf4hz9L/R6vz5C9SeSeuMV
BYDtWUN8Chzv9ylP1mTHsa9SiiI8sJx1dVhVchDQU1GsrpQv6b6Smak6uJCtW03F
0wwoA8fFQDMydtKnNngqasV9vuEpxCofM8zLTZGeHzncCXH8vLwPJ96NlXItKwZT
vNo3c9UxT31qx/VOjKTT2Zn8uONpNtMuB5qtHzeTJUrpqwbzESY4biDLyAaebqXK
MX41d9gHSQx9yE8avYPLwoeMROh49P0Bryvk3ythUaSBXN33lcog8RjmE8FF5I1I
YJM5mgmgKJ8mpNtlhcLA7XrbpRrGUAm3dN17lSsXCGuPlMATk61iZS4E+nd5kssg
r1+7c0vSHtS6qvUfNciYnINr13REyUxxnvzVtiZtpuJdBNQDDjIJyYlWF276SYsJ
KH70kTiggKfaUdJoY1sAe8K0NBYPwcrKYMon7a3MZ7AcsliRrCv5J5m5os3y0kZ2
j8HDNnO65RI9N+E1NGiy+cS5edg2QME4MWAS/n37WaNm6bOXnuX0+mvZEramn7CQ
6AR/L8kC42j2FYN5eJ4tgBldwaS2QF8IbCWrZxKyWL177qPNJBK0PZ23VZNMXMdA
TB4L6g8n0exghYwU+R/20cGzfeOKVTHThoxZZLNFOXt0aGtCHXFY6jrHFHYqkNaD
5Yv5Rv4NGJA5JB/EsSrUGJRpyo0gdjvkefbENIAmFvk1ARtfXcicH7fVTxZlvP0S
GGqx31UFbiueeYnt2F47Ykspp1jF4q6jbw8NaH9rjJImJXfLEP//Ez5hBsdyrnd0
2r0NeQiR2eD81Te82mWrkKkxRBNnlCTiM67LVKNDM+jBUifuAqZizmcsO8MYXf9m
SvKEd5bTMBYJQwjMSbR9OfUk67Cz/IzXQrxuan92Uuk8t6DNMSgkGhKxO69dNTxU
B/9n2FVBXvzNPNs9/jTOYfKqiW6dam+J5eVF0Xa+V2BvQQxSvERYmGhsv5r1HtgY
lSoDUw81QbR2WtD5p7gD0rCkPKyPE1y8CwBbcFCjobo6lA0GDS406O/JbkOwod9V
xc7jXzIB/3jGYHSl/thvzNdTxcJIrLM4UMamZZJdUur0RAF9nCYPEdUTVyA+dpmW
Hr9KgshmhyrvEYoplBD7aZHFBrOrfRCwm7AdKjUFXz1cbMy7SJgewcPOGwPaligJ
x0zjJReeU6Qkt7whaoXnWpy6Bp2/FVlMJmch0N1OvaBMaeAFJUilYXn4KHDlKNr2
fsCI3qBMQOUwFshlXR8ZdogewA18L2fEAG4fY7E4d4UhSZf/af2P+Y7z2edBs/FS
rE2cKSAmkpM77TwqqJ+0OtT2vntE7lhgn1eY/ZzUHG4W5TTWy2cAoJVr5fbvX8aO
/g7fxylyt6JUqQz2L5OeqtRcbiH8AK3CYZK8bCTxEURiuZeCM8asqMzIwgzz9VPj
4cazlI4DLhnlmVC5OpRIiBxFDpTjArCvrxIHJluMaPLv0roq384cCnIKMvSbC11U
B0GtFIt5rx3hwN4bwqrf5eg82LwH7dskQZ40EP56J0vdnPSgW6wJrqqyeiE5/PLP
71Yn31bxUdLvdi6xJndpDOOS17QrXviajmxtmD57hwM4F+ilZcrk5OgN9xQq9Uks
5OWvRClVGxYqpEc6ORkxUu6XwrAYildCT69v/aKydLTVgou7Qs09Zllmz48MILuM
tGtw4C44GKv/IYSrONLrR69whTZuvHyGZYigaXIDGleKb9nlcw6lvfHSypGtsrYb
HBsA6sKWY3ySmaxw2qN52aiJr73t7a8uPexN9vyvRdybVoti6tOsbNRg7yjMggCe
iZJXayCPC4BIB4BUAzdnL2A/MYNWP75snVUZ78vN5Xwfh7op1rqCSIsX8pWeypAJ
34El8CRtiSb8ttsuFzCLY3hxftmPN2BqO3u1dD4cn57GMEHVzVQP5kpKJregGMAM
BgHfVZzGxPH7khEKYKVvLHDGUki2PufqsI5amR+Yf8oBygSCz1VbfsmOjbpTaO18
IVkHR3EGNjI+J6cbIQCpIZd3s8QHJ1LVAb9Fi1rkwGneozEDdTnI7U/C8IjGlE+s
pz1JfI4AyNXYtB26IHYQeQU3Shdc/kemU3jBv4NclMg2zvzvLhT8oPvh2noF4RQD
NecS3o9hT1aXdIDnackC/W0eXE2NepIsAZioF+zHvCDtmIkXq8zbED46EHyU8tYl
Y1+8k1eJkdLATXaupsm5EO7v8AE5AnLVWOrvdI+Sc3Hl5mtTYTS6m8psthBn8Djv
5d6a7cBDKHC9Yw5W09rQk/R38haRGSTERyPXnM3IjBd0RIPSeA9Wrx1tDAVgkYHS
A9c+W/fpBJVXWM0HUnSkfluafgPvhkXxBLrurGTMIEIWnQgbA1lM1M62AouFcXSL
ukphd5h/wIHhkkZhtq4VQwVoVqW5P22ZYXlvLG187IB8/ObBy1+xiVnfPTe55lbM
oLkjh3Gy8cKbCvRrshUwzqUiJD+Q+AU2zphZrdRmgL/O/FNSc/4wocyyFo+1p79t
tplgB95R2HQXs8O05UUZ3xNe1DQzEMGVqwUM85nkAEl0FoPbK1xKwR6r3ucRWmQr
kDsQQo911sWFhPyEWmvEArZSjzFbIPppT0qD+XVsaH+mKQM4KM5+Bwnzy950/Fl1
xqzNo0aak+fFo4LLbMCCcCovK3WA4zCUcnYkzF+SpaIoUauCXMpdrdU0mdkjMdPJ
4vncidQXg3bjG/besi/GjzoyhQZJIwDG1EYF3enaz4lebfpwHWAMjTOJD16XBYID
Br4jZ/jWNv0KYmCT2JJkCDN3r8YzqW6jyIsWOI5UTJnnI8N5Bqoxwl6k72ajZuZ2
1JRYBLS4kTln3u3itOxFZdF1NDqHE28nyErxVBQMr6QofTfQmF8DGjssaUUXSBTr
F0lRnbXI43nV2YlS7CY1r1JyYdzg7KL+vRoEqQnDT6hqR4WAPF1JIW+LLcNwtQhF
ZFo+tZi9/IpERgyql4w1XuOsFqSQaqgBIMLuhJbLlduu3Hw/WgGTfTDEYfoIqvzF
VTwDtQT9texhL4xJ6PMKApOgbPdCMl0kVUBZxjddMt+QtDet6aRsrwrEKBxpekL4
DRF4z6Rz+/p7BqdSrcc4P8UdcxuLikqXypghMAvQWN0HOZWJG3gO0mwkgiPYVsmV
34TNdOEJo9pCHSgLfeOq+sCHotdSKfTLnKotEaHEQUqg5NVMoX0qcgkcY6s/2KLf
9YW7g2ytV406YxwUI/xTlifovpt8d1QmQhK7zn6pA21AGU7V4Xps/JmzUa4G4s/Y
ofi+nB56xdJCvQc5R0s7C3GOHyBQ47aoOmu/CrZVYdDpsdZgVsGNHxV1Pb/oGQso
0PlvSWlUKanvcKA3dPbALwWFT46c+cYrgKZXpamw3F8tuNcDSj1tX7th87SLv8hU
YsrAOiU8mCg4gMmUG5OgnzlBTfBZoh20L7tO8TCZAaDzn6hSH9k5YWRg8AhIGnNf
0vg4UvF4gVTMOdbT05aqKpjVSywSKEWqn8w3n8e6WZ2D8LZ0RgL17xrWh8/YhW74
7eWhMf8OzXls2Tqy1BF2yqWIvDP9VoRJZ/Fh6ldivKq4SJmxmWcpEcHkzn3Gdd/l
/E5H1WSYyidoJsAH0CPRmt8VtmvGZmedET5P0db3Q9PcGM3Z2+DMw85qWaov5WfJ
U9WwFY+prpm4rkwUKjxr5yrVoPjV+FdmtYIRHXIr9EVyTEOgYrraT6rV7R6sYFX5
Zm3x+XG4j3OkEAr6wKnGHOmMBcx/9posZEO7VhfzVTxvdDhnH4720ZQXmi3LjdMM
oMfTZw+W9Pq400/Z8WAydFkUeHOeTuoF1P7wiLW8ykWzMZ4Xzd2tZQF3V7EzE8sr
xpkITJc9US3DNxcWXvWyK4mpNfmojuPexxMI/zrH6o3c7QJmEcYts+BmRo0casQG
8hljW7kTy50Q4yugEdBYasL0h8P3gPiMYfzDpTm2B+rhzpraMHVZSlVNwIxi73gU
4FISRfqZy0D6v/1m0yQnLx6K4ZRBZNGCVD/set2oodl2pp+ENW1USXAjhwelVCGi
qCHBj++v2agZX/7NS2Im+1jB/DkfCtOjKhAqJ4O+k0DBIwKlq9sZRFyNE4w1UkMe
0svN/8GSty1mk5/FgcyuzLPjytlQAht+hq/fzgvjKWOerCB+mqrtEy040R/w2iu6
2CtXpr66wwF0JjOO/7g8GY9lytswbuwWie7MInI6H9OouJVB3En2p/ZP58B5/piw
+WG2o8iO2N3Ma4eiKj2r/axsMbf47L95fvPiiT4ErhnrJddY9BzhDbmACcRUkfpB
lUu7LVHzDkATeCUI+jiZFOLdVtTv4QFXTWRBUXFNQK1AdeFsq8jYXz3SX8+4zpVW
/ku9uNYqt+lMOwyJ/6uAnoTjx26NVc56muWSI+CUBrApdVM9LrK3q2h3v2amG8Oz
BVzy/wWiXvyrfPYw8MJtgx/GvBFTHh8I2GOrMh38DM3kEAo8ZS6mvz3HrV22pYV6
NsQvRI1HG7MZc6r7v721rqYBdFBbBs+AStcx2J6/ZykXdM5Bm5wjGYnBcSkOsXbk
MIH75uaa6kcMRDRdg95BH++H3kjzLBlzSBo1TwVCHeg32DyDWZcBAe0QtOCQ32iG
2gvKb1JRUWgjhzLie7L9FH5gWLsNs7xo4RjpvGzHrLRpPgQi7XQpkJecNAZjaIvw
RdDyX0zXzIkaPKJebYXQCla1eTLNsMpCmJqGJDSU6M/7xNfXCTKgHoJok8sR29H8
dFm/9QSvjZMJb93X7CvJZy+4LM4/pOij0goHR7Z20U/SZbjFD/ou5q51KVXAeTMP
tekKFrVUhJiGy30H2gI/N2DwDOoda41f1IfddpkoOC2rZ7z28mIGMMXYSv9kqWcp
I0e8iLqZXEpq/pR0IWTpazRxTFzNRUWzTdIdc4dpdoaGe0da8Hsr1Q5/AZN5VlvP
E3Aay9FohIJQ9HLABRWmVyRqkIVcQTMiBPd3oQPnuLZR2d53tvPEZSIbTrBseqcY
/KSksBxNxAbB+xlwfb0uXlUuEl0HFVrTcfWYXCOiNkCS0BVieEFVRgghnlIcW3OC
m2JP62HmuJRFqzlLBicPsP4JYK0eXHHRikF6CNb3UqFvXumPw9yxcaWBqy/0Pu1b
qUoZ4C/iGFlXsoHr+eckBN0BTvtRcC7Rvqdm8HX6YFuVw4V0KhAxY9wyfytUJQd+
iXoObjcrjjDD1jABCQ8W7ijoozRLkso30OlOy3xe43TULbOAWrhi4kUewcK0DnXC
46zt1rDNkCePt+qzXKeyt3ZJ/tQThoslWScx4oBR53pJrd6AYvFVXED+t+yuj/b6
5k/7An82rrptcBEVLAWJ3pCpHakXsxK6fguJPAfgmmHQIXv4o5gQca08rR1vQomh
OXYGeDqi4gX6bpFN/1ilm3j47owlSt3BQGBF6CSBPxDgrXpMpV3pwAGPAAR9SYVv
zSCuj7kcP2+gOjSBpfrh0TIzL8uSX1z8c/pbyYdU/QrMxtBKl54001r0bCbWB9Ld
fF4MYYuPYKmigRCYlFwyBVZpCiOzOfqdCgnhDcZsokQayI1EIa6wYtTK1U2wJqrl
b76ncdLFkAg4crWxCFantXSl3S71bNF/hlm2y9iI5nDh8DFm8wLDuAks6LDApUDm
nSqj7DcJ/pqbFoozmq5r3ZQP+mDBqjVn3bVAsZQs98qVj9JIKnQNbkxput2DVaSj
2OaqlPbND39usR9hsNe6z9QBW18e8bESW+CqoIguYscz/trDO2CsPZigIk5jGxV6
bNXx513IHdOzSAVuUQKyUpUom3T4QlOTJush+TZwrf90VFi+bovcIzmmB9m9J7r1
7G+SZatIMTKkQZqjp+EuvUfsXHk1qL1GbIunvv1YqPhd/fRN/ayTHUWQuKW6NbtL
erSMCbQUyGClLTJFzySFxiXeK5nOnR0m6ftrxJ0+IFYXD0dJgpjDYJ2B5A7UE1/2
1EesKaIyhSA7aju3g05Xn9S35lzCSFO8nfnsayA+CKfyjTw1m1GfZfkGW64oYWZz
3x1nFYhYzxxjepb+k6Yhb0uEktN3m2163aXZSVmWT/gvqgHA1hl1BtNS7tXO5OLv
eoBakzrb6BE2mAiH/dJWu46n93eyiXRS2/x0bKiJTDW8xZpbkBxh1Jz9c4DOygbY
qMyOoh2qET2L0Ukfh8U1dccOzVKZCoyuNKzsOg9lu/6n2I3BS7K9f15FmzWxk5Ti
3vtHVJsBHDVbv0zn645hsHRMa+FcJdo8rVOm9bQIQ4ZZNIXxqvAD+s8V7i7IMTp1
9vbOx/ZbcbnCrRLZu35gowO0zwQzPmqjxrw2a4w9/ahuGkgw483vPGYWpC7Tke0+
NJg6L7UNea3Bo/E2FIv0kNF8QROjX6+tSZqhVXOsLNpvIQ1YjYeS+M/6cmFx5v09
WU43/hWClv+vnBvkXht/PLE8OkVK/UVLnVFUh43Qb7SUUbp+Z60oV68awNNphqgm
HLvlkxUEd1cy1fgyjA0Fzc1S7Cvrl9AFy7LzZGG25psRfqt2L0XtgRx7oI/dZ1bF
vngM6xWaU1VCG8rq2ZvmB7fIY7+JNPggktT3fJXm7Fhri4Kxn8+hYtaK60JXOC8D
t/QvY3WFISXOXVX+p5u8R+6ZD/PlRrpvPM9a+ra6ofFGBc+ZCyTBDSAuFUkOE2XL
1iiqr+JT77XbiwFLEALx5fe7YVM+Pt7g71SFNBuKZWetJITR5fX2zlyQWrJGZ9Q+
J7oSNWIWzzNrDcMv3/quEKCzOuQ9J3/aoZgtRornnMbDcpd6Mmn3FJC+nnvOxfA5
yHrp9l1RD/Owb4vVNnI2Q+NL+siJYDXp9Wkzuafl4wFER9e+RXKRhnJwj3fR35LB
0BQkHAf18oQnyEIDy/lTD8QaE68klOSp9qHzo9KItKv3y90MAJoc5gY/X+8e1+NS
Lkda0VlsX6MobBzwShBdd2xNwzpQYWcjgPzaosMagmRkNLJd4itPsF+LiF+7Iynb
CcH/KiJWrbbsn1GcQ5UWhoSAqBrgdz8zbNGlPdXbeFSbYW1J2bjAQmc1bhSDBsho
Gv374ax/CJKB54j/J1XSeXFqSi9V/ZsjsyC2HBjvfIHS6fcJB//EJHlJYrgXXefr
FAs9qrQ7nGLWOOv7cdgw9SvJkYw3Xxm8Izd39QtfhHvHHYxe/svEag+jWAKco7zr
A1UV/d/bmFBDigaOmkLHMp4/EEme4q84qTtUVEvz69bPgwkgRC5QR6+UwX16HXN2
4+ZZHvDe9erp3rof1tbFcs/wK3ZDw39xVB/X/pIRsyOWZlk4bfBdfU4gmhvt41XQ
ShmyPp/vNfVId2e5upZG2cT/rTJA93aHa2oDDN4/h+bIIBz0oqEMXfefcE7nm0pD
qgdmYszXDpahO/Pwo+KxQ5I2AgOebA+qgQvZjmlSSsbMuUg7c4tF8pkfqrhiItmu
896fNlnED/R8aA1qijYSY8hk4GGOJu5pOaPF0NhENO0uUy1L8Us2ag9AF7H2mclP
xZPyTmgSUY7/3AOxU4zEzM6CvsZh9kTcBNhe6we32FvvCS9jbHoFsavj9DGZperJ
6RRK+qNQJlCQxYmQJeCt9DkmBgA6ehTJdSLz5VUXoiIHQo7F/4KrnPvTWsWaSj8R
oSYSzX3C7mvX+MQYBrVNfqdO+XfjB9a5dLGpdEFT9L+n7mlRfDNbnaT8LC0P7VOj
Da13Ny/AZEqsEywqaE+lYPw0aj6jO/g1xWcO9qIEuwQO9q8zcKU7w96A1Kz1U0rc
FMZMqQEXjHLe3a5aO5AJIVGN+0XwX8+hP3zFuGaTxbdAd5PELwxaTKrBd112e/GY
P/r8rY5kAAuUVkL8czOb3BrMj3mJlWLCSVhJu+392xuVjRFQvvKsQ/Je/Uh7LSHJ
PzBk0iGa13fsMJ2bcL8Gu4y+XGVgGpJh/GBxHbG2yYnriL7MJWzy/JOhk58zDRUN
EBXm+z5ovZFgMKQuNtqaB8jyQQpNDCtCVQezj4Yl/Uy0GqM/vCEJUIN1EMUo77s/
l3QEnFylR+VSC9VmzQMG/8Np8Wa1jkdFbB1q8mazUb0ff9sIDg2ndk9Ddwmx67zA
lI46V2SgcmAvfSmsKt9IfWX3UGfUy3UAgfhJF4dmORjD0sS4DuWtkOMbMxaMAi3w
PQI5UmgL6Ozh7YB3IKBL8eEdYOxbdlm2W6UnT9hpzDuQ6W0lVuFfcc1ewRG5A5qs
Z7kO2H+NlNxmDOh2S2dS0D3sCZXiDses9fV4b7o+s9NtBJm8+rYkVt7VOsP1vJmI
GlNkSDuib/hzkobYPP3XgQillGVzjlJ2LMOMU83Pc0kacaJOogn/9CgLOb5BpK65
XNIJoRg3WcTXNv7djcKQiSY/s4Z/EMI/09qZpNX2UMm644wJAQtRdHkf3BcNAneK
IXBXXZ7ukGZjKdtP2ge/IQKeyS6LZxiK9/Nhc5AdLfVtAr2D4ynWq8PPNvjD4V8S
EVNEc2fSA3ua0yTunqYs5hS1jaYffTbPwxJo3TzA4UtsNPDSmnVI4vvMMBg09Iuq
8faB5iS60IIH+Nxq1BwsoqpFHKrlX/T0yFqlHEpyLsWhcF+cp3Yis698MmV9XSsV
QAyw5BV7istypF+g6UmD1n1yPldNoA53mfRj5nLiNj42BvzDxTYIPDdKOBF6R6GH
qwPqqM//iBbMkCpBAXkbO8J88wF0HhshekxZ3e8hewDdtKNcFzAFm/jxuD9AojP4
/plmX8IXEmePJznaILOHQb6JjsFXlaGc9gWHyNN0M6u9++WPsYu/TJzCji3c8GCE
9Q7YB1fptxL8rQLDw1obk5m7C80mArave83Q5vkf5gKC0s4PPu22bqLibVLB+2Eo
eNsTJo04YgVvkJXcxBT1Yj0PiGxgyiOAvXGSCS0bxRrkTFvml7VCnEhn9RFm/MAi
DrgH7X6rBkxrobvvOs/ORVhCcWSK41LVnHbvx3OnPfzbDW4NDCmuIEhynTznfdpm
PfXmpe6mN1fAl6X8SiH+qUovqgKQ8Ngb55A0ZcZj9jc2NxD5Hbs0toMhDMdk9OG9
+9A5Yah8VBuDIE9KUvlArA2IJk5Knvj42P9kax3iYnqZ8omwGhP+DRHAxfdQeYrs
9T38ljnU+rd78y+6Wt/RJsz8nO2q5fiGxaU1N5fAMeMOjABJr3VF+HxULdwpxsd+
uqXZ7A4CAANI4LFjmBO3CPhLSntQIKAJodw6hmdXqbK/YXEgGiMJw9Bvael2otpa
Nr4xQYOIDP3fkkrg0IkH+kU3vWKGdGTUZiY1y+jI9i386SGE3olqxDNB5ENwtdwb
IRoIGAGn801v3dClTQ5JCVYXRZTCObfKFSXIKPVnQ2AiUtICMZMXYtxB8f91EshI
athh+ygqqNGeKtb7wV5fjVrq13pnRm7H81U59HX4VU+vzChWxugHfmWCwFG7uvmd
zfdBYW2Q6EDJBsZFDoyarer3ac8CQMVplRwXMMnGnXdo393cNz8XVpahWymLEy+E
3rLWcS5qWNq3VZKo+ro7kGdSR/Fvh+3tkQYmm6iWSW9KPr/Z7zG7JRJgqwAQxUgA
69tC0FFTvEDyt57dKnXV9q7cF+DvBIk+vF9OjmADXgAXFcdK41rOCUyJXivbO/3U
BKtlGqOK45mjlhxjsecstinkNj5X0sX9uH9tugOyV1/gOQ4O/+NyFjM2eVW8KNh/
rXDJSqnPePyD84AN/85AgZbB6ZM8tDCZ/L45vARujDRXndYdyCrwnPkpRlxSvlHp
ajLgbzChUEFaY9cKmF+nWoDk2TVFM8q0jay7NbV6sc9/Wc3xesYJy4dwgbiPH9BQ
pPSrvectRuaaQD34eOCAHdQsfngDaOxtDBKOceQk2YL9l6D67By0ap3SLPJ2DjHE
ZRn8JL4uOr17K9MX/a0nMVTatnahM2LZ8I2OL4IMYUZ7c0N/kI2LU4bkdkuAtFcV
qzP6lvOfzgWYqtFrizRBpNgFY1862j+Ehw7M2OSfsMLts2gimtkVEVgpXJgHxQCQ
kXFhOPcNjgLJEdMiaLOiQmOpqgVN+43+tPdBcynOs9XstvO+Hthyned0O/AZbWax
3s57x79tAGosUbdOhLWIt51rYg+GCh1eMVhpzutttMdGqkf9W0aW99Jky4gzmDMp
P1P4aElaawmI5alAGuZh8xZ8X6T9PUTtcRJ4u/fZycHyThEC1+dGHG8jLf0zHy6N
LngjKciEH0ERGOMAdXnmQpglpagdTh7W96yR4he9H6AaUS5kwjcFdBRNxgQb36rA
raM7Kc9HmHQofnUwcf4vbi8Yz9zL4+P7kVSc3sAgpn3ZVPHMlXQKPLT8yE9rJTpb
M/wmf+uqYPElmA2SJHVN6TJwEI6/aoy+/9dZGKN86paZ2mcn0Jkjgn4sQXaSbDfB
ZckrH/VPl65zhVXugIMYPLbgYVR3anmMcqysM7kHiT3d2bVSqsJQif7qGo/BJg3b
RuVZ5FZkPiRWE9Cv2WlfpNsE6DMel6f5tGvQQxYE1e6WaaynwUO5HSzQgIfKmepZ
QZhp3W+r3eEGPKsV2r5vfP0VQNeR9N8cd35LxJWqIClD/JdKcYo6jqmh0XdZIEel
/oO+gN2ZLnI52TOE5LDdLSAelsfyAStq8BTVyQzIDG1XV+BIq0fXrOsHyhKHpHaW
aniMIHxpBCIxT+6FTvuXUU1zEbyyBA9c+2HxIfR7WVhi15tBDzuhlhQQIhcGiwBO
jFg5de7Tt1iF6zZA+6pNGi6BqqPgeFKlK6LC/EUnZ1Y0m2bbk2Ss9dnNWRrSN43J
57QrMQuGeqLSoxWZonR6gJ5UJ+zYGmEFOqkLHtvZMS0OSnmrcrHPp7pXax9/4Bof
8PigmFGUTlXAHBL/gWL4sPtjLgyr55ROAfeMW+PjftCEMe2iNWJ96DH9vTtc2i4H
IzyQnREG/UlB/x3NDIgoSouxRLRNprxADq043Ay6WSM+GdBNff5z4CyeafgLgc0O
Q3cGKflc5jsbLaZpm83O8MHr3rV2TUUgxLYLX2XRKPOHujMM/EyODZ+nx9SfC+IB
LBKf0Z3A/fQb0K1+j0iHAI/mXCkd5YGT1S0ZnXVoEp9x7hY7QEsuSl3Pyh3kR3a0
PYf4fYq9Ga/loc7tY1jrI5xxWJh5SglkUKeYb2YgQLnbv9Ax2NGnfAn/5L/e8DlK
IrvXriprlE42Un4yhf3n5ri1ULiNGjOiu+SzjGTLK0wnzXrl5mDEcZynKt/661Mj
fqOoN8o+7bt4HNFEetgunHufDh4LfV5KpVNYELccwO6yGlAzKzLj3KR2dBV1HCjA
NWuwYIAmdtQtpAoHo4q/QICo3Q/ptuiWdL+PaxU8nEA+rdws2bdQ4F+ox/KWXCZV
VSAwdX8JD8erSgRW7Sn6BlMZrgvxpFMHQFmkSVjqbFnbJu3D8H+zkC2FwQLvzmQ6
fcUBym/ZMlT3XxF7BptYZnM5uEeMSKw730hNXpYmduNI4ujbwbhQlnNuL5n5s5hK
Q4MpMfAFF7TIMUSEMc3ZoRta+q3QM6d2o4HkPuESBVa6gdQGDUih2QdaLOa8616r
qs0OPPuNhTqYNaFXFaJzYAzTvH4eDflJcYBSWxdJxbIkR5nYHh8RwCHTr1u0KC0X
GiuhIBNkUgo6Pdb0BQTRlz3z9RkZ+VyGQujig5QLGDGFrMxCJmQ5JVY9veF4XALE
QbDAS7XsWooQ8ZKaenbH4ZFfaZt+L2GOe1S72ppATHNn7qbMeD4Zwrpc3hf5YPSW
32AGZ6v2T4qORB8r5lHSA7THAOPomLrUOc2wQb1XoSGu3rLmte4AWqUacE2Jeebi
pYw9kBvNnwVXsRAwfCRz6MCkTTmb8z1D/Ue1vrDc+dA7KfgK7v0mByGjLz0m5OMu
42WwEUnvr5jZ4OANhlaChL86JUvP7gqB1XG6Hbuiun6i5UlUOtvXunltxv5osW83
Qe0AaXrjxLngOzaqVqQgNA/m/urBmeF3NbdGyC2AmRmkLFv7Jz/B2NL3e9GIdeus
T1720vy14zrFwInwpPT9WE9BoaAI9UCumuZxrCSM+mb6DBlodtwd9I0P7gSZ2oNW
1Cn2aY4+nuwy40XFrlCsViOuSVSSFlZp7jGCn0Tud2op72KpNDFwwHu5ZjsODaWC
BsEZ6VDWmkzc8iY9SezHSHRUenEjsy0UR0phhPfwzRRRk7X0BErTlILBzN6n9mVF
fKbuLy2UMP4L8vCHaZOHQWE/1XmgrhMzLtBifTjexTbbJPvUSYfExFuP8HHmT/Bj
A0QJkyNDc8HUp1eRAiDAtHijcCas7Wl5ar0dXqTSSexXGi3Mk67ab51YMjnSdpxj
EOSk5mHySqpSbux4w9Kohp9OLRetQnUcT4oVwmXaCPSnZoro+Emcqzw4nqs1BPDt
1lsMu5qpxNKduULinFKFtgvC5LbzSWEOmBNyOtSpP8neaMg8wt2Nfe4kil75eIxk
t9ebqq49waO9nU1K+8s6WtltmdaZtG/Y9MhuSNEa2D+SD1PhO8C4owuF451maDHJ
ysWdm28WaUZl+QeOXpQY6S+J2FPc07g3OQ9XwicEFI0G+FmPIQNmKKvVFldHTiAP
tpMF9aJ2zGy9y19DKkQSRBSl6ykMr3Vkn5tLmHC8hbsFD0uuz8HYN+N+gG2Ryewb
m9jGOeEnqnwnDY40r6a9XZPg6Gm9P+URbVIg7PufPOJnkS/mYAYAgSuBBq90kDtg
c7Ug2/QuDAJ/LJfUq2ck6Z3vIF4Ip5ipdVGJOYqxGnUmSNfWiDBHdMxciNd11N6v
Ck5RrohY0GplaR65L4XYSU89qOLw53T0KBgnDaV6oKF0R8LDSnqrPuKJ/w/lzdMb
PEQPPpoU95GAunleHGhkSBlRux5S8NV9drxpnBnX3mPySARAj/AoAs1Iso5dHA9g
biK3FyVIPa3YyAz0sd/pU7Y+xBb+r7xxJ3Mx2FhIQQshe4wjXXu1cobEwsvCQWfP
H1asAL5NkGsaFuzN1pYyZn18tA/0P797xZhQG7nVvzTn32/YubR3P4ZWzW9uOEhk
CurcUJl+k1J6BwEuMon4Qm/0xytuGbQoja1JskA2CxbaE4jmiDgamCy1i2csbHit
GSFSolJ360AjRC+05IhNhAUB/2cJtwI3ejziydiMgUfj995vd3i3baQwL/A9Y9nB
yorCetjcGm0mWZk7ZFtRv9cAXbhgsNeOQWdJPdVnc9HzCGHC06jK2TazuW2b3koc
w2UBehWXvE/Ao5lBevjCnEsl8q/79DxBbl1vnjjs7DrEHh5hZdSLW3jpyF21ng+a
0M3qynr9iTgG2XaA0hHA6gGyKBSR8OdhyZBCqclEwEcYXxOAkFr6pHWeBQYYJ+H6
aYKDtAThsCX9jsLyG3MNWI+lI7e7Xi/aO508vw5l8ItOngzQ5XKWJRtq6CUe/BoC
+xr2lrIwEZgmqTX5+MBRJjevJEev6gZ0Z47s9VHE9AMz7EKdmdsVESb6mVRSyqQN
OxaDiIQqdM/E/d+yprZBR/Fu4fVXSaVyp7RrsxdFXZ/BabQaFYGc/Ugtf13MA8bX
7tG9BREHW73cJP00AHY9BXSo0yg1q1vlQjhsx+F7hYsCVj5ORh5GlzcmWYxBHW+l
KvatK58iWVtYwcdJeAE9kfBTkZ6YMdvSaC0htB/V9Da8ZDQn8b2/9Ct0osteMzQf
/Jc/jDgknE4WgrteEgzlenZwpQ19iEbv9yducUsJRDTIklK3Cp2AkIM19acEQEOp
rE1MXmp15k2xhQT+gyn0Q+jbcd3EdWV1KbthlHXWkt68QKq9NvBEF8pEnowQT+Tz
7nNk33FxP+duEkM0prm6hlAzyHJVKRghOFh8qttGNhILAL5lu8guDC34O5K/Nlqb
YVK2Uuc+zpZY6KwPsfJTXj7VsrvLpFXOeGNKU/0uBg7zhOdzF739TQaiR4heb6MB
vmmbZ65n1SuSEg2mtaly+hMgCj4EArgYpKGv+/W4BovHoCurSsjsUgBtjM0pOjqz
hQ83H8LAzD5D9aX24EtpPOS4O/5aeJKpMYgy6PorGxy+KeqtMr73FnobG04JuEpu
5+bWkTAwceM6iYNhdhvz+D3kkllfY4e4p2W8tE5ti+r9Xx/r2DgLtiPNkJ4Q3L0G
Al7dzQvg/Px40WgKYQUZHE82oVfTfx3+fUdNSNlUTsQ/kZ9HMrDBF5KzbMgvkwzW
f1ZsxfZP1pxZki2FTPzNPNz3Yo6sGfFrOWX2+V1fAqSO3aoY5hZjrHtbb8H/eVoi
SV+8KgOEQ6e7vEo8GHBz1F7qwJP2hDABPrPLUijk56c79GSa8b8exdhY9OnkAgVU
HmhOC9D4vhx/rVW51MVplRB/8TQgHf4bVZ9WQW1HKHuvTC2QRaRIdkFmc31A8+VN
or86QJkVh2dAVhcL7+M/BccKoXB94XPa6RCI0OrEFWe1p7BlDyvk1hVCMJF1a0Xw
rOG4DHqsyksx/ECbj85ouF2rPc7gGq01W7si/G3cBvHDqS9lbcmVz1w3fU8GyxIR
2bIP0pHklW1KTbGUVgBT+D/dmNLzPvtcp5ithhUJF8hwF7X9kyHt+5tcX/yQjJDC
07jcm3IrIhdkUUWLsiBXjqbgi++PuCFurrN1jpGtASB3YqUnWCCQY3uwuv0zULca
cbCFw8P7/fq53JK7nxSIRbvDDzRSxv3prl9GUHpR35QxE6VJAFde3XYbHROqWOsv
tAH2VIhyzyJpckT9B3ExG6n6wIaHeyB/q1OKtNYw7l80HbOzssM1hFVDDVsGQeO+
skQlWfNmzwCUjBgKrw13Oc77hodV/YTonAtwRwudSo+hwHdxXMnqxDOfEiF5QHRr
0fB9pFO4LRhUQ/szs0Mf2Eb8g8mx09bPO8umUXjZCy8cSXzp/Hh5qL31fFBLH972
x3biW90keGHvHfhSCOs5rfiRRkeE1UN/HzhDoAalgAf/iiHXvDe8ssOW52CBWSK/
WDUzTFu/NkiTnoZusbIksyyHebMp4Gua/snpg0EGwVEsq1NOF2rpFT+rXS6TX3H0
Azaj1xnbr1Yb1kGyoEi4DvGJoKczV4CUU8PZhhxmacQ89MSgmMK1WT3lYgnJos+X
v86LNCqHYVOJtrzXzK0JVhvHeeDIcC4f6yXY5r+NN7ff42jBT3Rt+0qhII/bsCyJ
0g6GbWk3MpJ5gHFQtw4WXex4N47FnT7mykTg3e6M7Cztt3TP+oLqKvby83Lft30j
OxK0HXlKzS0bjvwfFqtUcGAEN+U/0G0IDLrjl3nT0eGb+tQJXNHtE44UFas40hNo
oqV0gfyjLQEE9e5OjuJYtw59C8hnKR6900VQsLzh2p8m1vbuoRYi/8nY/ORQc9Xa
ECEGThESExIuPHcq0cGcjSXk1Vgxy8nmv0zcOMzoQDj7NdvtyB266MnLsxT9wZZd
5fViWoaqEgwfn8zMVUBUta439ooG4Se6ZjElWrnq+nrw3kZX5fYADnCoCGHi8QTS
6DAV616SPQ5t22oPZBneGeeAq/wmfu5lm8MTsmiF+GuyoEwh1adLLs7l5uhZGNKM
nVwLVw3mELr3yeh6GpXjxo119baUZNJhbfqQjWtuCg769sR5nj8FbgsQsydgyJ7i
UT2u3dtCabLWHilLHgweM3vsTj14gCE6CjZ5L+bpV8/aPqRcBC3DysqZ5BJ7KDJJ
686Ja+B4qVqDGNjc2jPxiZdetoBRvj5ppSm0Hvx7tN3/JIO7WS1nBxeNNHYkW2Q0
Yd+YEjF8Z6VBCC/QNMvtJcC2GwGOnS+/C7h1ivAcaksUnApbFcQLr1r+hd59OD95
R38rqc2LqyzIyXtesWnoJRkgTbmK/fDHbXRfS2YIxHV2/yH+orit1WIIF72w2vkf
zTc5/Xz6Y/71oqlj2LBlGBJM5FdGeoyoYdmk7xhSkmuugNlQynZz4s/fsIghBtAh
NsI7nyOpCBBLYkLddOhgJLFREw6xNO6FvV7NZAbCS9Cl7xmgd10D9VqLsV9U8AnS
PxFBdkihalZv5E7N/uVesadAFpfrGqtotStYyIXU92VUsmdQyqEIH8B1cwMqvBpT
6onanJvzbpVstrjd4XL5aP3i4MwT2/B4CtPbCGCIeenWqdDvN734XB12Skt7L8V0
MVo9OU06Ja/JoiSUf4s6/l2pCvizXDprakHB2UDX30LBQMFoh0FGlCst+VcLS1Ta
xQJqZeDulq4W3r6i4Vp7z+QYBQNC+cmmrRV8SBlCnEBnLDxcizUgzJG1HYS2E++Q
vdhi766Oxd97IknXwBfwKWO/guxLUKMNMJIYDnh9twuvsdhk+Ye765w8MakSRnxb
uf+q/lq/EnEsEErcN5AFRsq4qm79kYzf+A8lplSy0Ms7IzsOWPvbO3HE8gMYi7Ss
JygbcRh/NkEowEmsgreXuSm80PF3yuHBrP2GJn2IDIpPVbWlx0ryJl8JAOvqILbR
6zLD0B05Rlkorf7FPfI6Us9L6ancNCu/Tuw8JZxDd31ir+6BoQR1U6CjZy+tm0RA
LGZ2s9DLRUpochIVjsxWj7nU0tw5djMzP1yVFBT5auq5s8H0jHwUvRuBrrVQEpXn
DHsYPpHrbPHEQXAk5l1Qr3KdZFtzCBTQ7U5mHBoA+B1AagZ9uFFIEsVkizxZq4H2
KR4fMSOUgiV9xCCVyPwrUr2z3rQZcMOeJR+CHXl0NZRT7WEsmG5ZaMdW0SfEjKai
tZLV/oTg/BoCtjM7FpDrNBWqUqYDrL4MYnrmRCjByVjIRrujkJCkcQfXcsi5a0q5
9HtfsvJ6rs3QTjfO8TxK3x4QJcOQ3T5SzyGlYL28EhbG/i4yzHs4a+wkmn6Mydyz
a18Xs25EnUigRHQVMf5h4gkF3o6arRUJB8rIf1sHFAMpUF8Xkw71vEpqIDnSxRYX
iht09zI865KIZrqP9hkLcAQGb24TKgQV9xM/6p1f7fBRW5v2s7HRBFyq+IFIZICg
myuyj7WPEbI1YqV6NWCyF/5GXxvP3kBseO2EQZXwuN61IpLsuJ6GEuFMDb48DcEr
0hdt6eZLGXCi+HOlfYyHR/CJ+THUBQMzzbaULkG2FKJznADUFkQUgstFbky85W9E
qFxFmghBggiBRP7zEsmjS5Bk2wZSloKRrBC9hWEaraZVhDim4g2AYdZHGMuFiE33
UInAjxeZUgaWKVt/6B8EXPePYcA0kHXjpGTDZL3FCiG9JRZtoWJ61lD/F6gjz18B
kznMEczoyGcHCM50CjyFQqVmL4xS/0IIIGkQIbQMLngkCMbb49FwqcasPbTP11G3
qe1h8LrVE22FucBDWbeVP0aczEO+IJavmOpKAtpgypDJuuJFjZC2sOuamedaHctj
2OPe7jsT/80sCzLdKMru58Z8SDiMzT4y2K4M1vxaQDBQvW0PgF3GSt9RMQ5aoKM4
qxY0mKGsF9lW8G0KkPIF5l+Z+4k7z4RkVgwXQJUl/WSW90qfq4GqDV4icV/1nJ0i
A8CuGirA+wKWsMSKg+oKL5X8LXsqvSvrIujm6l3wfadZfmkVgZi6YNAZ5eyIk9AW
amlVuZIkdtvMH259NqHQimP0sd/8UQsQsej0qmCsYH9yfYgrc6hX7upotrQoWpnP
faEoyOr9q1BNxNZzQvesGOiDQ86UuQmRvSOEGJ0EyCzqnuqqisT3/AXMZmLZHvqF
vKCa7/bAMIdlPvQtkY7T+cibDfNYAJ6VODOcSSePIy+rsln+I/LMhrp8ajbeEFSp
I5GqrwX7gyi6P++iVeSlPsDe4XvUAKsJPmlNgNQZyvZ28Q0UMjugji/xQYjZgtIO
eqA7bgdPs4tjx4m+3NppQq5hAoESmL4PKwIqCM9NzPOVv4ak7v0TvoUeUzPOjgLU
7cUqooI4fYjBnRgEblVR2Dp7FGh5Rfg7UgzneZcp6cg7qFwJJJYDs3D/sR/Y52DF
4sKd4bikpULAIS/bW+fxLynGrvjLXOFyj6LC6zbkA8FQpS4mSQxwo7TgBbYCzgWo
lZ9deCPEo80YnxZzux8e//ETPNSK/KGoixB3sISEgpgkgYCno4tjfg6DKRaO5zwX
5LEZ9RYKs5j2sPJVTPRUD/4utwvRtVezoeadvkKF2fyPcdIXxBlUlhqBbdYCRGO6
sXZitqDoitb3r/Md+he48XPCJrgWWuwc2npJ+v31TDdSAqECJy1HAEy4nw47KM0B
bE/stJ3jMPAMhQXPG1fKbOnPO/QGFzscR3vtq8KRNCSG5qv5IdG6vpR3pYW0mSLR
Bz5WPq6IBS71ITJjJiIPWDPlRAwE1gYvBiVYYjkCn07SXo9cLqm2Wvt4wvyaB3Qu
f2HhU98XmdgCYWoda/x0VSPu2dcw6edv6W/YyxJKVYcTMOwcwnI8LaK2d6Kl/frW
AXY+mJmQcZKaeC1qwfN0pUS45luUiBcuNJdi5N8tNl55Zw3740Vh5YXoIOgxZ+KZ
V85sVpvDl/rSPNtmISBo9mWgGEqw+UooIur6jAY3sEHWg1rD9Ebi2MBhUDMGrlvo
BELNy8c5VL3g5M+DiPmIj7TRxhAYcldiXY46lFMlyVsmhyQD8FqYti6+5rMTvQ//
97nEuvSrbHbxiafJ/KXYjzfs5aLM8/uUD48HN6EFeNmEaPX5nh/1kAAvv7LkN6gG
vAFEkrxN2kdjBsduOdFO4lWIFo0gmdIn2ilaeUKAuzy/MJ9Rk/JXuQCIKKbsqOXr
ixJOAFGwbQwmK8gKJnQw9lKp3kytGUueoYlTTKGyFiHDOiHZxBTCZSLtVItXm7bc
x0zHk1+Egx9nrpcCR1ix/TSO0CF2tYql1b8e1qmNyTl63MiISS4d1fQNqnPDABBG
K9mhk987dcRNh/pcoLv6m2M4FooWf1c0aLBMotTg1Ii4P6XBZe0W5E+flj0utEXz
orSzsXsxm9tLUfKsrACQsM85e+OFk0uuCh/Jrn274Jv9vllcP7h4sy99hk7GzioH
Zq3waTX0nEdVulYQ1KVK2i9gySYe+YwC+aTuvi8KJwKbSUdsWqnHjpEh/q609omD
cBErt3kNkGu+HXX5CdKOTyzTQ5N5RxUNkBCDKLNaf4ya8iJtHnHrqTxpzn8IpXMZ
sL60cwh/73pJTTHaq/Gy4iX/swuYsJnvsCck4ZbLQsYSLtjvMnf4qVvZBJ+3CarZ
rTj87zyFdoTir1tigH/eqyczGS5NvRUOdjlwI9rLNaveyXyM7VEyc6XC628IC8oR
DhLc++AsYbeRntaEFH7WebWtXs4JAAvak9GJnuJqg39ChU85S5kqyJRcvzfd6M5F
wvt1wHjNT/c0mmObpGnPTaHLj56IH8bLLn7zT/kga6pKK1csCIweK+R1+cNgJatI
klQP3mo3CJ2SbzQ8871JIvfQZNExHWNB+IV8qASTbW5ZhqzZxHK0jRNcO+1Wr78c
vFOW3G0Y9gpElU86ISAk92lthGU1oKh494QR80kSu5UZ73WfG2tEzY+v9pnO27oI
eo/D38Sw2JDkWhM4r4e978KNfEaDpKGWK+O8snAtmM4Z2i1EyLaHG4WCSGbdDXXa
1XxnimgUSHUZk5wWhQ/5Bz0wUlIYH9nmaHAGqqTbwlra8KxGsTNUkHFhrusKD33o
Om/MbxvzpoGUp48/IXJReQQtdO57uoookmb76uyFpRLdIYttBer8zIX8sUxL5Llh
7zm20klB6HY+1ae3JgAJcb/bZdDFIzSqTEy/tivbZGBO9CRNGGpzpdtfe6by6cVp
FwvPAta+RPnNOq12RjGSF0mM/4/ZavIicOVQ+JeiJQe+ea5w6d4zzg/iUxqudnEM
wrBVrSh68sUaZVXVc1rRJACcB6slcoUfqPxJDfFJ2es1fSIEjYJbZmIl0hUjCwm6
Je37HIwv8NpzE1+Deut5KrXeWT95cYvPO4XqY6O1qNlUOurSvyJdHTqGGjN1T64F
HI8KlOUHtqYbmfGhxr1MXIuQ1NvKGIVl5Rrj8vAim4l6erJ1c/nXBWW04BLJvdDE
nKyJsda2egI6NQV1fJHDMWnmOkFZ1EmsisRjVjTzElI7vNO0o0n78wRjlI6qQnOK
5HiGCNguX43OOGVgVDU4TMcKQcCZcpanphYLF4Dd81HycIqLHSeMg552qzf/rxgp
HIP/HItCepY3RIknfveInjW0mlM0OGajD1LSvaRgO+XQXXt1Ogo9/OvUjFKysTVy
KAMAJ9hB+JleWD7dVbTUY+3RH2a5FPMcRfdMJaJA+wxCjynTQjhHLe5Sj4l0CzmU
aLgfU+nxPGjS+vIoNFwEmJEBlpczG/ou+7dWjb4N8q6ixdbwYcjDQiCWV/iVngUC
c2i+J9O0TDUX0fxKOA3WBpd4u7a+E+BJ0iaVhFL06so6oBiqH5mlNQh6ym4t8O7P
b7tRDsgoLHel2Fp2PYpnjpqcsX2m4kBTL8E9YrUuAehrPFQej2wsGyvHNiRL3Zul
oDiVMPXIZ5O5penKs54iq24kzs/s/c6Kd0xmPiZjmxlA41b+qT65usjBZIjD9ru6
SaCD6Tjy6g3RZ3NXab5kKPqF79htZlnUKDHaR1/QnOLmWPkQosNgKh1156Tx+kx1
XDojGFn2monLj1XyKAo9lCvTCtVdr20lo0w9wKwtjNfCRS+0VGa8aj9tx0sOD2r+
adZZPmEsZLnHHqaKl8MlXnh4gNP0ilYOuFMMnjX7zkarJ6c+6lBuGZEczVymRLiZ
OCECKrPankE6y/UvmzjcTGNY0UXGY8DmQNDaL1fvKM9MU6g0soCtjRWCk8M+H11k
2uuVkDFzyHVgkbeDov1ktaU44lIohDQxMKPClT3JvnmkKrTZb2n+2EqSSQigB1uz
ir6P1Vy6vyF5W20qY2pkdbt15r3Mom6Y84EHHkg1pYNlGAyvhwX6JecP1If64EJl
pBo9m/I83K2UUmH5yVpAt7EzUfZXWDFh7+EjmWvfCYWfN5PIamBNRPJu6Xl/uwEB
629YYjHahjE6yLrjd78sEtux9Zpp9WgoKGXnzNRbR8SZCZo5R7VCNATjoa+3JD7u
gudnE7ZgNroYyM38GetyeaZf/J1TzusyitvmuP5pcgVQLJm68jS1GpAc42RQ1por
nbOt2sSXinudhzHKHw6w3MoolIsS39Oe1lLz2D438poaWyOPlohxRFF6oIp9PSGg
ZBtYoDpQ0h2/FsY+EbrbJoHw48nhcLcFeYy84rEyEFJkrNzYE1jwOmXPbyf3+Tqs
V8Mz3Jbili/ES67TsM7cIpUkhIiwXRZAICJ6lCsRq1OEnvDTYE0CBS3kPWhTQ6Hj
kmW1H8l3pMxuM4x4ktJ7uBJBBOGNBuWeR2TCV+4ZxwwfeMBZniBuEQBp3gajA9RQ
K/1pHBGIv9YoBF535vid1p0XEyimh6kq1lBluEG021UzYJrwF3Qtq30Wsg6WoQx0
GNv8zYaDE9KW/vdR8p7bkZHMT+5zz9yoHJRh9058wfE3NZfYd+GkBuIpC31QZmKj
fayEvGTBpDKXFdxTs0D1FAM4MSEBW+zuPal1833hRMkDh+WCP6YsIxCjjYZjP3jF
4VPyYwD8YVnO7qTHkESy9KbynKKHQkRVjIAn3TrZFc7o1O1xGY346P70qiJFTVqx
nkT8KCmM5S9jqYGJcIjKjtxNRec/wBQy4JTd3gmGBDb9vtl5VFQQ0P4KurDePGh5
GlbP6p53ucZNGnL3pOr+uHXsDwwdH9WMqqmwG60y7Rdb2bsji/K6xd+VZ7L8Yb8C
h4np/1VsOZZCFd/FPh+owlRuIhoAmoQbCd+HjkDJksL6ouyJB4FGAxbwKao7Vy4l
FUn8aaepkiy5qBddUDOLVfe9KlLEcvYwTFQn4rsNHo8sECHW3iN/TGdX91P5dD7J
BQGq0a0DPdsIfuGOMg63kdeLFKItPwq8H4JnH73LEVIyh9W41sLi64YqqZWF56xC
VOpugyPqDFG+niNNpcFRXC6/6uwz/TWg/PAycl5MFNzegSsTeELdruXG8Kw/jTcw
F/9C6szH4N11F7BkfoquYThEX0BASouWUCKuzR6tFNF8fGfRXWnc+ADxdDf6TW6F
KC3BnZl7SAeHEPI14ZO1UUQoPzE+JV6OTzyQ3XfE1zcWl13oaV/FdvNGT0qyof39
1hUhAi0Gdc1csXpar0bYYn1uy9g1Ebw7/ckWb5evKuRYnVBykN+szOYJe6vzBrGP
qBgEn9xkc0Olu+FiFyk0X4dBdok/2TcYbN4McgSJl8hdox1uXkB41LeuCg42nAxJ
rX7zAN4bAocx8y1HODc8IN3RYfVtATu5Rxu3fV9jjgno7VJSJdVAZxkNTxUKAm0+
ZJ6ThaVbFVEmLMRdH7/46+3LapaJt7bHorRilpPDKoPW1rTB3cEA6rOQp2Fl8W1F
WmXf/LlNyG4JYGK0Ak8NjuX/aAGyoh95l8sNI7DTtsRQiRRFncWdzYaXSfqhee4v
7IzNYC+GvZzN7woVNpDb8cRQQBYOIRvI4C3krlvR4YLtOuiYDgmZTHRLNdfoQmYY
Fy2nIfcKi5/zxGcbGi6aePqbB1H7T3CYe493HrUFNqUMFvOLgam4IJaQ2DkkyisY
grIdr+yanS9vewDzAMTBwpHmkavDApXr3KRYm5+lu5R3w0WXlsfiW5hFRJ7kE9Rn
cSVD0Ei+hHABDR4OIAm+er6VsbpSiBSwG7XCdFoHqFO9S+aBEhE7tmXF5aSN5vMl
H8hFudA5olaaKOonMxSz14V43cNx2RqeP9QBLZuZF+c6s2a71Lm8GFAU0IP3YTyU
Wxiw7MyFXR40XzeIFB7mOzD9iZqygWinozCWYBeM7q8wvR1Kr02MRCnD3wkuDhPt
icmRcz3XplEE+QkZfq//pefgHD0hd6CUy+wMN531mE9uAH9f96W68P2R+ZT2fwbj
yz3nupDvjq7PxiK6qvHvqaI2PL/0RhP9SymwHuut3gW53jVFxKdX3JRP4YAUuZKJ
ObQX//glLfemYwZe2HDE6ZJi9LDIs7MjTKd1sE33lVtAWQkokMfgPaRq4cXAkwf7
gW1cFGmpU6wztOurCu/sg1eO3tekdDwGAr1uxWRRMP/YEpvbumqE/cSLj7phTzXM
yuhnLh4MQs+wMOkc0ntmClcNxJYOeIG4Mo9Ca/+zxrFMVa2787/2UuHvy/8DLK9F
8PZGasD58RaaQ/yUxhl6LiFXgnlcfPg39bwym0hEu43gtpEahenc19yKDsfqReGK
chX9i+6a8jj+Y/R8g2sSTi59yE5yiyfJEd9YoT9jzWjKsSZI5awGjugNaRvwvauH
h+r7t/yJ/HOqeIlqIfb/5IotTDJAoHtgPSt+tM8TQtY1xjDGXIYI851issgBzFAT
6zsvxC9DnWI63JyIGpuXGMyscnNef54mfqvCmzzdQC08DIeZyzpqHsx4JhZ3W15O
XMZcG8gqgnpekC6CLdEMeC4d1h9bLnCjwxyGaRh6sbiSTytYjMLI0mwCQS6M/Z0b
I5O9qExjzzqUfQj45SyxuTEJ1PVxOUzANslulBYmoDFG9L1FKvaqGRC33GOE18wd
QmTMyr42db5AmXSMbjercM4/yykrjJxC+NnZOVpj1Br9/jX/pGchGdYY+kZlQCIg
cL6KyU+YnhyIDcbwk73E49HTQEEMPWe2DiFBTz+x000usPDL5ObRyzDK96Xkj2xK
fEoGlmvdkhG7SrO6oF5yBUJfgdKe2sYSrf90Y6wyZj1DI067sE38NkC0ErVGpp7s
XxOPPZxD9mPWT3ebKK3UjqMVDfKDqTwK6bE4AWs27kdK6Q4NGFPolOHog4wN4dEE
iX+8qIX41W65CQ3oB7tz2QIYfMWzQUK8C+D8AuNrBo+rRioXdq89t8oXr20Clu27
/n1Z3tOjo3M9S4WD3XpNDHA/mTJmaXWVZYiN3T41iz0KZ2vvcL/JEKQ9RV9aOmAp
+HT2bwCmm8UFg4J5mf4ET9dcUMpDccZga5vwES1HYLSNYRlVMUxpv7rWHpeKuvfI
kdxOYyBiOMPnOc5QknZZ6KPPwkMRUf6sVbDgqvX+BYiZm1brrSVDA13yydiC37xe
cNBY8sqfA+WaVuADN8Zd9U9DxKjb+Geip4Grlk4e1LdZbADHtnSALApoNhaNIPYt
tCtRrW+bvsVeSnUzd51QxyWhWRSCLwUBXO/x4OQtFbmI0HAbHKBLqm1mKbXD7Fdk
8vZDb4F3m/21SAXX99dMZFxzQp46vRqrk3MXMpgN+mhWvOujX+sCQ2j4SzzaEnia
F41vHLcWPGHrF5K/JPZddzhX6XPRCIbIhLeEJuQiNGF8itSEoStlyAt61AKZboeM
8JQRv/GbGCeLl4lYEEzF0OTabO1DPe+njpr2MIBzQ784NZYSzhjCIGWspqh0Cdfz
d07IpK95fm1roAKV2Y/svRLd3faSK2piM5EbNFOcrVcm1Y3y7Mo37+Gbn1vPiBnT
3oqyJqQ8X40H5RUgqihnvhZfzb4zEXY6iX2Rgj24ZYu27GD5IEyXaO3t6JnwUNL3
AuJ7dWUDAzCHTWePVuu2UrcCUzi/q9jImBQT+hZ8JLhBQBB18D9dnBOzt/FKD5tE
4qeaefEyLiWoOTmdblpnMPUxIls56X7eWJ1iaEtbG3END9pLHM2y7iMQkweD6/Px
earxjna37xLQkjGf/VuT6BWq+EsJWQFaDpB2HG3mMRgmsaWKtiNbr1QDJG0zej0n
c9gF5GByLRnVy4626VrpueHIaj8OAia9JZwONTVIMn7Mn5kY4sPmp1ErvC0WuDSK
LBmuxLH3DpNvmMwmCJTLvpzz3Jx253RTlb7ds0fmFcpO4e8SLd3d/BDRt11lCI34
zwhTYemriZP9kEevMfHQJvaq5L/BOQQ1tDl5sbbphAM1DulJSI/jrNWXRk+kzCB2
TQnZ0Stm8Uoj9eSDFQ8udUfL6HksUUiQ2wN14IhTILOeByRta2qF2IAAfF4IfPzO
m8I7CpV83VcXeNdv0MspMNC6Yj24lqEtgvuk5B2CQa5gvHq720srjaEyBTouzjx9
Ka/k1km5IdkRCaf9bvymxETmLii0m/ATtoVZGnYswnfWjmw2X5FX69sM+USOpl/i
P4qBtie6b0nooDIDW4vKlfhAhdtgMKvjowftl0a4hbNZlGa/mkDpFkd0It/lkIBV
Vbb0HKnbVAOf9lIt25wy+krsUa+Mo1Cv1wKn9qeRLJrm5ghCWg7WliBw4tgOQF4F
541DlcaszuinjGqH8+dORHxdj/c6ZymdjEguGvWSOmMUVXdbyZVNESCiGHyYRtCE
MLiqoSjMBY1/jQTABD38YvrKLFDgAhRDVt5cbsZxeR6BHxdhuB4M4aWxNTyxOSEp
Smz2S8lsrzeZTcwoSBh9GLqhtM9jJuO6T/g61M3HUiXShbV3+OlUDidS60a0oGZE
uRrocDA32SkFK7wIEJHwUPT51LyK2RFecoKGnnwsZmbjDs64B9RQKuI+AHcOmElI
8KF2g/nLFXlHcKrDLvfjSpSTIXOw18QWfME4BOZHVB53HshWiEmmZTBqO7Gumnk4
JtpjEybNS7ncM/u7O18WhbErZ4ULK0Ba786ta8K2V3oKYz8j6pZRQeUISeGmAPFQ
vzOrDqwKPqH2L4wGsc1zlyaSz0C9Fs9ZMa1Ih8JiDeNPDeIUnJ5Xg9jGZ1Ikjl+/
hPk8Udo+N6XiRG5GvPwvmENyN3VjRZNx9EGhy+WXOTr5bLt2vsyEnJpQ7x3r5Zjr
s9ktRbaV6I2HYIpXuQQiCYVeHgHmC+Z/eVZWFcrqLdMrANWJe4o/oF8crogyrYTx
XAa7eYAdtNv+vXE9CTf1t74vUrU9JQw/OHTChtUE72ZpCeijIYiKYt4B/Q0VOWom
zoDA8YPSn6MHtqJ9WgjOsXWANFMyayH9NsNW2xG7gyTvxgjrDPBkaLhMGZhsfGNS
EEdQqe/7gPpSUSd0q09UhUbrBIyEAwqUAg87B7O689ZwSKFGfAOBwcRJIzYAT9rD
RWdWlj9/HOmhTSDgKS9VzU19VqPmJIebDgZDXgE0gZLRcqgVPF3pjSQ6/hPvIvyC
1wTkJzFn669KNn1YAHJuT5VQFbmgAQY7CqUIMj77z2dyAq8UfORlqNcAS8XRxkDT
8I51kD4BAxaIiKup3BEqlYmdHO8bWkomsKukinNnyuWSufuO19KyOuNQvoxUBYgD
tBOpuFExmoSOO6wLrYbbbF6h3N5ZRP9orezhwRnjCtuwjWYDV0P4tPk1p5l4O1Ov
EKXdkmBQrL9R0X8hZ9MB+WEexL/rojrj1Ctbpv2OYkuf4NfORwlDmG83VuL6RjWO
MzIgEcugw/7lR5L/a5br2/qQjmQgXcIuOQkLuA73BKnE0qa/xvpFRHUol4PdCMoU
6qgE1brP3WRXtLYRGnmo6Qzwles9Jasc7OmWulOW81NAqR8CiJRlDsbuxLnny2pf
viI3+YwoG+wmQhXKUOT7AjvPvfhNEN8odCdIgq+XVDl8V1C9m4nwxY8GVnULL7uW
9FD8RFP39PLQHYQqy/Tkjqhoc8Z3QdsFomAgfOM3kJcvF73CRCQy8zk7QFWxU2Yf
d3Wtw7QWySGfRuwIwRimnsmeIdcNQPEWul/b09l7glcYtOF+ph50EaycWV+J34rn
M9d5T+Algl+L8y7tOZSVSr/MTKQi1PKedehA2g0SsFUjHVN0cPVmD5EyOyz+aAJ1
jUGXvQ0IhD+1j14HjHbhPwStX12hq/wMsZVn+jkTJRQNd1SH0K/j0CIkDMdv4tqS
DzLlG6MzeRQHUmjuCUxpZ9H6dGcFJksfsM7zt2RSReu4LRTTk8rnBkQGe+DLqhkY
ibJeAG1HvLuc172PEBXE8MfAUIhZ+fZFBd5ZuoXA05dGHI+jJn3ofBN5uP0RBs2I
DIegTz6L4BT/cx/A9fLTa/w5QOs+Wa95isCwr/rtZuZcbWxWaW3Sucb6CfFc0483
CLTdcgDj0drtnJZrwtUj9qDp2G1XM2R/FMV/e7Pz/p9wG2OhyV0yW74YKI3KLgzE
0IIuaARgBjvvcsyjQa5v2IaI5Y34/bnHuEKNNrDCPJr3RMsJeixRl1KBL+uflXAv
Kpv5wTI6sZtn88snaf2zl8IpEYhRBp0T7TR125YkaJjJ4pMMCVJ5PfBEEFTK65Sg
uvCt2cGiW//rWXAvv1+zvjoNSuW0BHjlYf02OMAk9jsDHo1MBzzO53ipp0Rvf8zM
hmO4Z9I6dKadTnuL43NjJKm026bV3eJlkZ+IODg6M1PDIETtIbBBpt6pJCLQIhLg
wAoHtFvFDB4H3vBZjcwyt1QDtsGgPWvTLbxGiT5RpzJuwSpO7UZn7nEQ2boGuVrn
H4xg/SZXgpw5pBdvnqLIGoNxljNE1ycFBqHoua/PbN8FkCbeo5KHUja8OPKRRk6G
DKJ3UNfzwx2obKjTr49UeL2gCkj3ABNgIqD6n7Imv+um2nR/rrsCvanMt9czN8pN
486nfibk0UX0iSjb0gFDbcLlBQmIRl/RATNsa8K5yAobsCeNyd+59KdLTB/PhKZT
BpdOxiEKijhza18cR0ZxQLb07untWMszCDtmLEEm7jqOUv3Bbt9V7dFxO+jk29IL
mhGKCzI6/kbPEEHJy6/a/X+mAvQEFw3p2a5p1WCsMcsejbkPbCMCoyqDnQ7bp05R
yLnxT/3ihcJl9Z8F+3U1vL7t0PeX9g4toTr7y3NaIh9gM6CKtHZRABDW3ScrC6Ld
TiFjMyikoOCIu+rMvAdTwbfcjtk4s0G7HX3uqsRsZlYA1XabZkywaPESlfcIFUZ6
Mdq71eMvOxjCKiaJRJg8NG0pgcMHEfGbzIDZtN6wIixOjtWVejXZz83dmllZwJ9P
Q/PIvcMbKH+vErsxHC5ghRR8xVy2lv1VTz+8lfVN2AG1XQmsJ0V1zyfHnpmg/ii4
2SHswJa4RugCv7u5nhRHYssx8BWHGtSjusX11UguEaegJmL1ZTIBapHbxv1iCDWP
z2+voDFJh60bb78k1RjHgPJO9XEJv1Er70o3PmpEh+SnmdQkRrYg5tb28Ol1vW6W
FDohzRoOntAn8rRsAn7dKrNCkevYLXZT5hR2HM3n3REnPQZ6aKautjcZKOL1ShXk
krUm0ggZ3kkI/DGaW3y0ZToKnVGBEBJRHT6C2D8IVq1As2BmhDcR3OOzFCZiP0ba
Per9Rb5b20ELqjELPh0A2Y8TM3Qu5Nc63vRz5NncM7YHHvPlUyqkp7fvniD9b0ir
TXNSRqDD+dEygV+yWuEtl6UhXDqHo8eNj9u/DbNHdmoP2ILPEPQYCDgYQ3lDtCM1
4uQ6gX+an/vCvZU7Xzi13Rnluh/UN86ZxIMBGH06R60hZwohOW37BVmj4O+d5Nte
yWRJT0jOY6LigXHOtaSgY8zK5TZsiu4WIMgQB5FcQF6Y6yyp4RbYC3dJYfkzMMp5
yepp2fWF/lxrxmxIs35XC3ZeubKXskLaQi/sj3g9Qlomqia8DievS4nKJLpHxWJD
XOzciwtKaLG37bvAH/6lUN069net+Nn6+qOEOYs97on7R0leV0gI6WjWPcjSM3SR
HVDBwXXHwADHhI+5ZQ31+XgK8FVCw8JlOAltY2lsx881rNxH6AcaIifAYYhAIICl
D5XjkwkzdMOZrKXOByn6xbpKKCx5gUitTfret+Wp3DRvFtG060f3LqiCYWM2DfhN
S8RKErrB5jrzYEIe+u51nmTlDf0nJGRz99YGELaI74Rs/HqqcpHUz+5WfREHQOP9
LNOATHICOUbpuaSC46ufBMqOvqXBDD0L+/sUbyMeeHbItXppMJ+SvuHvKYodA8m9
mvKnYGr5iFzZoN0fSLREb1zMxl8HJB3LqdGP0/KNNKMQGZKAEOzSf0p4/PEHmAo0
qz7pYblAMOZjtUairkSW+0LTCjVRCnWTwAYKkia8oBz0doKXqHSMUfpwbSQrYEKK
5F0TWCv6YKaL+9G/1R4V3l2Q1SNS4+c9pRny3mNksybm15h56KA73par3gMs+HZJ
y/FsvuyUDRWzQG0ANPe0QVy/2K/t4GU0p+nRPmlPyeUN2xY2CjliLdqBvHh2X2vF
ptJsL2NdCHxgEmeWstTIznoK9eoXU7l8wS2W4PaQPWyfYWhXpRbO6Z9R4AC3VF4A
dC7pB+0uWyrYnY24AWANnH36Ig2LR/sxwYZYioaQs/q8HlTSP/qEPN5kkJ9rGG2a
QQu05MTzMHReVd0prSxopuRaoJILgqIkn603gAIvxzlDZc4g4fafcRt+8qaft3S1
fvkKxCuO4Buxm0cYhizJTwkI2/KrJZqf+dGbdvjCOy1x1TL7fcthxyIqV2Gr/OiV
B1puaiPwbqTF/04f3c2fPEKKXL3KAClapcooy10436FuVBLofmMtt/cGiPpUpdJ9
Y9vtqNKWQ/COXh+WQIWy3A3ME3E7fhs6woWYQyLh6s61nuDEi/v5bHVPJzUNn/oQ
wkZBG6ajuyeX67r/SY6Pfg3HDAetrDW4gFiGUHgFwAhmLxQ3BLv3EWd+ntF49Hrn
IxXrS2eGN7RHaPKWunZI1f6aF+3+S7/MHBCqHAITqiyXgxjFckYgM+bIkDl3D0IE
cmrkb06nNbX+ALbMtrULAFl53/Z59veIWsN3mqlfnTblIRULABv9+90KOfJJCnay
taeFaFsndWGbmz4f7Ly6/xOSMYs5GAytauwhJVoZ7eKziMwNkUH1lvmPf0HdwbM1
btxL75R5CYFwyrcCKraUuA6qyDajPvx+lXLcEY30oGQ0WZ02jNUJfBa4wLbkH5zD
gsYh1CKIcRAmmwjpcSMc9/hCjsMSl+onReyHIg+5py7caeJcQpoethaKcsdHF5Me
FoMCsonurYGX+pR0EH3ucnQLqs9ae3/95hT0Qj5C6TDm50Xrv0C/iQZWikruwHtX
btoTAnfbYqKCtL/K0Eb00VTwXyqxoVoiSDgSQa6z2mPTrpSx81FFBXx70hZLcC4p
kZBxTV2RPx3zpHexMEkD6C8ashECHxgOM3dYD/5EnIFDk6nW4D3KviXDUkujXK/g
FYtO7SXZyt1R3jiJ9+JkW/lxWz5Qhb7VMYVBJs1wxz1yQ0Py0rPqHee2S3THA+0Q
5r0r3Nzfg8k2aWFpYSqv+CCnf+UBlIB1alVsBkBLbbwaEZepWreed2kfj/wCReXD
3Y7xXwlgtKW/bMxC99V8d41n1SXtXboYMVTaz3bYMrPELg4hYVHUMUp51QLhuoxc
FKKoFy2L0d2ZuFutY4Q5Xws8Wa0K2WwzC8NFW2CYtvPPjqWQP8eoi7U7BVk8p+FS
nKj6x11S0ncVxVU5n8xklSzIQyyUMIW15ZKNz9vMzM5dsQ+X9JQ1uOKpleFfPGbE
Hm6nqnaXS7jAmBOc/gx213aEebwF13DotWLL5EpdjV+hwckjklfv3PpekOrbGYE+
4RURlazGcmLt/B5Bvu+GwknP6hWTXPmChw+XWPYnk9WOSUwCYPWiCL8Nojo8eiiy
DH2HFTPIBR2KOhUqXUlA/qgBZhU9DslnsCpqt7LnmkvOwUy+YQheX2DKoJw6L+0W
hEbs9AX8PIqspsDqKGC5sOYgQXbRG3KdEpzQHCVjyIskwabpKqVc36/J4SwjiXk7
OLdCR6lmCLs+pBXCcwXFfiUmz572jY8t4AhQOHBAAv2nE+u8tVZ0pzwPgzTzcaIa
92OBnRUSe1dd8ToAkiasUNf0QYtMyJAI1E7Bfrr5+4yWqWk4Q652GLWr3wfnMZjV
0a5KcoBE0WT9ZqMEUAh0Tagwh5MxDcv2krUX7a76OM8tDJP2uGateWtUvF0wuY8d
JG8Di1jWhjyCXZGndbXfzzYXZl9UwtVw2pl/Zj/a7X8+apzNFzq2mZ+V/hulJ4Ix
kucsq+S3ZAbkeO3V/msahNxldiOoO0015/5bPuGueeCORiG8EmqVGKJbAJuZ20Tr
weBBUEodhHcwe2UriGGki4KtRXJGc+3zW6h3w+AESy9gKUSu+QUxBItw8xJjl6NO
XbfU5eKyOrTYqImwaNUWka/5Fx4ZpkSVqlSQ6MlO3H5K21q9C1PXTDR+py00iAqn
IDwEgvEwgZJwQ0Xdre20Sg/8jDl5ZuavboyIJlFbi7TuJbCIIsIk6KIZvlvGQZ+m
T+JPTbDaojOg6GwUyUDMB1yDiI8jDThRTY7TwrtU6GY7zxPWoWGIO5gqUkDb/daJ
Lrt1qSzZJLNABoRMU4WR6JoLkApxEjW0OCF5qDX+ms+fsxetKCzE4Z1uvHIKyZ+V
fJCJxuEbdMlwoqPOEHiq4vjuVds+kmn5Rfjj0pBki/3b36VR8rqjSct2aclBv5Q5
zbNmMe0h8cERCdImiTK/GORgpepKICgo7ILgQSYpqd64hjd3r2D4qdWDGmHN7YbO
cUVmYF5QyqWOAxVPrL+jgp2ggx+bvFmXiYDf1TttQy1epPfizYMkB5JxmhnyiKIe
Gd7fMg++UUpHyxHMzrPj+kbXprPuHWupvWIwFG5bk6p+j9NsvkDX4da+sF0ATL8s
iumw7QJ2kHTDTpnfBx1vm8UFAKZBFL/JvuRplK8OXcKYZ69vP/0jjOdqFKVNjW1T
07IB4HAr7mTxozpXJvK3XScn5/vs0Gr8x/plMuwQKQwjcsN1WDECr8ex8BbuLCqh
HdeW1zd6Q4V5BTEeQVVStzuGczL638YlGdwRyI1tXVEl32SZk0pZ0PODKCtGuXzG
MWX6AlaCZP2JCM7ixgiFP6QmbrgS0CeaXmz/g0OkQyKlK2GVG+jeI/u1My0I++eF
0tcxuDFG7mVXYGhoBTmuONw++aWQsl6+E3aIgkFf3tVPhGHJSI+mNLgEn9610gna
uwQFwwt5uCTRjdeO7xSm8y5x6ifumUs/1N+56XEtP4tEm8OBwtEcsZ5MBMxWUrfG
ud5blmqfALaBj3LpsmQ84VTGTwn5QFGS0Iqe/qcw0Dj0ADzycFIoqVs6Jwvvir3p
ryPJ+1jwVyQx222obc6wpGLmZD3bd77Go68SHjCfVmgYToco/Gv6YQMTmQOo3wRi
gdfDGJZoqsjSjPPN1L5KROpYzCDv8Y1yUn+TRz+N1vEcabUS8fMjyTOvrHk0tavO
gix1hhwozuLGDhTTQ+w/CmvrPxYWlmfaSJ9W/sPmuaY4V6rdMR+3jmbWEjDSfXOm
gb57fkQ7CpYF0mkFN0m4TyrWO0/PVE5NUG/mFtWkbbyC8Wxhqo/1+UQ9Xqdyy68L
rmxFiHUfyLG7jP9rTtzn17/iIuaSPIVP7kStHQjQ1puAFIlPZKFUNxEazNCABGVG
SlLzSAOaGvpTv+PkQH7wOSYlB7PtFKY6vDqJMo8oOxGNkJ0ENpL8E15NZ6FkKbPH
ypdXlc7b7dHMoB+ePi3FBO5aqCXklkiZ7BwrI6ZU73PvX+APvnX/FriRQKnP8eQo
QBZgWI9Nsfzst+4EeG9ZwmJuzWOR1XZokCwoik2cg2UyeMIAmC0b9hiFUgU8psgD
9TKOaMJ3GK7cCj92l2S9oF5/kjFmIsm6pPeS1nAhOJ+FxFgbKTTIh8nPYAsly6Ez
bl4XoEyKCYW0MWW+Sng8AZhmx/SM8yg1t+WW24xSx8/8tS8EqPrctMu5wcQ7IK+r
tokp5+LlhwQGFs89V9MtkTBVtCF49A7A7K3RMwFejrCMhpH8ubIAJ7e9b2fJVww+
GEOT2DIHX9PWq98XYjhBUCHTI7Q3bdxChIwKeKv02vDrxFh4O44Ijnmcbsc9HEZY
i1kao/aA5lbQxkKP7dqHnA4VPhxlwxMir1P1HS89DqF/mm1NFa1ENf8HEgcTx3d+
rmvtNcoOFjlRvtBnZRF1ESeY3W1y3KTDhNxkWPibmdpm1s9IgzG92ahG4sS8FQbp
/laEJLIx1cKSGRiHRu5IRtOA8RbkE0xUDm84Ei92axt8DP0uQciFMCwm+Dhvdldq
Ibd0mCcN4goUqpKN374whEOIC9iMLhhBG8r747mcXI+3xC0QZe0abtALW0sbfP6k
iewwvvY7AqzPCWoUhY6vzjjI6k04QqpIN0g4Y1AUskomzHKThkb1WAG9Ss1srRBX
Cn0uxRFzsf0sud0L7ui8cckCPJZmtxw+SzvfhiDrMjc6bGyvKrrtD8umrIXHRUM+
2gsk5UVc4ke3Ts4yRZ2s+zneVqPToiOoMz9bJe7Ojyi9yYkENAQPvz1XLrSoMnQr
oFc3azyd89vvZChDkOeWMB4bduotOCs9svw2VfYgle39DqqP4zAZewowg6bTk3xA
LQtXDqsRMiuE9X5oNZ9y1zjVHbGLF27qPnirq+CIuxuR5hm74pEs8rdHGqo6EtmZ
UQiUHHizO8/FJhhmIOdiXB1izaBodoNVEr5oKdFET0GCU04wvUwvdVx72nTY6ofo
ryI71metOiQkEarNrQG1wNsBeabkdveYP04RNpAzVJa2adyg8LnDZRULQBEZXdP3
8/AbE6hQdWsWZXyKsemZw5X2Vi5M0cUA1KWxTqrtX2X/klEdeGqs/Sivb+lt+86w
gHrh9EeJ92HOTaP5ZYEDaRr/Ewj3eaq/BXrhLb/8UuZgI0VaH1Ye1eY7ZBtQrW0H
x1IeLlpqvD5VgH9NfeMaYfnO3R1y+NbrVa7HYzA8sqZftQjPd49RgG5VOkUWyasA
SHCjb0xMe7ZOLxrQhsnkRitZqWVApocOCTlbj/pIPNvpuejJSiCpDOc3wYR6HA7u
hehUXJXcCSUjw6S9Wrx9qoqlrpSGtAN+sbLXbuZvxUmhTVODFFJZIM+5SWxms3YK
zoNVcFMzXeJZQyI/3LB3nBDtfQm6EGg5P/jl7AFjjk7k6HSzwFYooa3bA1xaz6gk
AG5QPxShq02B5MH5upG+0VFeO1fAcTRj+K1a1IIHawL3j+Ce/O636aroL1L3ZLe1
LyN2D+hzWCj9lH7PNGmGt0n5NJ6g4ptNPdtoE5FKHdJqXM/9lVr7RToSRVBNPe6x
vK5oh/3k6TwzuATSzIFD7ijUsBhfOWc2hVoJMUS5Hi/UtINROSYsUnvMfLziNIeM
fayfdbCUQyS/hPH4kdpC6CrycTSHxRpzshxJHUs1AalKho639b3r7zy3+N1U4+Uh
bkpBry8xHOAX1F8nMxk3IkO3hEjXMgNO2o9dsy2Fv1kAAOImfVBn6CPU6inZltUa
SBkJAuyTKA4eUS5Xl8U5Cd4Jnkp6Xcxp2OqP5Yw+WsT00Y7XsTMmoyIGWzShvxvd
qiFNPSemOKcoGROsejNh3yKS/7jZ0tyP+qzEj4uvqaiSl6e4uquyWOkmY3vV5SyG
3A/+Va1OvJ6hBqWFdIF/URiqUc73/NZMga/H5lW91xBBkH70n9MXpN1obw8bDsOZ
08TrQ2mbnIJLxq54dyS1q536W7+LJlH5xvmYm3UVBx1QqYkRAFHSuAWRHFwYPhjl
+2UviApnRni+AKZYPk7J4YpToOJPI/UgE9lGM0dfWuJNVwPsuiFQ0+WNs0cCgpwr
TL8ROKlXHEWFCMmmolJHvEW+x32hFkcgbYX0k3gdS3qz5h7En2Q/SXy533typcBI
7dyAhN05r5w4xUBiDxn7TS29LBly96N8Sd7iVTUEKtlyDPJedN6WcLyDs9BJdxnu
skZFSSAsMp00pE6qpxWSIlQ7khBkOwxiMkIegjO+TCdBRS1/bjGBt3bk3zIQ43/P
eiCCgngPMJZJea2AuNXTKjcDcE6+Jtpz17MJx7pO9rjrEZd3tS+JwGqqq4WK8to6
rhzlJQDaA1NahRkLqAkS5ZQK1YBNbmujSZtm/c6Rnplrd57L5zTJnZyuTWoC0m2x
lKALR4oZCxOhyPGhvfSVv2/Tm+oUXP/DXOjDpgGGTAG2CjQ+aoudN5AgG06or/e3
IGLliCwNvfX+YNiY8ac3ZjhsCdu/eHi8b/Eqm4luRyHP+Kgl7smSa1LlDiRNokER
22FLgrPmPSI2hE76f+zxtEDJRf6ozor0mjrS4ONaTnB63PNOVLw1Dm5sbpiFmW9H
d4MHIokbyiM9aDIu8tC2Vi+CEWZG8uUHkcXH9sS85F4OieS/4F2MrZuBaMIeslcb
/06Xg/Omtamc+RECtBXA/9D7wBMGpZHO13wmDxp1wUWi5QH0fHudCx0pHBDS/NyQ
4vbICP8KcWuicG9AYkIIpCdW21QIsJ2zwoq9XeiWjsA39EPhCq1uxUbAh8ofdEJP
NQC2+gXqoIy+u0CwkbM/RwwycavkbAcTMZf/2Io/IdWcSo9lqOemTwyCil/+K1b9
7HYuB5JrP5la2Hj+SM30PPDSmrAP39IF6woccpCoMXqN9hrOF5BBcLJOI8aN969P
KYkoIAjUlY9Ypxh0TCMgui4qChzYIFZ/aofErDq98Gx4muiJgvim/NVaP2dlbppL
2OsuacIFB+57kx+CaedqWc3pu7h6vgmGE25YzFXBVnda0QeAgIQQQmice73Qzhvm
XQ8TZjY0PqAcH2vAcES335fpbtkF8epQ/OE0kiHttzUiajdXcsmGitYAb7lHY+GZ
EUtN70/aY7kzgrWnzRRf81OLSYeS0tAsheYrvG0Lxl6Y6JevVPQdRqy4LYWvDkZk
jfl+8To1wURyZg7BSiWLQ/Q2CreuM3x8x8NCSN1gnV0PN0sYVFpacYabwfUsSvqM
UH1jS7pDbonWNt5IHxGHRCHbPWbMTCttZxlQSuH0uysD5Jk+8gCPKOOpZ1vdBeIA
YZBzrMp4VCo3mkywQ9oJF/Suqp0PxwDP+2dO8QXkgj8manfvwuyru2yN8R1+dDVF
9OR9GVvzFKic8h208Yj0orw30QJTfPhDqlI36azQHRsVSzjrviolk2rS2+q6bv4i
J0GjwKz8JwftoQAvLbElsLqZ3qM0QvnTHRq2clk5aHHJiUJiJrhHp2+K3AMXjIAv
7r3s0ceqsqimwkc/Ct9n52eT4IJmtdyQY6HMwdgE2G4FKuF94fc4LibwWpuQihxw
KlSdcmlsla6TiyUzQIYWofb1mrbovYgGIluH+5F8o5FpBj+AytEeeiLE+SarfXPM
v3V8i/nwG+iUm0M/rQAWhOOafdle4rJFggvd8ZRBq2YIQON/Uq9awD84uamdlLmZ
d/L/H7slS0fF/P2JyCRGIBQ6eUw1XccCsvwiP0xgEqJ50uNaP9k3ktbk1TVqJkkV
3Sj17wm1yFI9JStd9vTykliabDENuXST69hRbaRyOGfQrH30+utea3aEKI2jkItL
e79gKdSRS0mZkH09ZeDaN6zdWACLCr8xCOY7F6+TycVlTjJVibaJN+2U2NT4VBD9
fwr/IUKVuPZUvqy7phxo/3OtTEZp/iFbZSl+e7BaI/voJPhxrkKwij1anh+/T2iC
oh680OSshXilu3IBjAhJWYNJ8JlTT4KV0dNQlucBlMPKaOe1895Z35+wl0Jt8FnX
cAxUhTZ8ZFL5bI+aaXx8DrD7tGqQOY3rQeLfK4yFlJeg0ZaYVcoSV4FpmcHNXa7E
5C/Q/rj2J7h02ap0B00jHL4EoQHobUZaMtmj20rxeCdFj5pSf0/qW7Gdrd8nWJ2u
s0qJEoFYPRKZUd/DoFFJzpBJS3X5ItHMWef5JzXfhpuJ0788c2+FxBB0CRLjC9ia
bM4vLSOPdTOlrhJtFkv2IkA51mpp3fak+DiFnrAnSd5S8FuLXrUeEEL5j8d3tD37
rRjAlZaZz1a7QGbYqjQoakWGI/cpIDKQ6xWNyp2Xh6iDwf/NzH6JALUlrsyVMl/p
THQVZ+wQRAJYw9yynYTU46og2lMXfMkl4CQztI2pQ8haCxDCoieEy75d8/yyocj2
Ct1Om+do1uBH5hzX38978Q6QklgTfWch1q9WhoqgLZ5pr05VhEBV/Q3W0eD8RrhK
UgHbMQ1lEBYMOrqkReelzxyWzgb25g2kYhoNWDg4zix+B83WthOhDfML1FlABI14
UXwpKxxtO10TrhRDEhbynCGrsgOAtF9TJpw37v6lY6NgOIb1B7sXZZ8dp3mlsR+I
/atkhVKZ6Qkfm2shCghDzABXmHBpT0DzCzkC2Slt2lTTO2F82lQVf6TQZvjkPP5x
0WBNU/qjf6F5KaUyQi3Wsvq9FBCewejsjUwzHXPyhWawCii5WQgfHTTiuWIjLYnP
aPLQ67vmc+8gbqZdfUj14lyQIkhW15c2rPTis2FOzJ1/Q6zGFhQF2glnHnO9ivu3
5U3BXxbWeSAOcGX9Qhdwb29JhZCsWsWUPhhnJPWBXsHEvvLuF9pM8LpGb9Pv/QB+
9NPpGwk7DZTWqTWU6P0CWwr4FBapUOH84+kPZ7QY789E08b15QKGr6Nyz058JmMo
5KH7shxmT9S/Ms6fg0ZQB60+eQMGL5caxGhhH2EZdJWTHuy7zlsce2go+OQ/I4Oz
ON4qBzBafE5GjoFIUhnxT6vqOtkqR7AkOnanlUlndXc7XGtdVK45SvSY9hG5/OtX
Ekx3IVwkceAsRnQCE65m2yzs5rOdYyOwm+UN11rX7cMmC/Yk0KyFvqAuhiI5l7W3
9QZ3QZsVvZloDhUWI/3k6Me+a9DtDmCPGKNkLLtSoYDwJPh5Pp2aT1fB1LAHqr14
fTNXk1EaRwsBnewd5H3A5vvHty0iHBWU7A9QUdy4o6rmMl3EvRUXt3T9CyFMelPv
p5G9bsnkVDWeOWStfKxhWnezQyfj/d90qpE6MDHoQI+SAdjYNqSMVZfTqbCwsYCV
XWXJtrHsWAYdHvFBUKojX8vHGAsmoqD52PqxevKwR28p+id9OoAbLbQbuqVhVVcR
Fik9bY2c147YUSSOlzO3Vj/4N7I2ydw68O1stEjQTpo/9VLJfPAMeSOoyZU0+/8U
G9Vs1Mm1f5z4xmhHRIgR44yolpbmoV5BYjRdC+83lwmjnZ46j7vJlw8x8EITGPXG
RoBDJ9brkHmFapoxObszkGGjHDl6f/sw4rChgfJA1Fa6LZDowcxfHT42p/aq6nwU
fLala2h5b+ziSglUHltbe/E6R6j2zwredwQhJfrAevJmC1dW/8PIUJugRPNbPKVm
hPxm77D84/VTsGiuXnwu0ibjaWo1bmZkw5Fa1zzeZYaTLQPd+tTi3fIA7Bp/c9di
tAPx4B0w/zeuC+Le+VMwVWhi58IxcWJm7eCs8p6f2/yru+bS1L5quRfIGrSiLqiA
Q9MYR3014d9hQZgm2OQMSs0zx/+MpchhGLO9nkYcD2/Dj/XfAlOuTUx8kYWLFRec
rYc3yv2nKnzmrrtrkWJdiskE/T9PVKOZDsAp9mELtRRJG5Nb0h7DfYYJVBB7j0Vm
9Lwp8E9RwMcmqw0V8t4z51k4G1UeJecEZYbEub3hoAFQ8wQpzoHFqwnlFVLaf79q
4f4Na53O514FJEtXUyvX9vDgQow3OaAftnyTWKmH2oOPPZAcB8R1NWzobL6HuuUT
s4PbVU9oI4oNuINa24Ly+Vtu/IT+jVXS0nVSNfPvab4LMWSPxR+hsOTX7+4S2I9w
jhhu4mspkOQbUodIJC4FhL/CCMvG6ZtyzlsqGWjnWyJP5QnFXFu3LaLwgUjg2G0U
3n+thXg85XjP4Ut9XQ2QSzV4jZZIVWUqTS26AoK+XfJ2o3HcF1Brj9loVzAYL8ot
tHM1jEirvVNEqzK0eZa5brSPmkign+OVAFh4M6ox+so=
`protect END_PROTECTED
