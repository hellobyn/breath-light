`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6sBRBbyjt/pySxinUv0K7hJt6nem/nz9i7RkNSZVV19yESWntOwv7iFcj2ude4XE
il4l4SQaj4FCZxV9qXbZGPNs/fddxQi+rWYl9dmm1jXDLnCuA+7fr9+t9fUeZICg
35xt7WuMv+BXW33meTaT11bXJEUSa24XRH4Un4bS6/ZVgGz3GMTP/02LQMAMbDlU
srYU+06BYmSv0XUVGyCvsokw7vK/Xh4R6RK3JFcVOXegSQBp/3QIOWJ+0hldrqUY
oAup5iTP2zA9OgZeARd7zBn7qUzhiIRTm0HiJ7qgT02R6h96LRtlqC93zKRCiXxP
2JX6exWz+8VnGdK52yK1MUYlcU+lzDYdX2f9juJB1KPWHDDyZRN7MZ68+PUV0f/q
bZ4fDwLDfYlxWmwGzRUarpNph2H0T/HGUu23fM/eoJh4Vip8cymQa6T2Hiv/ImyY
Q0TF3AqGGtabG8dDHTE6jOnY71prQZIaNU2gSNP5Q90=
`protect END_PROTECTED
