`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKbjIm4Oq84StW0gbsuGIahGH3nMRXHiW/XvvUznAIxlfFtf7amFoYIeklur9lsj
C+yxuT8A4aNgqa1dSHOwWAfnlbn11BE+RkW4IfcrZ3bwouWPDJTmrPhzVuFcT8Mc
M7koIOe47TXDttqvN8DtGnRHwzwFi+WP35ZOX7BN4otkF9DoZErxP6Js9d7UyGXT
YP3zZDKtmDZQ8y5U+Xisu+FqGCAd4DZ9PV3hXU072eRrjN32VRSkmWUdkwDZz27c
cYDyK4StPK48V2UURfMEr1mXB9NL6QPRzfH4saWWRhb2kfAY7zOQ71pNWyaa3qK1
Uote1EESyKZgS4WYgmF/IdIxCBVz6r0b1eMGAyK6/YezRVS2/DFIIf6iYA6peGuM
WG/Ulv+0uLbT6FzuEBxBNNLbnQqCcKZf24NABA6qfs7xenyEN/czzL4QaNCjWjXT
+en0gGAZNHN9xW2jUFN3mITAs2yax3CD4DxRuFOUjQ7Kde6nCzGEUTpIQh8KzGvZ
7sK+sh7HtiW6QZP87WdcLez50Z+G6By/fSUkt63ZfvAVWPj0/Nea32mUJkOLiTFr
sGkd2BEezqffiBVYUIxi6FGa4j8kJ/rTwFVdjYBAzRRLpTuycW68ZSJzwg45OzlZ
TTBpZjv+RlyKKo36YeNBhWqdar2dayAVoviGPJBx5fDrKuE2pL4iKWN5n105jdXP
TDvCL7RiAIvgiV59Uj1KmEZI8V3Q8v+lTTuJpjY/Gbkf7V1NWvKwVeaUWw67g6ZP
puaNmkqfYa315hyjw2TCFcpi6Y3aTBlpW66mEyP/235m3gFoWvMh5Y9nQNT6N4x7
F2RLrNburM6hncden3zhP2aOg2oPMSiicRGVcFMPxVVLHxrvMJhmanXzYCskcb6p
GQxMG4Uw3seIG4VBj7Btgp2EQu0i+0+w0b7XBg8ttB9xRFP4fomLIR19DbiRe6lk
Kfa2CLuOcpJDKBX5IlRGpO9oDV0lmbOEk9C1u9+lZTLdkOYuM/++I48P5mkHnABR
2H7wCkyXcEXu+wpsfceGcUBym0XxWPTWVhRg35/T2wtoDxAsrHijbYiZU0w4pubE
cRINizGQN7S5OYanEZjH2Xy9DZn0To/Rf3fbRb+pPTtYbtw++zuEyCXqE5MfxILi
lUzsQfI90eEgTlQUZo4HdhgbgVqS9YvPE1tv3P+EkiQD78g28f2Cj1pSIsYy7h/a
5xPHQXfNod5DA6ebZUOc8KnamF90MYh0J7E5P74h4dzEMDM5almQxNr7RTQfo4pA
zTQDrRZy2y7woegIa74D1UBwd+5b9+mlWHr7gZrMSZ3WIrfqp2Kz7USqE6KYj5GC
/tnohvTXUWazkXLRBGZN5RXXnEuMyTPSdBrbbJAIncUzI5wcyVgS4H5A7L5zdwyF
MJFtlZcMdZ1+2BnzO75a+cUDZZf4yqOp4VGiTZ9sF9pvAFSlHABmGcLhTUNek+uT
H21uch+e13iWCecUtKjOt+zky9wxXRnpotxagXeSFXGZU98RQYTyZ5o3ouIYiCS0
wTFXKwS3liCDtTUThXJ5qhuk84kPTCrQwrK6KnaIp7s3c/hLXrq7BIl+OvHhgqUw
GLjk27V/wa/+A9iDkDcUFc00alAYJcXhjXMw2aVb8MlEQ8LF5ILj5d8LKubMH+BQ
fbVIQFemJmbg/Y3wA5tZqG753nX7/GNN0kRnjnzvLYt5TnchpHA3vqoCkPmDIYHg
XwrsH4s7pkBYbo6ciblcT0ZuAB2+feGqN4Psz4Kns9Tf72yGJ3ySh2gQPyBWrvWA
D5MdITgVdpdvY8pm4QqTjwsFTMyMBmxE3iTeiPTmvF+0VRtS9q8LKVJUyLGKK/0D
LPsba8IO5ltDhk178W2w0HIB1+V+xsTcwdYL4/OgH4PIc9GSCg5JWwfZa8TcDuNs
uI7pPhdp0TM+emI4HS0BXuPvbUC85tPWQ/+7UmeAC3nKOWqJ801lYWX8FuCcKAH2
1QgsH3OJ9KK5Hp6+wW4KzNzDiVIaQ6+IvODp1chg2ewUoErcEPKJP7LtI5DMuSQ9
kDDQbpipxsDffVCW+gOyvOTzA/9PhBP2r7RpkgT4dhU46LtxC6MBceYjS7kQL5ba
UZCUaJUKT4+mqcA096hH9S8CknnPcQbArIc4vKE+3/OyXGleCjVwsZ+GNIx/m4KS
YvBTEG1khfEIYwxSHO3335L49v27nzEoyxU55bTvM5Ii9+IDBNZyWmYRGxCjg3Fx
iPTIKtCA/bL80GFsvznpOm9hZ95Nf9R2MiJXg0JtibSzui/zCMrO0udN+z28lYiu
j1FKv2pGEx50C/qfqLhpViC6UPciKCzoE6Wff0WpjHJDMyCXQQwhK90iEkkjLixI
eU0isytttoOt0JgYMZ7Bew5SnHC4SyCP8PenXcq30Gbr8qWx5tOmUJlqlaIxohvR
o/Dtpin2dRNlf1al3uiSb9CjROsghtGiO1x/08jcKhgsCeupycGSlm8kwt0nIpZc
DetZWvsWi47TVOURtMTSB4pZ1Ejxa3ntyPDEySMe0SEGhVwVwICa2k3uQpXTGygk
0zMQoDvipNzZXOGXCBckbFcYlFJ1uK5gAozCSByDL2lU4wBw1DXZjOT7aAgcAhe1
IzT6EOz3frl8uH1pWifZP54UjG4iAV327fV8dMiUXgCqR8hno0fIcvDuGODAzxiu
Hzpd7FQHJYpmHAGKrUtDru40J2MFjAAok0fub1X9sr/rLBERb+XbRMWzQ78NEs3q
1jjSLiS26nsp4Ut1/3Xv02rx99UjSL6G9wlazhtgsDr0In73Nbi+lqfTI6DSyaFc
XTYADPMhbLyTFVsJ4ZcGzlDCbNfzAWPnS16tNfOvucSXAanXSQb1WBgV3BDpMzFa
SIQSjlI2zVlV8DST4ajZZMlMyeYBRuhpTtRujuJqZhtL1VCkawlz524kImiqVEt7
ozI2sFAvy68GnPIHbQJs+VVT6dWbwum8QXyQ4tgECDulv02VC7lcrGNG6TTcWZI8
zeBV8r/aUrdKXGopcN6jqaGX3krAohnjc39ooOGgz2goyjWdmGKEmXifplw0oO3w
NUylsYhOPlW9K+BdNoq2Hs7XFyPAxa30QGuSci1wYtsBA1hgBrNqx4msazXeXMhz
pNa/Emo5nZiGp4h+1FnP0/3qPC2akm7341SiCc80jBPOWdIPd1nj+4TRCYTWempg
gGOz61j2crkLwHI+xN4LGYRIYXy9OVM118hvxOwzA5PpHSDSjFCpGm+LgktN661V
PTMF0qU8kJ+DioAEsaq3jvxAMTdyx8PhFX5P0jUhRMqKube178QPOWND6m03bNNM
ZTstK6rRkOQB3xmIWSP5R6yjl3/UYV3Lo0X53f/wPuPeKTkhdeTXaERZoivUHdZ2
n2RCntGR9NN6tE1Ix4rln1MVUuRykKhl9JHXXEoLv/RrXGAA4o/eCWU+cm61hu4h
Bl2ywsik/jZLQfz1WPWsX4ah3Vrdztr0uvPL37l6oQQrkCv0CLIR7zh74f+3BByz
F0WtfMYhX60PdQ6N0mVikuXRLB3hCYNVMEbVa1/H6WRK2R5JIjuD8wPf892Hztn1
w73cvoauUkB7AUdKzYkWtit7uKxPBHCb5RaHqrFPLCea6vhPQHvxV3+9DZnoCzfE
qXg79YHMqBWj2rafzCBQdTArC2hYJszQpA+2qCi8+tkU3x4/mrx2TuRG3lb98HcY
sDQBQIZsPj4E90m/PvJa3YmAB1FlygcLFOJ92bSj8ZEqlI/Hu+f5gTUF1TXMg40l
K28jrSJ1LPbPhTExz2hgTTt3dqLbejPJaHH/nwiriE0Z7pD5lxvW676gJVkk67Mt
v//iB6h6o3RiCBcTc6YhSM9khY18deRDRiKX0Wqez3cWoEuiehs8VUfwIX5YPHsZ
g1hm5LHp60gcIz6kqTZKRfLyk+AqkVLh5PpSHPfeMl3YuCs73Dvs74uGN54wcTYY
bm4AKT1WQw7MLy1RqY1lFzhMExW9tzQCFY5gYVLS6DcnNC16bqQNuFC5X/sAV5oX
cMqF7xq4biopK0Zt7h4ZQThnZcEmXfOsIVq6uTGp5di6YIx5Ev96WM8uCxFvbd0+
yGjS+PIqRpjZ/Is2mbajYHXu4bouX0dNmcz15HTT2BEibzG8iXK70yQdnpb7RL11
ION6mii6xO46UkJFa6ilYU+NZbg1rxjJ3iwoBbvKQ+XMQuwTSl29uhRMwvXT6/V7
9ukTK2clKgJr+mjc2713I4gmk20VI/Dxee6G4aWksgac6w88p0zD1vjzVs24EniZ
lUQjwKEijQ5h2z3eZW/G0FCEYMTc2d7DV7EKH7fn/Kk1wnEbm4h2xft0A3GbxO4G
6Zc+m/K3A48yvLaqUL0FKQCcZM1+0r357WM0XBm1ws+4u48xABF7NAmfdgdYero+
cQnCdbuWJtn03aV4x9nJl/1G/9MVTdwbMDuPEl912LqFAgY9hSQWskOul9mjqXgL
JyMn+/p/QO+Hi6LE8MZH7QWpvZk3UBPG9slGzl8Wb/j/L+byrJn3Igb8rnpwxRxb
DTMYlMVBR2p+eHr2gE/Cnm13z3Mx0B4x03JiHNZlnJG2Yb0tK5TdRJX4U9pX9dEn
Lfwj6FnoNwqeVu2iSWdi4/74WuF04BEiDMtEpEN3zy/nyACijEW/Ry4G3qDzOPE7
+98mQM5Howm5cLtdcploX0XCLqlIszOuA7rfUB5iKSSDdAnBDD/PbXM1kD2br6d+
9mBnUv2YMUl4mtVhv1OaaxTDcxezW2kiKk8IrOCQvL4jgONWnyQhZTeaXZ9mN5m8
R5w3Th44T3TdPk04dXuZDeoFf4u1Y/Dkyy0GCEe0JVWFtqMa0Ye2jYu5n4Gi1h9g
XfA+ht+iSkl6Qmxi+b6oJnnUQ6Sl8fYqdXuowdCNLgt7FnFGlwcaPuyBYqpnGLSv
PxYevVlXxtgO/gBuDMBwIuxujKx17Nc/hyVgSypbBfB1KcfWF4Uosbe8a+6g+aFd
vPywDoyQhsQNMnThHsHCMy+D3cjBVT7lQm/1LUGndkI5/GL5rhXejFUCUu/ChqNB
GF0Llj7mx4q+7zFCPN0bk2JOAv1Psz/ZlVCf1sSVfUSvsqpFjh3uxBKlPP40LtJ5
3zGjyvLfuHxl7nZW57KTJbzfLFFJ9dZN1I8KmHQhz5eFa3Z/I9mM0mNx50kwULyl
NTNFoDj6m7JTkY/Alklkk28sDozwzmtAGiNfrdVK/e05L4+hMVlfzsQ88cBUrm7l
GAln/6jswucU06cWOk/sW8f+Dg8UERbRtLhYzR/4xSYKMK9w0uBqA7rEfVN+2DzZ
deVm3EwvczyiqhLKtS9wGLBpRbGrmATOjwQ3kXiEEWGRMTZQg718dzI880n6VAvr
qadC33NfRFmWJ+OYrK3CDWajdHlVLNh3gVqvLVG+u012Fr+j81lGe+HSP9Fm1QHu
pgyt3aOVqr/so+zdl/0YB+Y/u5C7VbRjx63knrcl6ebb3PAiwfkV9RvdnkFbI+Xz
StiGkTkwJfLP8hpR2v6IumYUaFmZA3vTp0M62xd6h4C5imTEItDad7D6EPCq1BO7
TDAoYpMmClbVOrxP9rNBc+ID9hXa/QEM9FnCP+mbP7su/V4yZR3nvNIAzaUwzFE8
9KKcHsVEjwgPl01uECGQ/KTH+3i7DHQS5FMl6vwPMiqZpzdKclVY57OsX3Y9a7Ie
pU/vTdahbzcpEX2atfHg2dxvmG059UZSgMfnEu/Uq2eIhmHsuJ/2bv2IWmqO88VZ
7kDNksWxXquaoW4QuGoRSOOaWsxFweXlWKIDsxyNg5y37DKHsChp4sys0V4o0YC4
EQSJLiIJSe0/RLzSqM6/aptNwDvt+q4sktz5zWZ3ENMoLbCOZJ7IIbNYOE+CXXW/
R+/kTZ7tQwBFP1hoxtXMb3jRM+m313JWWiTYjnXP1vAlEKB8ntzz1xpkSYcvvlKL
rlKTBKMgM3zhisYVt5DhdQ6gervMzVAnl/Op/ybg1HI7OYqduelVN9++T/VU7xl1
icUPEMlOy2LxCYri7DTFfyZ66xRnDZAJH5Sa49yNlB6LioPzozPpFnw+BlZdFOM0
FoKzNuKZLTpyyo5FLgclOwMbY/88TA799/f3RGqZ2zwlIFosM3jeEVRGMt7bqE/Y
z48ED2kuRyyTMU4ncTCraMq9jj5A0Obi5jc0YscydCEp5vrGATeBixvIPUIby4Rq
AVkJ2u37GocDRYxgbU/KJFWDeUooWFjSeerlxArH7bscMnpSnMKNrjnqtmZn5jAC
SL7fKxzJ80+hyarSQctUwkvfZf6cDVtN9/tfHiUn7DJA2V5e7mburH8Kw0t2+aLs
mx9da4rVJHOFLsfDmX7rmcO2dPau4cvheakxsnJT7uHhLAs1HesWfeCGfo55VbdR
dmqpXS6Yc+SKOFAIb9fC5WFra3AOUXUhuQNh7xpm1sLteB/1ylP6SPLyEVc5dpXk
OHdtW7r24YuVCWhdeT8Yhccjt+UOHYq2ycXOaTNcUAX0H21S2+HbHsfayB+/qJkS
dU+ZIZyQxilLclwijIChr32ylAdNLM9ac/J1j2RPBPPLf03o9BDoFtCy7qM+z1Z0
CRMUO5LmB5Z24BghAFhsLhuMm+tN8NVG56kzIdJYeTDNxMyeDv9K8vj+fy5+4mNb
0CscxD5ZZpWueZ55DftSxaVeUbQkC3d5OTSZLWQyDYC63ZwKg/rhLwS/gp5pblbT
pQFJcBbrya/lvKcNM7jOGTp75vucCmLsLiwsN717y11unGSojJM/N2oEL/KweE/o
8AwVTliJH9/HMUgC+rE4Ne4xgUGhGxikCVe5Ynt9EvcY9nqurIyU8mn1/nBT9K+c
segUY80lRyzARgQTc93B+bQXTA/ywMUD77RJdCgH/KlavdwIRykts+AXNPkLwtWd
jczo61/0ZbR0YmtmTQbuvRa+ysY1fzR50sONcaNruUO/sVMyHn+MtIv7I6C51wiY
aOwsXt6ABD3SOGbMO+B+ZiWEKqalPjfr97bYqy25Ce/2vaqgoSpx6p3a4iJ5PZfR
UxpaKF01QHe9jG4xwLvPIZ3jaWdd/erZu5AxWFW7p9/Shh0E+R2TOVg+31MvyGQ+
a6ERELiF37I5hgQBWn6uEZApl25RcF1cQIrzSkM/0wxEiRBD7mi5KSoeZmiLR6k1
/kDKWeCPeI3nM9sd4BPg5BKHuyTb/AFpIdlEuclzr6RoLMMHsJJHvYZdbdoqIa29
Q4mKAzqoC7l2EukwyPFk293ihSh/Svo7yt71kDE0MKtVpPIoQxtoiVS9dkyx9EO/
gMrjbotd0wXRX1f/CjBpol4ME4zPehuBsTeWQJB1mX4a/AMa7a//dlz6zshL/VVR
JRHLKE6RJGySmg9Nvj8QOVc67wv+ACR3htLlEtsTZndHQhomBqTFKAmvf4qYoPot
nyTrNzeiQumKy5Dcfk39lVMUvrHcxQlj2zMJlGtrTBOmVKwNlRwDvQ8CIzjfHwVP
5ojM/S4O0Ks99FxyoRh/il0XMVbzhmczIViWIcRd7OGwcx48JWaw3L41WhOYuXiP
CLuygvsNRn1RwhN3j2XL/4LI/iq9sVQxpcyZiXbvB9NjEVI9o2Wb19U6WcsQjFLQ
pNhIlttSlXycdClQgiPzjJwM7Qu4/b8Y9+M/s/22GdgK6HFMSIYGG9KwJjK84ZAa
5uzfLzfbwVK00pvn9muDuG645F/TPTvgu9KlthPhd3ai3pl80bqZXkDxyLyb46b3
niCbl6W1XtMP8BDYm5Tp+vFEP1Ye3ya0sHd8oFXos48eSfM/wm7rw1aZw5rw2tSJ
PsgloB6N7SRRcQtHekmANAd5mTCwP1cMIw1/2YdNwAasrnVuCk5kxdoK0KcBFOpQ
6frCOp/sa/eOXwr/kUKZD1DH7BrenAvteHsTcOm8g3sgGm9gaM01mb+qgK2SwadV
PaPTabi3zI2PH8HUDhL+PuofV0n9Z2NTDMC21Mhz0mBIv9O5zARKINgEMiGGAvNt
JQGz7RoP7z3kooknWWXH1yKB8vEyxq26l4JkJlL3Ym8+wFtnBnTaWGRcDUOTp4Vu
vEP7SLiMvmHLY/7Kjgw0ElP82Baw46rQiCC+DaAWjWnF02LJ5MjQd5cT30WdTm7K
HrQnULV1kDhqzZL3QoU4kY8SuMkorkQWZelu2Z0NchIFl0R9YNzADaIylOxs07MI
eK2nhx1cX1lJ3EkDb44XqXfDMJBx4dhXszoh1kKIYevvGAhFhGxwrd2baKaq61Nk
0ng+Ng+eaL9+B8YeVdJv6b4SQToCYMT88aROrgJ5UeAnhsst6tknlIzUu6aXgiZA
WgDA+RaCOjRbwaWSRkc617JLJ36B5VTkix2jkwADFgvkPjDmCYQdgnUG1963mhmL
RkI1wGjZXbv1JJU/o63m2nggSfiW4oVJZsnEjZEBDcrHxh/6tUf8AdTWoBaHMX8d
jzBUzYY3WGIRAzX9SV8Str3iEPNpqg47JBMQWFD6+d1GPFHAyTBK8SB94yOQxQie
UkLxc9WBeeSVMKLuJnqb5t+8+LFDqd11g7WNyyLo+lYg2QqsFrPuD1ZWwMQKXtbj
nVSjpOolEoQOrZE5xt1wvNPiAn/1h0Vu50fCUBmrXuJxuJ8BiXX8aOmx4dZxr4Wb
T8b4/EHtqytzcE9nGka9OmcY5cp1y8M0Krxl8J8Hv0toqDDvAw1fz2Z9QoxRvLnS
d6fw1rkr2t6VGmPHSvLTbAjkN8a+SZvOJSQtPQ8Ua/05L4h5Jre7Nluepu92kscR
j8/0e4XOk3PmI0FX8TbRgcfwo9fCzlyHqDU/T2zVgRzOepDDMI48/kKztvm2VvN1
TXcbUav5d2Gg1n50GDISA6YAC06FV2SgogzSkaKevVanK8bjWd81LfiSTpHjrKPO
Moxnz4fJtKArxUAzXqql4mMNEdl8F6U+y+0/2n369nTSoNvdN+YKjjT2n93/Qe3C
S/4C5YVM7rTDS+yBroHeqv3kj2ucAM7YGSH/vHVF/nrAqvOIvtZfS8UNmYN1JQeS
HIp/hZzwMYmXqdPbkEmZeIzgkTZ82xE3RkccM0d2UxDtJRauzluwyDeQ5DqNlpmS
Ir+t7E6WKNic/v42t8R1wBKdKsDjLOXyhqgZgt2/X54aqbdsuj9GqVYkce6pv1PB
n4loz8bntOnaYmVuaey9xBykdkcXBgmwHgaNJ/8k3tn6DMf3mvZvB8BhZ2twJvjo
K1Ecx9FvvDj/mbnmrRG9XWiuCeS3yR1McadcYRzXPqxD7dVATVdWGiHA/pcbXh0O
0x6aYI5qH0OxF9iIyphZW5yXcFgq8mdZ+W8XOvGked3P+9ouCM4FQAoYdPx+3QbH
xdilu07ttzDb8rFLb1z1EoBpxnlYk8f0PwDM6SHxa50NtmwEeC2ZyFNGFtSKzMNa
Ud6b/rvpZ+ZtGKAe3P4+Rn5yyKiAN5ljI/WUzksNvK04IUfMPxT680Ri5bNtdeay
PAZ11hYsBaAPzwEjrIX/ha30O27xB/+CA+BLb/LLLCuH+k1k5G+Fdv6DljrD3XzK
La5CqojfToyEkp4ghSO/iOHGnA8dpWQv076SX7C93W1jOH9pD5qGIUsLhu6+Lo8S
+/B8MV5USToPyw8YF00kwInDF/3mNmA174QLo5Z1jtPsmvwp6CAkWQr0CK/nXlyf
V0ks5CzLM7tRNEMkPtNjE98CqvlGqlfCMFr0g3X7Ll6Abe84VQmqbZnQrCODnfMJ
DC8nvFBudS34wLaheTuJmAWNSnHPmyKbTtY4T5yVY3gRxzER2zHCLdI0BSXn4tGa
/wSrR7+lNG2bbU1f6x/pTWbB+ThiIwhZpQUgVT3HB+HMpG422BS5JW3FayzVGCo+
cfmdJmS6ZfrUatyS50WpZ9WeZr0Yt+J1hTFMLPJmZkmfz9D+GM1mGIE2nMZh4MAF
k5PliGULoDhwuZPfTa2al25WvYhKC5y/KWcEBXKzMUKJVgT/qsYufmni1+W28+ag
xHNuR+wVCirGs2sqB+pO5GcPlGVRP+NxgK+RuGOOdYA06JThMHPF+0kH5aSKVO7Y
UgoX/cqGuVzHmvqcEBqXetm+9T3naCwtPdeA68KWMco7Ql2HXkGxPMp/BWibZFRS
DN/EEtyZAWXBpUZdCc85EiICh6tXv3EiJTpCTZf06LmHycersmCiRJ2bh/YKAxJB
mjdjFuZ+F1tnD1kEmDJF49fSYCQtjB5flQOx8acP/7ZJOT5gLb8AvcL73BWc7i4l
cjtJabmbsyHgfXkPF1SSuTJwZvGvdc0/aHftmMVxqsEBEHFTQ6oidAtKVrXevQ4R
9rFlzPRRmj6PGfhlclEZ+oDw4D7/VUrFdjrUG7LZg/E7gEdsNfD0RXsSM8xPX78m
LLhkrIPqpiMvgTA0KvznrFqSEp96Im2EACKPC0XOPFmTVVOoYJwXNXpRfquLpLCE
pL7qrtHNNnjfzkw6KYh8iyH8ChvRpEQZrjmrJRC95RAlc6r3Ah7TGJqvAqsFSdC0
xcwdp5RjJb4o2VaAsaSsGymsJXc+bHiqmgKqqvu3H3u4psxTA17rqt/PM4DRDU45
8nrTS9EsuYcGFPdjxKAzDQ8ThVaGvk+/XgXl3/Pto93lhUhVyWHyoktWnxXWrPbh
sftvBwYhfT/kv5SiOMkCPrGebpcNBGeG+cMB1MkSZoskw348ySnfxsuSzRI22yV8
2sUSwYZaJ9pTsYwpaoouAhUzj+oTWRB52e4Ej+MbulM2cPRZ5rxKTk6gv3bBODko
yEua9M0dcK+s1aPPAjubHzktmDUDS80FO39+cvwEeTTaQNBYv/IDfYn7mPSz6OX+
ahqX3lSzjKDyPpUZ+KNGoA+mCKfChi5LremFP3xTtX6zYwPdtjFk8RGQy1QUmamT
g3E/pv3jnBi9cV8qGspwfZqueOAaB9ggudRjN5otYxuaUBPSfFIFq0JPc0jQwuF9
+phWE1LuDr9WmL8LjnVyYeRP2QZRgnyqFBOK6rDU51uUX11zbPgaKni1fjgCRsfe
5SI4FJco5Ypncd8NCAm22ZTMWhvcYHsIjVVsU1WCwTKruL069cpqS8EHXuwk6l/c
b+40IHGzpEY97IPZNBPqZPgniHxdTSqKvg89pDohvmMJyPoJ6o62GP/s1Eri7stO
OLT0chdPCr120s0RjJgsPrCNBeNbS3VJ843gKOawjRilufr+ukLpU32ZNWjcNBts
5cUQtCAmLr8jZE+5NzsuC9Vve9eIn7dqHFjqvOUGtnL6lZvoa8XblthAdJj9pzgN
/8VJy8VNRpNiQkadqTZeM2r07+r+/hoFimLu06pFgCGI5ZbPzaUgS4oCB5wn5c1n
VLgf8tJ2VXhP+Z8W9igVA+KaBQAqzfM9en7S9d97mWGiNAaN37i/FvNKDq7H1uZ2
DQVkcLreCYs38w+u/aVBceagY8eWSqOC6/9qWmYoT2NGMcjcV+QnVKVfL4cQvOBb
tf3XWnOK6N4O+9cRNc8d/6NCVuQNLBGHUPN23b3iG4KHuUXdgMB2eztZQGE2uj24
dCKRJBtFM8UUvzOlqIVVjsiZOLfZQlCuQmv255gcjlO9DB+iO2XbGhY+UTvJEDpi
KO1PkNwhIJg1PqULuyBV+U+LYe7MRyODTorlClVre57bh0NMCzuAHj/ifjzKypRu
L1NEi39PyLcDQlUH7dCZaN8rU+2U8PO++KBILWZjNUj0DePmiwB0YDgUZmfLIQOB
MwCFn6mjxfoawORcvGe58tgPeE6dUi4aW4nw5XWlj29pGy9A1IXJq2UC3NSDlIfu
nUFyWHDLH/KvmP7AgeXizBGVnp78GA2p51ckVQr9hQU+IktYPSYoA1s2ykCCSAdL
IEacrpKU3RFV0iJ0UxRbj0D4ZfF8EwTsXFHoCKtWA0bZrdL4c+fR/TCPEzYdA22e
tn4D1G6BOA/xwWz+pGKcgRLQN+iKDzLPiCGh+rrxXxpA66+ao5QfNnyMijTnEpw5
UVwKxFOeJxfC/jfbEaojXHWkir1FVxoaDCutTHvWBFOzpMELvKJmtsU0aSN0QkLO
sr7XMJofHYMsNQgnFSENCoTK9frj0b3z0AsO1G6dtBVeLTblpUQr0/LpNrdWVu5u
owV/wiV9Xg7xLrwTy6GbQcMDambsKLfQATZt/Nx/uzwYtoYU9sd6T69JhGiYEy+B
jswx2SUknwMrgvqJm0rLE9gZ4OamwQGTD02y6/Gb4GgEzTrbIhk5ZMZ4a27tonPS
gkuznDsaV5vze6bIjQe43WhLrk0gs8SPFmupV7hgpuMwBWCosF+69FgXa4ClxQ7g
7EybJkZFHQ5VoLz9iwq/Cew/dbVI6S8J3u5YFwZy+DjWeHVVx0eN8QpU/lQ6ALII
9aD/AC264xEHtSNQXxjpt4m2s8VOWTgT2J6crP/WMdp0b2f1DSisKVAz+Hi5TwHG
OgCTzhm9/dmVKbqGy9SjL6Yf9JBEDoDtIMCF6+GNidOPnCdo3ACaxmP7ZpwLNpxw
M+nfBgwm656qLO1mDmC+ciYrCgE9WI+P37NZH0l2F3wfb7aq+VVftKYO2lYiRK3M
uqO3BFpjStqo7+wsmVKFFowSyh114FZnuJ/qtinWbesI/XqqCoh9Voh0hkQVda9D
cR185I1nbip5pd7jLjPTZvP77PbkggmuLluQxzy5KC9wuKTF4NgPmvY6tb4yix78
gjGZL+xuNN6uXi1XyYIuNNXZv96KS3gJ/084ab/mfJ1UQUBIGvcPN5NhDTIdTrTB
GYcit8Xvw8SyvfRpq4/1fxIo1w1hYFTS/NCv1ir3vcwWacLVX2iVMnnDgzbJFuIr
fvdgtnClaFza5LVGSxkldRD4dGM/uRYmd84CMgks9spKHbrU/WtLgAZzei9pd443
efK2PGijHLNw3Vir8caHAX9WeTb2W44bCu2OJiOOd92VpDyxW54KwAXwydopUb1J
p7txycXcu02t/Mrad0qicqTMJm8ohzl+W6jCLKJ6oAGfQ+w/yTDED53DVd2/gzk/
OkyEDf5uHRza9iTETzPVjGTjBgVaGFnQzP5vk4DJMXFqVasmOIQab4fg9Qwl37yT
yV3CZzy9wCpRBfmzajKaZFvCbp8eDEGEgl+8UTbAu1IMJr7u79lq3d5eCL8dZIYt
Yj1fkEaPvaHqd84aEUIdIVJyRJC6ZU80/ELPhh/FdNGWKFHCQS9ydzpIk+9CEVCT
T82pRQ9f41zHxaF0QjYUbLSFuH808V37nOHKkg9WvMn5TjcYzSS+XokQolXPpqJg
DIgsDTtEO5xV7n80o0cr4C+F2PC4suTusgZJCO1vwfWkkU91+R2+SCm4wKugD08u
dmVCsJ5mewkvEVvH2SFJnTEnWgB63Azfzu3TxxwsoDNC6HSyqHOQGuh6cEIpUha1
q9KekqTiB5GUY5tzyWdvOTV4mn9hC+ksJxMjp77WAPRRxg5HuE4xCeIaROSelubY
mlDVgx/TRBlnQ4toYgpqBEnpP8zwwg4VNLMWTLOEHmka65xyYOhUtEdsYMgtK1XT
TYavUoYlzW6SIenZaoA+KXDkDDMK/6Fw3/zRMY3JOOJhptVx7/0URHwHDYmQQcK7
Gwb+C7b7qQAE5tn7x7rkmWff96kcpXUj9nGxiaxuXtE/PMqU77/dnSE479DGhjRm
O6W3+jnZz7nwU7vTNVrdr5SZGhgXpHf6joSTD3zQuOG6om2R7EuLb0OojhSl8xyZ
psKkN/UiK2U7j3AuM/eJy+5dd+u6oQPtpPGPeyGOvF3RlfSyK9NAffl2rhBhEzLb
Yh552D8UjhGqfvgwq4VsbWRtYBj7oNNWFmWVaD0pa5CADIf1k+Gs32Y6Zz0Q/N+M
38siOD1hWt6h3WlvmevwS0C1FBdJmNE95qKIZ1r0opDWKC2WbYEC5gNB/eXHTeFI
qsbwc2HZVADyi+2Nu1KIY/jRGOrT6yqtPXhjxFm4nJsqZpJwqbc6Q3oc8duDnAiA
70owG6Zbqgdm+8/hyNvDXRaIbkP9QLAW31kHDUPTxh/TxhXbrwmW5Q3KNIvdtAxu
Src0d/JcWCQgkRSkUr6DGAT1xWai70mW1B1l4J35qbHb3eozfI1y0CuN9Xvp7lS9
UgHVsjcJpA4JSitBiyuyBSxXRozAiT7gSm6BHBU2fjRGsT0cr2i55BZ0fYJ6qMLq
HdZO6SMJnEvxk4F0l6MOVxChkRaRsARl25QLdjzEYqCRueW2tZnX5H80nDyLS4NC
vXTCclqrSU08RcsLiVtylCKpUEd+PwysPw35xauouCfsg5rcJwNnGEGsl4iJOOPA
nr+il5NAlcMZn4QMwyNbAI826f6e7LdZQUmJVJShKkyTrG/tcGuXZHY/3uLxwG8Z
X3xFLHkcqoWZIOauP/VWpD36l9EiIkpnCe5h79XqYNglgSUSkQoHrVDI8HDhRC1e
ND9/Bb1Cj6MEI0a4eC17q4c8V8wqRC8t52Cuy0NGRn3Iu/eCz3r03RJMe1Xotr8m
F9GZh4gaeI8to+xyxHV3sdnYNlme5i1rGblN751wLidVyp+2I9zpj7g4dn2GXPCW
WeVY7Knz1J/HPSXm19XhRGz6pxiLk+SplmFBx0KXEsmtmC9QJrLoF8R82+3ItTXY
W9dfkX2eP2sQnhRVvumgwPzvQN6llMlVB2YvOja0yzjiOgrK3GSTqh3DWyODB4a4
bhlyOo85cd0ptv9racaQ9q9BET9d5Q6agvD5SYKL1T5AhX7lRUDitxkvWbevybY9
u5BNJjTaDj2xHO8TY68/eB+CalEONpfzARCKp7oRGy8Euu8NtILajgH6YV4R4bjT
Nq27MbIzh6QmJI6MIurT2yDUYpuNOZJ0lJ/MNy+CEZn2muHIU2zm/4UOk0e/Y70O
PSdUnhBNIIodjk6yMf4Wrlm5Jg+FM78fdA6ohYJutw9AJIBKwSWIJaZIKfqRFD2b
2CO2v6Qz8vKVwEmDwbR0W4zG3GOZduBemiIM1Mi9xDPDC2g2/Uatf4LWvU79JUYl
vkE0sVCBrzpQM09PON0X6Rv1SbTWEp2jP6Z1vOHajZUGeFd4s6yiqMEFhBGd51bA
cotFgOiWFMbbPg84t306p5b/j2bH7OflbPaT0zzOuIRWEcbbC84UQxuQBCjobuNL
blX9Fi0wg37LUPt3e1J7uzPXtzjYmBcxlo4bR3Xbk3+zSno+eHXNWuSMNTK2wMl8
8HpTN3Bl0q4kycBNL8OTMt0o/QpAlE6UoB55QnbwUFvQrZogL5ILEPoebt1CRL7c
Zf2+SElp5SunlVoshTqYcWPn9QSiV4sIu9Cxduoh21ztZUFQEzDoMUwFO/sRAPHC
g//D6H3xtcKGKDgVh3g4IjRt3PDFnK/ZSOwI5fCLnIj7j9zfVpIouLk+PpNg/5tt
Gwm2coYnQ5b7OxkuUkUpqKuj2KZULiTIseMVqX+QBptq0/JcQRWTNoui5YQh/WLy
zWHvdu65LhMfFiUKyvPajH/f+U9+VY3dyeSMvYTjuxGKG6RgnRKC3g/LR3CpBqHz
pCLx/z7Dfio72nNrOPBbbdLE98b37XQHNTOR1QY1pM2k0bLAVnZH6ywaGMTSFN/e
tf6Xz+pfIIVTusPn/8SClU+fciZhVri0leUIdyAKCKHy5S+zAamKTprytJd+Awo5
TCetgbaEeLz6Fsb9pPjHQVL4gLQzJjCsQRfwWOZJAgRRRdayPGaw0CF7HVTPNBQI
7jV24db2V+tgB+vJkzN97ejthGJVBpaNov8ScyRjZuFw9ZRkH2VWzHovqA8XQ8XE
bqNVNnf678b9Dt0nZ38vYCvMYAsE4PSZcEVdJuH1dWGcPedqXJI6QxUBLPM/T7gA
JwKVkP0QGq1FWZHeNXUqznLPnyHSu2SiOtlQdpxEg5f2PGxpx6bJhNNuF9ug3Kw4
ss9Pkz+Rmn9Qhhr57k5TxlnkxPhzLZ1Y6NE1Ck4sevYHkfuQXTUf/Y51KRLc8dMC
JVj0SHxwShIJmqAGnfQsEhSgQMGkmmtXANms3m++R0vdwc1MsF70CXZZlnx2zQKM
uhSUzikz40MvFVWCRMyjEGmttIeP0REzo2DXKGG7Y+z93fBuJlKdr03dQh3dsUkJ
MwLAQGQhSuwI2to+OFryhb0g6y4fRmByKdX5tbYycG7Ou2bZvWLogGhd8aROmdG1
NVHDtW1+MzR6f6trI1DpViKLUfSZmJJRwAIyrM7i6yQJJ2vRdFtz4XopzW9iHSKr
loHDb5bRTNaNCH8oEey/6P1E63ek8Wr/xtMIX+jAENQ4vu4kfLtBdahCvIr2PH4H
DpHK8IhGOPABS4CKBOQEfAqVQ90CFUo/WtpIKPWOuACXsGt+4pQVlfiJCqPQAwvr
KF1yxKFRXPk0US6MGzhghE+Wo0IVpg3i1UgA/NozhlxBajO1qZGq2Vpohqyd0s0O
mxnD5bHxfNRCB8+q4mcBanJYn9qLob1o4FvjdkJdg52RcgNQTe96cWG0Ow0v0nSg
oBZoe73sPzmL+Ch/EGIATFnbe8FI3ca5K2rz9QVWATRWhqCY9i7EYLaFhm9aLdiW
ln8EUoEulTWfpZUrukVFTws6d0MBgJtXwPlxnhBEqsPaBtoeX8aMmiGWBS+2MP5q
sVLDcEqTtaYxWSfCY/sM5B53oBzqJhSsCnwM59cbwg5/Fha00VJ25mCrM1Mbb4Cv
WKlJcjMpHdzba40NCikJXZ2Z2cGLI6Ys1GILMYj7+M010ztupJ6FNtr3Fmh5Hisj
JFN3cbLs/d8lyYDN2YG1I0mlzL4AkRXvUU1w1bDZMViuNhql46Zlc2DUFAJwJOtA
E90jfr6Lr8ke2cuARX0GPqnWFIvuBP9t+QMp3ub2E4tdIjNUo2bRXQvv1ctgDdBY
1WTQGGbzbnuEjkgA3UkHxdISzzvqqyi7zHyoyxloIcPIa6prC+1oN2CcwYDNetyT
9fMdOep+/qYoiKzOxJUm3ac9rZiCKw8mjBHcdXq1kixxApnbvjHm5mk7p3huTylb
0mCf/LLwDsfqZ6khuz8ImYtUVCF17epDdOLSdTqC/0+ybf+/8kRFEdQOJ9qVYUyD
+Td7XnkBgl1wfOThTJx0DkX1bA1z7QYDk6Pdm6EdPL6DatBo/pKUqB3eLqm/32gr
bvBhdLAO2L9y49EtgSw5FuTm6y8E9+Inx+gFK+ND0TX3U2dH2OGvo1B854hjM7ac
vjU4rLtS9Kf9Ndu9IYEGz6LBtMEalOsh3NwnpiGXwhV5fyqUgt1qMkVMvAKPMVWa
jxDkmwT/ZjBHaJffFo8focSJFlfQykHsiQ53J+dIu2IuJ8x0ETr2g9h14fDbo0iy
pj1+D+6Oo/SIf+AOvWz8uykAtAt6mu/wqpIlaYSet00hSfUTfWCloIhYN0LCDhgp
hv0nUT/Lg7bDv2uYV/RsKrWrI4CfYxx/mFZvNpwtQQZo6ZrTwkkwayBxWLMyv2P+
YwDXlgUimzDEA9gnnaVnvfoM1T5NvIYSvrXe+7bJth+CpRn6jIjSfjcNT2mZj0S4
L8jDKZAYKhjt+v0ufN0Xv8Sj6eCRp49Fj3jZrAv6NKxZlhF2i4U1RGEFbPNbjSCw
YKnoeH1G5IffTnCQ8thOLQDQ+m3G/8DsDkEBBjZRR98MY4r7LhJhmlftwS32ulb5
0201KK7xkIhBf0GUs6HWa3g4WJ+oApPlGuxTxjQP09UtHQkjw+UNRZjxZNXUv4M0
b61MkMLvGRHKPaeLoAaLgfi4XF+kf85LeqiUSr2bdygJ1ErYt6+KF4KZw6RPJr1E
B6j9CrEuKvUg/rMHoG3XXX2m51dNnMa7m26yUyB+DvsBILCZcoEATd16ssi2V5mv
2rp9oP1fwuy81aQz2EU1dj1gDmugeQAb2J/7g+rOz0fN+sFhqNZ4xp6opTM/iX00
+qjuNvvkJuG4PZAJkmn9wt3oQoLx8Z1GlsgRT2fe4FEHjXAU8ysYdmZGpiEHuBU8
UxrXa3QAcykmpmSWA8/LadlhQgVphrxWSNa2gQREsLAYToVeUCbdpHUe1/uGJj6F
oUpGBVF6hjhAxX2VemWc1NkrjoFkfbtx5nLRhNs+WvPCsCV0IkP7e3xtt1vL0BeW
BKpXyMn598f5sqhGhsb/y78Bpz6NZh8XyjK/kJtLU6KRCHRnttOFL/rn5tLpoN30
THop3C2OEdaajDXew2MoesFo9+f+11JdPiLZhwGQYaVBz+JGg9hjwv6hNBUgd3sl
K2fRSWu31ohZsvbvAzeD660b0lS424yCIDFttwK8MIRVWZDLW4XRrq1pAdsI7Esr
dKj4HY/7+S1bqsZkDaelHGpiZ6Hv7fG7HpMJNU8MEHOZ6J7vyctsFBQtZm+ZCJ0o
CosE1AUpYBvp03BIdKMeJvDlZdJnm2OeAh4xqFf+O3OgtD0v6VaC+LA9V1l12D/0
9+mSaHv3xVRn2A8pB2rcF36RmcYzvSBx66l/DlgPsOhVRwWUFenYFN76n4AoWgvh
Zd82/SjNvLY2JT/itaTdNjGm3/4aTLnfcLFigTgtK4Skp1rA9UdrcC5FQ33SaIhZ
09a+e1ZvBh5o2zFv4SpRE4YIQFEBnnCpguDwNyMhlGc8lzwNTs/gbKFIBbWeoGuF
XeR+s3bxN8dcNxdv6iZSunT31hbKW//VUd7qI/cjJjGF6C7FpzbRzCHMf8HS5NF0
lMUXVoacTxIag5lKhujGtEq0GkYIEZcKizcwxyduMSASbC2v2FQ0uJwbM8vdO+wy
OTn/ZQK6kVIbl0p7xgS9ghg6zU6JCoUddBpMaxc8LMIiKk8MoqcptBIFlJb3Q57F
Jf9h/0kLC+ln45lYrP37x1IDnZUxDXlgdPPokX1iZ99mtpHol5xteqcjRDUBaN/A
b+aQHzRqceAIKrdFsrxI5hSGe/7XV8nCmpzMcdojymlgvuTW156gJw4r5FMbcwrs
SkRbaef/FwNPI5nQCBIrztqf7/Fe9XLXizPFqcdrLUB5YA6I52K6FkF399wsaMyY
BBrZXDCQa/YpoAKgS2FO2BbI+OtB51B5YAKdnzz5E4nOHXgM6lMKjMNRW8CNzEwW
4+0+09GgQkyelPtyr48avP/myvm2UK4uvui7mEou0X2n0JwdkGVabqywMGk/Hjqr
EhyNO7ysZaPqy8rmm+h0eQzZzy7d0oV0RPJfBFEth5+IBCLbMFYkJdA0++BCvLjE
TzEZIzjM+FwDY+fcy6pudcSUfghJcC10d2HSIJXSspEEMFRZbyXxv4OvByG+1FPj
ImCyfk9o3aJYbAYOp6/4Y7gwIS70MNoDUWDEEwpHI04fcr1OeT83TTwXmGYXGI7k
E8VukYOx0/P/wlHJxSSpSdEHnoNa5JtHIsaxFCN/qg8ZYl6cyLCNPf8LEMTa2e1Y
UgVHKi4iImg9sL7oGw7xSo5ROHmzw6tYYpda/dSs1yHSvu7RVsNzAI64RKO5QC/v
upgtLNoQpn6xcz0rSUKHdKR8H8XMFpuVQUtsh5u0qrcox+qusbeI9HdYRXK6IBQF
6qO87NteMxO+1Psp9OBUAk6SPPfFCNuK+yw8UGwgr5KvgXv0n5Ctn+e0nbea2nOH
w7PnlR85YcFXcepl/kGC9pOzqXBlGUa3aJ6FPRC446t191DU+LukAIHB8CZMDQvP
Sb4rn1ktYFyc5L27Ru2PxHrOBpsma3BXVC4Vjj9mq32/ek8+MEUpnuRdeTmANjZ7
g5wLyN89RSj7Vb95alwsVAjnKLk8Zk3FJ434es6JTZ/jVry6QHzUSslV/vFGRPJX
x8fbdexa9UzpXdJDvSmTSrPnTO4mPsCtebyyqAcMSWxqNKEP22qh/AbJNWP0JoME
Do4AjgriqpwkXFFnEK8g6wfq3ktMGYNp2Wff8ut7R89mGXWnd3WfWDHMGmy/a87T
`protect END_PROTECTED
