`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypyO8lL8dyLyGsDxCNBpM2qOg/6MGxbDVPBS3H2Xp+JE08BhsxX3dbZeZaFTKtHN
VEM9atmXtUyjK4QziqE0U+aQ34YbCcAyCEslFHFXTBGQ5/u8fzZ2Nk+mmWItOumf
3fpokCaNLhnl5J+gCgKwBnJX6PI+lPzXiPgov5xnPSG3/xiZNdJVKwovOis7uszq
91faeVBOHvtGjYpWhDBc6fnUirmPrtKVqQ1Lw24+lqRHBzml5ivk8iK4pmDVrszK
JllUFHh33jQmpcgmJpLy5R4sCySl2M0DtRDUvMoqzatqL4RO8Iq5RORB5o5k03VK
2SajJsh5g8WmFonndsE+e+b8AGCzwtuEaG/c7+LsJAWcu+/u/6LhFsvNtI2YyEhm
IPw5o0qC8O+b+ZMMTWkQBtu4cQiwWn7o0K5SAtq3uhTaeKNHVwegtGizMrHE1/B7
vMOb2dHqFbYy3dYM6jfg/w==
`protect END_PROTECTED
