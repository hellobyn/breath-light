`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmSq2P5xj52EwekbcM4UzTGc8KYKC0yIvEAXNSefsPpdehQlLas1P4mTFLFmzN82
ntQpm7nnm4BHeQj2KY+BBnfq0gnbkZL+9++cyuhIFIuJKVZLWnht1rCeiG+O5u0G
M9Wb1nUvdD33eVzWDmE0HGZdTshiEWorwTnX7qQkwNezxn4B7ucPqBO9mCCihSMe
gYSm2E2RHgaxkMX0FUCwXKECxFUJykdSA6Ocq/3+Xx2h61BRigAmfu07Z3/sx8Qb
ijo6bXzE5hME0gnHftzfnvl996qwNFFBGxWzKBekrdMZE3eriCosnd47cDgeU/wK
q9zrcRY2DNXEEOYfZXU18h0z4fzl11YsIOTK0uKBS0bGxhrJluqPwsN5EtLFskkN
CVz5e/BdvfpbQQuW8xTG25lRKZGDuI1jJz6AYzg4w5YR57hiDET8wqiRDK0jv4+e
J6KEeR5cGB/OAzzLdVO5zG/IsI64T0JMYC7sVKV2jMZiLL/E9mkFXUcg3jxjTnXz
UpLNRHXOu4tpibOUNi0Mw+kO9TrdmnMSlJr0+Y6R6pNcO5ogSAqREd9eTNHiSf0v
ecmX/UPx4JVblGpI7uSOG7uBYDIDNhdJcddRfJA4biTXJV3vYskxqCYW+VqOVUS0
8Cs+R8AmT3t8pfSJIre6LXBmbUe6/mhnlKyg2WW6ZJuyXSPtEIXlx22vd5gyEa+f
JcD5Hx1WSdXDA4nhN4FXlb6EjecXeek/oS2Soh4ON1OZen5mnINwGq7UcRTD4Bl2
n5JV0gdff+HmuVSyHbiItDTa1GywVx42JJ3mgEdC9FeM5ZOXWITuj/5em04b9TZF
sUHnmaAzUNxCrGQlfthnd1ZoXU7NSb7KFGWPeODOzHlol7ulSly6pZjqFZT1q6sE
zdx3zUM1MdWNWRgwAhBdclKZV2FMedg9onrqehXGyIKtv0ILIRbygPz8tAN/MBDt
RB4D8Q9IaNt/rvswxTVMYC1zFACvOUNdvh803AcwrTCyGTbZRV8j09h8HjvPuXav
c6l2R+aKl1lukSF4chYUQtRze2Wy9BTeNwbo48jDmTbKPCJSrYX0Z3BriIN7WzLI
8aRYNEVe0/FJ9IDXkf2hYeJD9jPxYwudnaU3RcsesjGlN1QibZoWOsA2Tvy7tYG0
p0w9zMOacMr/zRzpjntRHxOqxbWN5+aCh3VtyTzWWDHj1WfDG8LuVlSMu861QvDF
xsfECMjH3K+Fd90lwOuX2PkUsHRnLHMhzTQGc3FBpTauUhoEMNekr3tXU9BauLCV
lF0SxVoGxkKozrB5pZa4di0/LY3FWCqWILe18f1ke9ivikDHhSRJwLv0uevUtBCJ
CudfYXylcniHj9FiJFo/1mUMqxTeHTSRmKtXs9ZCToBwIby65PCjmdY9yio5gBTN
IiKhZ+p7qHxYUFkDjegLgzzCFQ2HN3d0Iw5xc4ZUrls8c+qLWGdJOw2n9+BhGdad
mhp5X2wwrcVCxshOsQGLeUP3A4UBmPvIBN+LIuc+sVRfeMh0bGU5ppjWK6Wew5D6
Zg7afnhT5Z/ewlpKwrx2JF1XFJVsmS9BV+VoUEeBr9t6ewJ86srqBKKA8jgUoKPJ
BwoLaX39WyC8G5adUH8/j8gxoiLzki7JnAYknZ4F1wM4hzwYnBuQ9vxLZns0vpQQ
uZKi4yOMqsjtV7qicXHmdsULtJtWQY18jXqoWA6O7SGp47W7vPb5MGCLVH4MkdEu
77814Xgjn4khwiNDO95ef4Uz0gPAX62Zyohn/XNcTUkkNFLnME3gQX6HJ2F3hX05
tDei7xN0+Jjj3WSd5sdCYx6JrmWZy0aGgIR6AUHxkiawJlUyQZ/fgTpYoEO6LWoK
VMSmdJ5xEsvh8UBPzIE8+rDtPiRBsXCyC1fvxzQBkJjMjxrO+P/YOiplTGGmGvpw
3ufF4Dpp2ISAa5DnxTxnIdJEm4OR633KGiJQ+cRQnTE3//cR5EbxNW2MygWmYpzV
GlpBrBHvYaLJGC9AU8F8U4+Ml41Ej8TW7qRxNQwLtUEq9Yt7Z/Ey74I9f0nMOe0B
H5GdOU7m666NxBdC5FfybjSG2U4va6C00pJUuHAvv6NN1mfpjraKs2UmlO2N3+ks
FPm9xuThc22rn6vCzkkRqgWoVY5BpBgjicCByDtmZO+HsrXwTCjjgXRGZoom+V4C
CgvB5Y2IasHo6UZ5snhVhX/wGuhzm4uEdnYUKhPyC3lqWZsgNdSP6c1mgUISgZR5
KXo01bxRc0kGSNwFegTpYu3lmLbp1eDs79AFxDNP7gjB1yjCbv6xJKd1dcpx0FJh
1zcg7YAyQdglpfiX12Usv9kd9E3H3yIgx6UOOaHlhPXGn5iSZ8bVFxsBsmImgfWP
gCfnPnuhfPfKjH0cTxGXxre1FM0diuqx9D6I3CVlIbTTx6JeXlHmPdto9ReuH6Mp
`protect END_PROTECTED
