`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nfh6gX0z+CGM79MUACoNzZW/P89UWg/pSMU2+CRBtMjArX/p23ZiCxaVtU4TAzvw
mzB2zRNT8jj3TtGCXLFLIDW5ket2+frgA11Cai6HqQq3urxQekLY++oELfX+fCiX
Yohv3OkdfLfNJ+IU03oKIts9mtUhuhwl6QcWjWyU/WDpTyU14rkAgLaOz/othAs6
WSAn/KHKPtCYVgE6ScE+RZ0e+i1SX6eICJKXds9vNd+iZon8K3B1Z9HJXeSaNVvD
v8pZJ9zkfvT9Z4J9l9CTrZ9WHHO4wfvbANIljh/3UlfLPL1G6tGmfR/E06hZ5nHS
dCl9nahOR2Q1M6zMzz2wMXNOtlsg1W5XUC9PemqXevt43J1srvREzQD8BJaAxIsn
qnxfPHkA5tIrBcGK6hQ1IA4GTnU7CPfZBIgda2kP3DABW4jSQz0OAc6DRwShZBmS
zkT3km87g8v9Sfn/mbkZWB3Ozz2Y1D4kfhFDVB+WutigfhxONgtECZnPsyaOTwrf
vl/gYd0wqh8d08wue2Ve8YUwcd+HP6GRSuT2QqysrryNVkWe2xoGTZBtxTIITeeR
djrTY38K1WgOCH3qu2gKIyU1eyGk47vUz5p8wQoTTQ8VSTlm80Sx+dPBDskNtpHV
fJfTy3bBvkAOJRBqbclJSpyAOC21UCHcueqwGJTHzzVYzKLFx5x4ABbwhp+ww4Y8
hpYAHxUok43oDi3PZZlwglBZFdl1i/vfBrxDi5Uoo08NXVcL4RneSX2qiRHBw5rP
UemK0JFSVOQ/9+EAqpSvjryby91AXjzcrx+n+S/k5z5aZXcb24pHBqgiUEohh1Dt
1EpmVCdHpWuOULJoz5OsRg==
`protect END_PROTECTED
