`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMgrlfyNRsEC1lknkCvw0P2Cevi+r+mroW58Is64qISozDHuCF1wUBj3mhxe60pq
mWYhwefkWaDsvKMVvczOVtL5PYDn3Rt8c+oTgfYLjcpO50fqtlMHSgqvosRIoSdS
mvimrhuM4X0vzN+1n+yaMwVTfgPR+UgLDecPPJNTJXZ7UNe50UCvnxmIUoodntgr
+vARN8XV3+hRgM3IotipgOUX2cf+YGPx+bvWloO35HxwnC32uiODPD5oaHGMbkCG
WsEviLKlv9r1k/M1a202WLlX95Nk3wlHgH8YoolLgucOuJNLZTYxdxR0oLnz1/5I
cKAXOTmnz6VESR3WDPCPEpYJ+3lzeHq2OpDYmY94e76QCQwnKgwXwSkzcv96YV8D
zOENhEL26daqn+bOYizunTtkHDDh1IxWx70t/f+UlMcG/yPevpVFL6vPbiuEZptm
oQaGKjfgqbhpweuMnHQKu3bS+tfAKhBtiOO137MFdTtT8kFUSdKWpKhmzT2LXaFh
gCzsAeCOWPbwiNNoxnvmkqcSuFIZuP0E3n/9YJLGfyhvVhNVA1vvXg87UunCCTYD
DzIxPpz3N7IsRzqpyPqSFG14V0jo2hw30/Ns3Ufv835mADK6Jbsx2MuhKvtgpLS2
IyCb09hPiZeSW04+NyaysxAuHdPoycR24BJ74bY9EhFqjyPje9SbhDQhhGCsa1qz
3NxDHGZSB0vMkarP/keK+llAWaWEPpZp4RCKcrATA+T3m/Jsot9O0v3bapmQgvrG
1I20/eWw/QiFcFhr7G3o6s6nzhFM4rZMW+58mL9+dX8xYMLECfSD9bWNa2iFjABb
Dqo7botCvj5Usj/rVcUkBRyKaNrnXzlWZPjQ51E083esfqDLN8ecUcBT6NIJ3Kdo
UrAdZfhC7AleQmOq7v4IxHJcmJtfziQ4v3ceEf58db4lZs49klKvrm8HcClFnZT/
akcGm0x4UB2ye2uMpJ8LjM3x8Cog9zgWrxGX7K/wmn7hwh3VErDBqFXfodxho8c0
sNBuH7u3hJLm067sNKwiUA42lBq6mILstq8dKpShCbOPA3KyQA6x4OdmeLHY3sXH
QWPxIzor1SjrGO0QyWzL0m7HsWgRodNACw0Z0tzzahc+89WGv4UFwRaID79NOShy
63QV//28qICmeOh9M3t9bknWCTJiYUr9N19fK/faKaIpN5CnHuLC67voPLB+Jg+n
MNuAByBCdOUYd9peXrZzx9cMZcfmei5uCMmKDk+iYqSEs3C/xmltkzCGzhCz41ZO
Iz0ZQnISVb/NlmCLGmVHadbin77ttfbh6XjkGETXMFwKeCTjAqOYXCY6/LZ9g+We
6HD43W2rzVNi/GT6tek3xVAeIm3uN0tlSX4Eoa0YTtyzFNlGWghBk7oZfQjs0ACp
bbtulIeH4iDda85z0SVVi8PehjGEIOZ0LX7zPwkgamsWHoh5aVEpH4DBIYtv2xtZ
SuiH3LlroQe61LXJR27O0rTxnP4G35OZKfq0Mo3D4873XS8t4eNq066DwBVUvgZB
WfXyJpaVkGX7gnq36uJyjkKzMqoizV/jwoKPRNSU5PHlum0A+2o2fHmVfY6ulQen
qujfBjhVyxVDpPi82FlnECmmsEclf2zCRgtNsikhLDu1lva2gF8XFmsLBfJ8WKP6
38fHezy4s2gASkFBV+fLSw0BCtP3RZN/+Pw7kwdc+5w9nD1ukf4y9hRQNHJ/B3w+
PSWeBk53za3qacOiU89jhAy9CweQ5M+0YBuZJvI6qJo6UJFoGt/auwzXUlpZsDdr
hs8Jb96PJiYqzDLDuL/pleqaHWisEf3qA3HK8rUTYDdqfQ1arG2SAtPCN3Q+4C0z
4ML2tTVt2P/Pj9uUwaFzSUcwAIDxENF4F7qfZoraAKWwlwZOKvtIyLJM//LxxWWk
rBbAzjS1D9xD6EjQPDHMycOEWjRtRKAVrsbr6MX45aYLkyotLzHjGyJRDqZPNzbM
SbpfPGi0HPyTJqmR+ow/eqNFL4LehJty4XQtf4Jt5xB7UcS53zq8sa42Ek7QzrYP
AvC+BXwuOLQi+9kjz17WAVZKtQ+5SCLEXxgliXJkDvXqKlEMx5dMi7XzHMRw2sgW
4ZyBqGVnF8QyxK2g7UcIYIr8hPf78hW114ZXYeEqNc+KKcUfu5BCw9sZam92qu46
iojDa6jcislx3RVG+wJLb6o5CwFVvVOABs7VRdFOxG8m4DcP4uxZ2Bis+mljjc9e
7VYsVjqTcNEHFKewge6zAjHV3lY6QSe/01UTADHmbTco6Ckhg8c6eke49FGFBUk2
0Zc6zreWxTlja3vJqVymANeA+FhZJ0N/TIXXQee+05F9ORh5SXxRmO+hr2d8SsCl
5iB04CrPRgraTj136WhH8x+PtGA/8OYTHSBYUxFt16wrtB6/UPKCtz9onxHm8vby
k4UHEl9fh6iWWlFQVsmDT1cQaSM7l5U1TxGqEXrJqyUe/HUsIopCuL5e3wz/Ib88
uomtQcqY8ATFxHEgyRKU0/Iee/PjLwXFZNx7AaaT+SopwWsWH+8Q8eGpkCzwmxlr
4vAGJ+JTBAXtyIF+bQhFnbY7BcuYBZut0p6FcP3SuAVSysF14bYMB5ZOgj2/eL8Z
thn6YlhAIZAGqRz95zRSmytgG7a5eiXzK51vhCLmZ5S33PZvEmeS74oJfqlKp6Qf
N9hKXswPM6rEHcjcQqrTyQ7N1Sr85uW2Ow74DP/VLxVerlaj+Kdzrk/LgnWhjKV3
gSspiHENecTfwKoEw/pYah2RC+Sd7z3boS2jrmj4VuThMGoheP9atsf1hmKK1x+k
P5mY6Q04itu8fw0ER1DuFipFAWtkPvt5m4jcba0RCFadCEjqxEsEKfgCN+8KaQJ9
XjfSeCcg9y99hqeRP4GUmRIXZHTdn8WV00QPlyS0DqbGTG5GOYkySIoPpnpNYzlJ
/nH5+tE611ADsbj8RL30X7zk+X8zwmHCtxee8YYDF31d2tYM670XJCdQYwzawS7L
f4wikcvZOIY8lusmJ3FHprqDcMuxAp6evlwiutkWIbOA6ZAEswfDt/jcV0IBo2EA
JHLV/i/N+fOQsyzwVl85SjfcX460oX93wEkJ8XadjNlEatyEO4djMKhBfWkON5XH
HWsGchk/fqYqpz8YLLNI+K1KOKbAr6yZxQsbDVwqDphTvJzn7qKXA7lZHuEP8e75
VvFGlKJ9qs4mbufuwIQho4+qATItvMsNnUYMbhIzeA0xvZo83cBl8TDgd1+xZPiO
Wf/EhRlzbKXG/2+zN72bFxcCAGYof64KS/Gebt3pxoCcYVZ+/Lp9qLmTf8UFm9q1
BlYMaboPnfcBRLTDuncjTHQMcAXR0xisCOWvCKzojZJ20StyLIPbLd+qV5AXWMlO
TDnkYjCCiFG4x7ZGuBxthRqf7Qj/Vo2gzD9gAb4XLwgJSHapn7ptfX0/bTKSV3AT
8zkcAur5z91+Jw3OSpmckOqhlkbxPJ5PpSm2hcq2jGpgXj+GJ5Cq8vNd4LNcgdAj
TM5EDZgCDIeXUNDoqqG0D1BuZ/Lyo+YhtFqv/BHU8XYR2bCMAjOZfYokKNnKqmC0
fTmxtI8Kt83OyKQ4kXbspU9goWt526SqXYOStkW0pR7mDFl92RXCZppIn2x83bNj
GZyZzWm/GTgym9ipsCWt850NF9kfAKeHjYUp9QkjhJBTORuLnUMP0tIzGJq2Bb3P
WMjw6R4rjRp1MlmSG4FEA1WNdYYRJ36YBXK9fh3p1A/ccVkme5UOC+VsNnWV2rfy
CiIJ7ZiFwBQ+w1ldL0NXbnVOqpcTCiprG9YR01GTBQaE+9mHATQ8KFtXb0ClztX+
tQHwqQ5ElWeJ3hopNbUS3AjsWtv4v7MvW3dblXv7MFnf8C3Yj3ItLIa2++M8iwLO
LLFyv27O+76Fy64sPPzNRa25s3dmSxsHNXNLOA6vjvtldhUvmxXjA4Ykby802N/6
sjA6MIqpZJFcpOwu+AewFA038yg9YQN5Y0Dgz5m5VbnUiYmVNjcPFhGrVmE/oLcv
PWy48riPmqyQSzt35Ol9H9AgaJZ5mnGrhoo43AUBV8V021Fs+LTuH90pCSkuYmn4
cIqLYACTla1ioRIKZguMaU7rqLFK2EBH0yfZIHDlqfhn7s6ARZb83M+ZopOpOa6o
YZoQf8PTBNavjznHnKCBVcUKjrGA84QVYYmaV4fuLa8agHsz734mqhWuvEEkz090
4lAnBk8Yjj3eyxTHMXf84vs0lMufIRtsrtli554XoOWTMUrNygSmp5V766GvQPCO
VuZUfyJ1FCkScPWhJziXb9h0CWq9R7/WQzo6AHBmIPl5kLfDsbFakImyGOKxeb1T
2KsCnvuOa/+66a7Rm72dpfYx8jCpXD1kF1PfPaYoXkZWbFJSt1p1qaduvWxpylUb
BZheMJrTD5RBYUTqKsvkdArq3IknfPwVCukhemfWPj8Wh4mTiD0x6YG0lPtHO2Wk
WzBeM8fPqMa/WifBsGl9MjmW8IgvjbcS0G3uFMATIMv8o1XozUqcLEz836V6J4XX
FQkCcds68gUrst1elgLE8QNDGaYg1EAYcwXDPnqyVRAHKWrYwG765XD4c8opI5lj
epbaYrKDpQVF5zI5dUC1sI1j059vJdplJ4XeC34exOFaeoim40/BWnjJ0aT0qyBq
mcnAKK13pgk+hSZr/68SOgOsty3zUG4BlWdsxBM/UCvVzQu5WIgj0TwWf0r/FvD4
hP6HXgc3q3RNMm4pffkEDN12GfRCzVrdCrXIBKAuv4D+6XH21Nel8wROafs7JKUy
i3AINE0yf14KeapcZypvl6J3hD7UwaovQDPMSLydltgjv+eCAp4d+HzgmSngyhoP
mdeHla9GG0zIWtgkxIKC0MJBpK5lt61JC8qgll/Z8QL3LNLAUshsaaPQ3BobEJ5r
gXJpR6z8loxAJaz13t49BfpHQHIqP9+KybRt+MGYSxnLNFx0+Q12+RGU6G7PiNFx
lJ8hgN3aRAjRSmlpFV5tuIiG0w8YnHkbX5m0eV9eWf8iziX3GGX3ASXADajdEmnL
t/4xgnkA7m8pVMwvH/yxFX4IBRwhlrd94QZwuRdGDsNfDgUI/L06/nq7hPZ+qbt0
G+N9mbo8tmLMRZWdfg0lGZ39YcElreG37leAMMBHbyRySCXqy/8COYsPGHU8tQzz
gsv0ATHOg6JAFxdNXZbGiXjbab0PBM50qHA93y5ljCc04Y30rz+Un4o42DrG/dWM
v3CSy9opn4p8uxrMx7dSCdeFndPx4GE4WHIhG10nF9DTKCA5ETmOrNPjKKFMRgba
NXBrityF85Dltm5W/kRcWBjERF1c40L4y7ixEd3tS7V7UVjlI8xMhJMlq9IX6i1i
3aItdG29ZO6uy3px3Zmaqf2wA/pfKq/x5PYovTqWdWNWlRWF3tojEd2Yn4Uvzjky
pKutbzpr9KlS1pRg729PZnN8CSyfeYwZqL881geHkFu9KmG2AezU6CVx96SMH7Jz
SHf4Hrj32Rv3xo6KiGlLfApzqzGriN6NTUxWUIFm7jV2oOC9ZbzH5lmXT06hGRkT
uNs93SGZ+6ur2ivq7GoVsZD76Gt9Ri/tcPD2B6MtAaCUCmVWJ1bnYZIZhhOj90b6
OQeAVfKZNHp0NqB2wmP74E5E5wkhEdXiYOfVBV3N1QsvaGxXhnifEctLxgbfvjXg
g4AD9/RRiPNm5tHF0QKOYWi0RDWpCK7D/0dh3ydB5p4uFB9SzBdQbs/UcVgSTjLi
Hw1x4TAeW5C41jvOhpja2fGO925HUaqqps5bAbJZ1hizlkIN5h6+jwKle57OtfcG
FpsP2WE0T7+A9I9IXPByxjX5quunmZ3Kz4Zqgd2IHDNSumUc7s7VyR2BArKTxv5l
CCmfTzQHKSwYLm02de9BtjFmq6dKMS/i/sgxZnlyDkfKA0YX1+2+IlIlcqt5fOgB
4j3IGbkfLOIV+XkYVtGeDNYVkto5ZrbzhKNKDny6OXt82N4PBRnWI7iubYre+nlK
l/RbrtR/5PUN0a6z4goIOdZm3hhZXs/WENrVHnWyghC529d+rJciX/B1teuR0cx8
5p5qdcwHb/Tu48bvZNfdGYavMv2WeD942vGBfEvBBSguaBHd3DdV3w2suoVR26oj
0u5loe8t67lm2kA3bpTU1kmNPgBiqy9kKdq7d6o2XWEs7yRzQtZfwj3k3gC/CaL1
EiX1atavX5srtLLmQUody+7H/OoPOtsEHZ+lsy4b742TF1nt403QFkhWdT6IEBXo
0LDJRWGoKYyvL5iwxKBXgwKHH3/Zka+oQmONVy6wgYWY9MO0N58TKS1oILSY+JpL
QPd41X5/Z+aaZOPZSi0Mk1CD267wCBu2jaeZwAwtjACCzIJ1wd19jH0uhbxJkWoz
Bj8fhTJNKOrHU6QPqDi++YV8MxtQmAp91fbUpQ2I2Y4leG1zduSHnf3cUhPj+fFN
vMTq82WMWIsFQ7uKHymdGu3p18tx8KGiy1+Ug0u7WRmlmJWWfbqk33IgWOspVm1A
95xxDIvLlRcEznq9LmcTMnkVbyeX3mJDdFyjsKSyLJ/rp9GlafiBTX4A8V+1Dqq5
MNtEV3ZNqeW4OS4DpYjiek2oMVpkK2O9yYYJIBALY5uW/oeSAIAM46CouwJ+jBAO
Hqof9aHA3xw/zmb7GfMXwDQTddBpZ1QjFWF97h3C4wh9hPJ1Ld5eau+0UisZTgBJ
K/nh/douImkcttgooIwJFHDKF8HmoGZK9qWLfzTxqpw4HA+w09a6SrEEri3g1QF3
LeDAS9GF/tos8nwS0T293yGuxCZmj+lqbhalkJdqVSnukI5VjwrL8b9fnbjMHXLU
DqAMMFALwldBoHdRw0XLvSZGU9uuqPxKcC58MRfdh7FTLYU1JB1sOUHIsdIn6RCU
3uOiyV8HF83ByVD3O0ckz/lqet9w9RZC7w6yQOyhPD94/6BNGOcTldSAsl+s7Oi3
`protect END_PROTECTED
