`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KUXCjTdpnhq+j9tQ8E9ltA4sqYev9vjtbDHk9RGCbUQgINpV90VH6yKOdJCehyX8
YkoAEQzZBTnaxOiUogmFAOcWQb2IpkvS2p/MPxQByy0slCx4u3Z/ZT7QwYWURt2B
3z/ovkdWKfPWSIUNAXvKp4w4SpkdsLz6cAK+8JygGZg8A2ugBXExEKI8N9jvVDQG
DAtMTyniHKSiwkjV3ze6zuD10S7AIWznZnKYouazpEPI7ASUChO8SAsuMPh7B2ul
VUjexlQfeCL/SjMJKRoRLO0dQk9IWT4e3Ijw1jlPW8BUjf0VlQw4dwM8v2pq52Na
uFBkWLNLjuqByfjeItWqGEbIEp/nBUcD/E6qreWnPWEtbWz1g15IoXOv5jL7ItUS
gp2iARdK8lxjCB2ef535tE7UhnpkTUANafGDIp6lCVauX1rlB9BThcyCM7JnlOr1
tkAQm5K+VSxGAsyAcMYxEdgnIP+pnLJlgzsBrcFrsAOOG5h1wyap+NpZcY73xWy9
I9izZ0COpiwtpmgwKsaoOCRvbfgEz0wNbBRUdgfL+Lfy1MUe7ELyZM8++asNO9pJ
EPk2cVFYPv0vLfBJ08lgThcxsO8s6/oBogy4UL/gaSoHmIS50+k4oo3HhtY0D//6
IbEnzqZWGL1xlz6Q+jWveVf81OqyH3ooieMJEIhEYvmhRukTDE+2/RyJphhnYll3
8qn/gXqzs1PaOz3OYwL9xp36bH2mwAxRQttu4gL3PcXSuCMoystiYur8SudvkqxA
p7lyT7Fa1s/3giYden5mIabXxib6a6HD5MPyWaSPDMm2NGdAwPjJS220tzs/lL6Q
/So4/nHy1A+CDLXJNF4vMfLKLB+U4uRMgtYKjwMd+5eJi4FZQjhHR+wNyZIw2RNy
f3zkT0vXOEYWtfJY1G2hNwqYpJ0hLi6fRwOcX6rJa5VI2Ahv037c4zllZ/7vcqO4
1AKzR1bwmG7ip2fKJe9MZrp3z8FRtplVOafBVkX7PQ8lbnBSuv5EhZqlvNMniclm
etK5KU1zsW2nLRvyIisLZKZwzh3NTQuGqeheXnisS3oYNj6DJytq/H04nQbQ6w5q
UD9bdrDZ4xQTuM39z6qbNlRpLCy7JgQuCq6Sjlp4tVf8hac5oMGeH2PiM7x4ynkb
9TFOvDsEO9ZRqbvrLBPriJtnwKYBTWlKxzb45aboVlq+tkn/rv3Qki7xb1LqBJqs
YbcdhPeJOPmtoLUIRHhcSat8I1Nxwxpop5k0gu/DYoufUj6RKMW3K9UFKyNVrIyv
lT0cbGspSZwIeudFuVjUo6qn84VERbt3iWnukNpOZI8DcP/yIGmHS2ILhRf4KjVL
pzLDWtLu5/WMh/VF2rfWfqj0eB3KIfuf+J6rNIMczXw3QHT3DlYeHfJdzWOgejVv
G7u6CbMPEeMr5AbHdlvFRoiMaHiS6VDsrvSugvkuCFWRBN/6CLpmBc4kzKymYKpn
0qhsXQwS4JpwRQFaZa7eD9NXFcoUHyFkxZa/dxOmShMHI9WSTrs50KH01yMu8Khz
ZxsRfaVKoZSVB7H5N8+lfomw/ELX8N0ob3bms7XfWK9AL5/zq8jxs/TYVX/mC7B2
faEjSreGyROf7kvGGoiCAm3Ol0jMeAekY4U9F4kbEdsNV2n67nrBhSCq7bz9/Kz+
0AFmX0u7iEk7+g371vGIEhbM1HNWFgErMkgS+91IoejVjybdYM+D8XLIAwHoyti1
5p5sz9pDiyg+tKz47nagFR9wquNfuohqQAfWrWSUayhjC1mUDaum9j1UJHhB9lnd
sMcerFE57GQjaScFHgjNklzDNR0H1inAC/WzOdnOhO66HiJG53do/hxvdnP//fR6
Zz0ymMZd9Q1tqG3w+5OFFdkHRQUPn7avlgWWh8fuE2D9rrRuqEbiu8Tgc+TyqCCO
py+7zxzs1DhFtWAfou49gA==
`protect END_PROTECTED
