`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66zqRy9hnRPTE9vHSTntprOzeBpVSWxF/ctXFESRhhZ+71DOpRe7vb+b0KuPRc6X
8eikPLJctvdMT0jzZBdvzVDPwTmHk4Y9y84o2GZDlTM1y0YBzocN1f94MclhqjzV
LGssF1ywC3LXefIQdIYwIFfqG4OnubRXswdxTqFY+iDXG4b3bCI/1cn2Yhf+ZssB
9wXpKrXzGXnlT31HnrQhAfuvNsAHMIyeSHTbXk2+YnhcYTKatDQ2K3aRvt9Po2Q6
mDDzhL3ZDP0Fs4YcSxoEub0jVdMLOc6LfovisU1zVFhAKUJ9D2wi7GgDIn5d1gcy
F2DVekiDRfUa9QfWYDTtBdIumeRLhaJMpmJwDS+8OLw0JaSMM5awt+y54teO3txG
s6ycnfcTVPXdbOEWodnHvT57+SWzdEQ/VGT/d6UGaYxHKe895niJyzTp4tKFWp+C
ptLYf15AiUspAhDFQYV5uj1pEHsktuq4qfpt93yQZgjL1UuKdkNko98Z5Y6NsyNY
HBr26OPbRmDjPcpYox6tOIHUGxEpNElsh0/C0X/pmxl6TZ5Oe2O5ruEFJU+rrGzT
13XlzNk3Yl0t//8x78faQWjvT5As3jW9+6eB380JtsVes/ERHLo2+4ZgB3DuRAL1
0SwqOogMkrALnf827qC5Qt+bxCvUfiv1BSvp0IpU+nayfh6RDCOVudsJyhi+whjW
L4ES+Uo6kB3jy7pqi07sN3siYXwSAp+JE7nB1Km4tA+rdpbxb3SsQYJivyI7exhM
EfSR5BlTKI1Q4+eL5NQ8KI50pN02ZzjAysO6/nqzv1t+UAOykG6/PIqtBWcMP5My
tKVjUK5+0C2kvPd3FxbCT6fvHindCQuUHm56oLqy79x1g0ZIcah7fE78lho3xn/j
bolxDLRYinhau2AZs5O74XRMtE9IMWn8Eh7MjaBCf7sL3qRgCeHlTcDwgO71fas9
IbjGQ0f9WBY2QfsA/yMVsed2FWuMyLLIbI04jKSve1WPfgHmFFouS3h8jd6dxfAd
fZS9czF/A31s3revCY2ZKcT+dma6FHzsvOmOhTTnhvxkKK8j7oQbyRaPEvW5Lh9v
3EOljTorgjL5OpZw2WvqkfWd0fNXMYi7kfMGYbmpZkCh75lQzNoiBPROq/qxaBTI
QMBMHtxvfQKhI4CIM/8alcDc+X3xgUUQRqAqQ0PoUPifcNFjHwGhDB0i7TcIkw8c
a2T18Qzd5Sc4Hq4SGIN7Hok86GQQ0l6YI1KW+edWIEezyU7I2ng4mkR3Mmdaal3M
EDip/oJ7h7l1zM8Xn18hu2m+arObGDgANvSqD3V0rF3TTLJSn8pdm1j4S/Pk1gaK
VKdK9UwH0DaBh7kLkZFwbtg091nczYQSNL16yExLbI/6mPuvsA0soUXXbaPeoUID
62krV1kXI7V1bRLO5IfZ9pLPJ70e+fm85zI6j9DjSNxvYLz5NoMmUt77T2xSkc8U
wwutHPSOQJN8ULSqxlqkP8B1GryVh/pmG6CNGQXHNZyq/6Ho6o2jJG5kLrznw5cZ
K0kYwW8+MWmtVwkkycWX16qM5/Pev12WMdLWiyxQpKXt8rwlsd31s4OMok2bo95P
Yeb5MSQ/EFwnOTsc3YmfJpaLlHypUiP9fidRna8AWVJqWChUC1FIgzeseNUUawYG
lWwoteHq8GY0CFLKoTFxIjYH+ZvTQqyORQqfn4wPoE7ZWppK/zzmqmENiGRayWvX
qNQYjmyIbM/F3GevFY0/gyAFk3ToNOScVE8lraaYXnFZoiigQWCpCMoYPosxGw73
nMj1WfBKQZsnvYQT826N7h7nlFTkYwBVgvu7hZxlE5c=
`protect END_PROTECTED
