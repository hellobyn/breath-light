`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXkw7tNfLCYNcg8Da5JF8WPI8n5ZT9ckdkbnZwKHBwGXvDSKhAjPSjgIzGmZOgkn
BrW3YO1ZDNZGVMxubpdcWe9izEvj914mtM6M/lH2DZ1FD4mK9ThHOYo2rYFYJGby
FjCh9dvsEHld6u8OmGatC3V/y/FpwMwUthVNLVMwz5tbUS7t+yPS+dNJPAkflLvH
ws9aTUpD2hshPi7snDo3bpH3+RNGrUKw+NdovlmLCkBURUJVvCaZHoe5lMXc9IJt
vxZczxf0bxEYtDEzzKo5nTzkR3gogSatdr02YNN77pwEtBSeDjllJYihEMvsLLnm
+cop6x6DjpACITzCGdylD0PJtPxJTkwUgFBdu6bcJxU0ysR4I/p6dZ/LjuifolxL
V/B7bDaVh0C7qnoQvHot/OAhbKHU40u6sz/0Yije9xaljOf1Qojv6F1DaEXZavwt
dNYLlXm8KcQwvd4KBQHAd7F92syiTocahVyw80Nd6VXQtOY6zizn2kJSIlvlzkK7
ZjE+NBH8JTn5wHrDD55lFQ95xmRdT2f0Ac/Wr0D3lknARvCxCAxFos0NwSAHWp67
54+iqAGPGyDjU83k3zvfVlN4LHapd3ppLfypt8VuuQ0kSJZ/FK8e7hMOjP3F5OCL
3UXHuiGGyGS0hhXzbGmwuJhQazsAcLeaKEUGocUsunrVC7iXsbdB5R3P7BQqPdyd
f1W8nl7Be0MZSUGu/W/fRf5qfMz7e9sUh9ZZp4jNvh1Q1dIuiEkm3dPPM0p6+ei7
96kt8Bk7frtzDxRlLsrMPN31I2KEZe4DGS5P3r8Bagvk6JUD5qa77QODfk9gF2mC
`protect END_PROTECTED
