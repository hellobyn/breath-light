`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/tx7GRlPYD12Roqw8BnxpZxaOEQTPAFEcUmmRsw35txkRG/u5agd3o77aoldLa1
xp8c69xLQAslSRv2KMUJMd1Kha0SsuvkFPbiUHXaDTffsXSFsToqKhVY/q07CmNP
T64wTI7kBcfcZQZd70RdUnA90PpZ5zlSQWQUF+RM56weZaxrj6bJA/hY73sPYq6+
rkUtPZYxKqIQYncnyO05AuRyqgFUww3KYqwWFzwXlTtn/DBSjnwFUyxXa2ZPGecJ
WSgLCwimUfaaNpnT0z5MdfJHvaRdrBUT7BYTYmultwkhRVJiNg8FlDz0gYMi5KFD
rosRwXR9D2iksFNvEg3T/9BK4d83ACfS0ptYwoSwcX5gVcl6gxHufZRTTFr5BfK1
j6ofDFK09YdjurVk9IvYOXMUiorVqV1vcV1JI2IMIsvLPaCkWoV/KFSWfl1V6l7Z
QvuQjwYWxIl1DvHBP7ZojQExTZzAETyzv5PYyuvS0s1nVcxc4nmO3diUDcdqpXVo
YEfJcS5cMltlWJlJ0JUIgDB7B6c2tcdh1tZRy+m8uzF4ZlSBYhIWpOSmDOjoN+zT
B0I3ngOmC7DcjJ7t16qAuw5vq3JA8LW07oX3MPTT6YNHLF8J6ytT3baoL7pPVNVy
68QozC9l0SUtzA+8p1ES1ORmqkZRDLPuXBiQ/svaUrwyjA9/jYHYcxKsIxYk5GzE
UFiyWGbWRYiD+3lvovSQpgbkXWpvRmFw4wrayPtPVJHKAy7Sgr4OeBnXWci4jI8G
TVByLhQ0N6e3laKAc35pbBJp4n5SK/aoBusruwpS7rP3a67+lXU4X/iK0i/p++gG
BcXo/FMTw41F9HEHERcV6ShtV4mx1jXKv4qIJy2hwIO5LEwhte17hHrSBM66Cd2j
p6vCIT4QgWp9VR92Hw/eacYQkiDI6q7jnNGRBZ+nbF+LednrFW29xMeKF0eGDuDN
q8CUyAc6RYnCVo5TXVOy+lU57OVaR4dh3om67BdSZAz5rfN5a8efV64dk+/oOeKb
8/nTGMBDiMr11oFnOoTDS2CCy1r5D0BKXtA851Y7g83ZWHo7MLJqFdTD6FmRUkxM
Xh974aURf+mOnpT9VhAbi2OPDx+6C+ZyEuTW42cFWgHY8m4Tw856/DyajBR2tzjO
bkWDZupLY69AU67bZhR4f/VAqNTudXgKHiOe9fP6XfBvcWL/y1XA+yfuL6YfLXe9
Nyx2EXz8tdsheek5q934+81ETUpDImeDjWCcWKmRkMT/i+tK/3e2a/sDmbW1PLel
06tXvrxsaZnU52hSQyHlCuo2gGNsBEOeIpwswmJYPXNPhGGOKTqKc88DSnQ18+VL
leTjUYVx2vNYaIfMZlQBFRfZSLr7vyNkYGafVpicOWRx2tY9J6sVn/yCugt24E44
QcLPdUI7MV7nmWMPm9NbXC1lGrpy8X2jfwWgeTBWj2leQZtVvQ0m15xNsTWgIrVO
qSlKPMxghzpo15NgJi5iUuxKMKhV6qYUS4M3HEyqHHI2MkMYvS0pQib2jHxLz5KR
MpIUeCe62glcC3a33Cx34GTczo/lUwDM8rqs8PPR0fALgcXR8ow+B5r62JwE/5it
`protect END_PROTECTED
