`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VqxTyTAU+PFyoNMWSclVRafMTZBmsWnlb4gvT83uEohTeuKRtYGn2k4sU1GH8wk
+lE3iiEAqR04yAAtLa9HlQznoj1X8ejceEXKZ8evFMEx4W9l9dkUowiQPlwntBYm
r7NYzcrnkzyCMUdhWTwJ5UxfxTr7t93ast5bEPdGYdlZIa2llLXiQkCpTFY5ShXU
1cs6a2zHQNHZ8f1JIf62KkLabCGZnE5xCBTqsMh5eCfjjA8qNoxvS8V/uzeyYfhd
W/XhFGoLNwdzqimbcT5kx/kOxZo4D39PbZrZ9yZidZs43/B7fDaMLtiASjY5WGQp
n3LxPK8GC3ZRmEn6aU6oWPKjIQ8hRThIkuurtrpzQ82I5hzyopwNLspQ/FnodWHp
58zkHtf1rRHHKrD94sAkF61H8zT7gM6OboMME7co/h55A5Rpd5uk09p5EBaynqeZ
`protect END_PROTECTED
