`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEz3k7HLKB+dLIqZgB33Dj1WyjXPRwWMMF/D97j/jnqm/tvqoaZtStQg2GN18vHa
UM+KdpSyGN5QWjM/ykQj9dqkW1tkL8hEKhoRRs4QY+iwsOxYWtfukpBpS8KgSuzn
P3Jgwo0rl7Jbj5AXhOgceHbDKsbDMpeuvcOBLC2zb3zbi95gdkw/9u/n9kTYRcIh
iaVBXybo1VX8aP2XdD8hhapNiMfuog+cgCe5zZgPbyRk6y7B9lVmYHL0TNcwLpeV
RbNqS+jJ7g6fSxmDPouK9bhY8+sjzuAvHhTC49875X2JWmGPi1+yIC9OTV/xKdhu
stoFWcpItJSv5ciBMXXZzO/qQDZhvXOlLaidFb/w8wnuGJOxl7ie2KYkJL6z7RKu
kfEZVlpxitLC4RdvuQht5SDl1iW4riuy9+IUoprpzI7nA7WlTtbcA8PNvXWnfq5E
bLxqkOpCzUP47QXfrGRp0hr2ND3RHb2M6KQP85is3B2E6XmUdmPD4tPzxZHogWh7
ROEYnzIxOmZh6ICC/F5dnCXzEUjmKZrfLdOy9QzAMxlR0fYFAPs1dp5WkTaT1hBp
QrDBlOKebYRhYtWDXvnUqP4BJt8slSFUaJd4jb2X1Shilib7uWcjP9j4ym5LjHNB
sAWHZlUPVR+59aHIgz0CmA2A0x5CZRYMjdD4r6/nd71bizT6xzQn4zosYzChrt3D
NKyl6WLQKKd4F2eLNUuanocUpL6eBHiAMZEIMbehNWIVsG6AkpptJ/FaDymNYygA
5FaOK776z5yxDQycVADXkYeCqOll10YZ9g7FX9pI41lhubNfje8HI93EPKiKVdmO
9AWDDR4JeUwTcxKTJnMVexp6rarTVcUvflhQsIfGKdJQrkjUIsa31WtfwKFwiACJ
IXUgBqhN6NFVVHCKAuGuYP+CnUCKeVz3mruiQ1yxSCm0TBI9X5X22PD3Ezdi1TO0
a0fCXrugQHP2+Oanvbpp3XuYxsal2N0O+KoGZgn49YE0jhkQtkvCuvvQJbEjtgfF
+boMc+IsGl/y/SwURwRDCc9kMZZh+k35iMOQKORc/+f259JhY1osEc9m1KpxHDE9
riMUbHRpKTuOHVQ2UfAuZmAcUOk4A1VHsWq5+MUp+cEUOCDur63C2/hnCoMFP9D0
mSgV3W9WaPP8StS/GzJHeA==
`protect END_PROTECTED
