`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rYymGZWI51/6y/NK+g9BmW63HYGCPIxSeiyHMEfdGVPWNRSx1ThMJK/Tw9p8NrB
ubNIakA/GnZPn190HHhpTrV2tm8vfvXHie3OO7sXNYwnbRI62RdCIRlhZ5xhcVUH
CvvIJAKUUkNXp4JvLHl1PxNroNqIrjZDy4XGnsPh1p0rgVe9SoXvL9K/X22AXESz
ZEuT948BXz6E2mzKsN+HS4MzwozFpG5KVVIXHqdBDBFq3B6Y9GyIO37dCu3POehK
eOiOsBgqQScdKHNB+VRlhxJNrYwOpLmM9Wnuzknah9XyTqGFGpp3uDcBWyv1VkuP
kyaLlrVMgHKk9R2U5dfGqqR42r0O7u6GFFE4Oj5q5MgAPR/kceWgoNmgyq/wjpPa
YVoTX4ve9HJc0SFW7EhCw4qPt4Ou2d4rczWfPD/G4+9KfDi6rZAPfBWucGNEEg1D
nMqnxwZUbjkSa9cOinGEj98qYMZvhReN/xBHxJZoiTJHO6S6PufXlVmkW5VUONTk
EKsyYeWRaUm/lvr9GNJzYvHe9QtSzsuW2alQbLnirAH23otvgypK+ia1YzKICTnD
2ZB7zRPxtCA0QZ4OQ8Pv6D8dGtFlsc6WMKVa3owMotAwPr8Oz8oaNWmIr3dkYYSe
EXnfo+lzrnqkTrgecv9FGT6aEled0oG8MhIQGfy6NwDfop/lx6Wn42bmXi+p7f83
zHUQb+86dksFY908djbQIjQcPo71q2pyppZPMgLBUFuiOhHEMulhAgNiM8+61I4j
lebvtoYx6RGeiR002JIw8CwJPzPXk/TIAS/leZvhu6hcvWPh/9Awxa8d67xtrF56
H5DbE2t7jTN7Xc5d8/DPVutIGGK6uWNzmyWZtZiMs8zzL9JHgGnKjcUGd2oc7Gir
6kQtXnD/fyFa/e/FXC56Ov6vY1bEMr8C4WDNijpUxicEPfaNZBWFyRqAXEk+qqk0
ai8/vR510VB48gohoWGBoCYlIhFm04YZnMJHfWEdWRewdOoKyTgBnpYBOr6SbqMv
UpMOknx4EIm03mgXe35sPbcgHQujvmR6BiAfqfH8kA7mgWKYsLI3NlTt5ACWDB9n
Bh7j8mwaEM4eWEecuV5CvTUTq/UAcvi5Y4Xw7SUHtBw=
`protect END_PROTECTED
