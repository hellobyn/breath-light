`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
APYxSqlHzAIqSDzH/V8Yrjiwk/BDlN7t6DfS2VfO9QZNQ0NYm6+M4D7fpCGHTJ3K
aXnoVJapajAz+j8b5nf4jLPDUh9//l2LuOBQSEiTub1hJMeWm5Q4PyubIaoMLZ3E
IHCOaGiCsTv11OTj5C4FpNsTbuf6M17MucsXryxk6h1392quvsnb3SlPIQAvQiSi
hGn+NnX0TMfBOHoQnGRql7fshlhtovF2qcavm07zHUZjaSN74RLbDX4yas+zS8s8
0cWw4WPqbO9HWnIYNyPf9EVQCkZ9uD18pnQCAMe6cA18/j71zJGeNWZ9kHmC8unM
JZyCGyBR6M77cB52wRoXteOyf601/oVg6meW6rwBdLevESLfhw5QaU+J3AsvTxle
rDrlAhUXF0fiEf033grnGbe1l5WXKLP6gF4J139D+rrjBqq3T2OiR/Q1N9/VaOI/
ruRzbEXhD76ybp1R5ctrYv5O23t7/TjDeaN605T9pcpkGIS3ZFhJlGT65OpIMQSf
VlAT0PkXZgXmLs9drN4aR6VDwaUr4CWCnWILAfu9f3rKVZ3TPP4pTh7k8bEq0/OQ
MxeMnxuO0NYhMCXZETyU1GYXUT/PP3O5SVuB58uetDYb1OiaIUk7Ib4xeISVqWnR
/X5vKw0hvjCVBr3JA1fvhdBqARjUE/XLnPjyPtbo2Fm0lzSQoUGuRayVceh6TOi+
d3XGintMV6mxa8hzicZess5hoQcoZoM/fZRW/q4FsEixQdwILk9CkAIPvXdZVARY
mpMSxCQuYxXBNJgB4DcUJsqgbdqYfNtxf5gnJaoS/AyPMlQkF3qj9WBKlDGzlZnZ
F7knMbkEwRyfGVRLKrForsZqXbYTb/4y/ku3UYhDODx+Z2mKibCKulnoUaw3DWPi
DH/gcetz3wrIP3F+pN9XtOJtN2E1dRvlHuAe+H8oCthhsFIpJpjXtrtnuxJUagWE
AeCEbgcXpIRjZPgb7rnGPiADQpwDhnwR6TWRs9KpmgQ6P00mcvhvPmWgp2CcWx41
gO9wQLyk7k9ouBRsIKTwFRvTTKQdb+LoVi3vR74tr72nLgIBtSFIG3yXZAjZbf+l
iDBYIy9uB7tU4y4BdAID+D6TCGqUzejX59H/S2Tljfwg8tnHfTGZQgzLnMWMVJeS
SqTpVEN4XXclweV38BiglIF3vESmJZohofc68EYlhKjArebZOCUFhUad2sS/ARwS
+B2B+rJftWLAVAaKVIWgrZwDyiq6sGIY+wtsLnAMQPyXNp5WPM++tNy/cXb5QUXk
QR8mQnQr+Qkr+2vxH0U6UsC+knmkaBjdMCMij7Cv1+Ppeugl48tbbeCg2JhhU5Q2
HAvmfLQfkce40E6JASqgRlKwMGX5px1K+WrNywH9BKdmgdPF+m4pBNb/DyNfTigh
4VpK0JTfsZYAkwpvdVcaHeYp1Tcv1KdhQKQ3bfWEKZfEGlsPMcitJG0jkBsCK0fR
VbUNU6EOPD8XmdNXRybAjebowZQq/4JwEbq8V9LY5mPXN8pJFkQwKICKc6WHv9m+
szLauNLDzrduL4mjyPzeJaLefbVaK5YQJ/DdD02Om+DRqJL+peuJGzjvvoANDrem
F1MUA0FaO2aIIH6NDKd5829NJtzujqQWglrBSOQG8zEX5ZyfJkNMHTi9mcyDyS+E
Y6BXd09zuO+ZdQdPlKyZ3UbGR+xk1q5e4ioStCE59SkzMXPoQ56eHtGA9g1e7q9i
GugCr3Qqc6QfCRAoLHK6voHeqaYX298eJLgmKJKAid7mFJOg4IbLymByZ5SnY/Jw
MBtns3hdPq7beKIykyJsOScAflfvjgTH9J5C+19i5wsEg7tS9w6ubFEzyVqf6+//
zEUhZMTud9n4KSjhI3QRSWR+0GmmQ7q/8o4lcUuE/ZJIj+gkkaDDgSemoy0xvp9w
FHPpFpD9mZdjMRcM6tpEJKMI5bpMWCj9U4EgqRlKNK0zkwKjBA9rvEw9dgfj5h+Y
JGVnht+0knmy2YvLeDAJY/N6riHKBOh3wR06jdJyYkrOSzrbXuKxsPfA+DT/P4rG
ZrJl35emBOry7/044owjJfakVwpr6jRZ/VDB3gOELEIyCoHyyNtF0yj67KIKhyH9
4Kdh4Rx0sljUcHKRF0IZBdjm+MML8FJMlupdEtHKF1pMDXlVK17HZ4IgSQVth7OM
rk0Dzdsr3WfjKRXBzFC+hSguF9BM34yO7A5ydaD6fKPc6FF625r6V1tCSqOmc8oF
eHRTmdYa7pG4U4LJHOTd+ZZFnUQAUTJo4UZ6hnINXtl0kMj2/rANNh7xKsn7hyMC
/oDDJg2ZlilFUx2go30ykjy+K3d1zIaTUnSjc5h/uFoogqtC5zaIH6vmeLo6+qiq
p/zI/dzXLS3kmdH7FFTH7lYinKGbUJO4Aq2PnAkU78aHFBj09vNYLZkszAJzHlXf
vH2i39T0leORvlpCpI35njzdsbsNK9T6T9Y+ZvUKL3fMKJXwV0e2ZtnTvm8d6FoP
/0bIwBk8UB9Q4O9/xHLcMT6SDAiI5mTgY0O9JhyQckGBt7xHwU25reDvZdp1L0tu
o63xLgaEOIYCfNzw5mTqsI8XU8YfDga27wvdVvPLxS2DP9Ok1DqdehZp9guc9dxg
U7e7ZH9JvZmFNFraWh/pK2MKqar3d4mPDiEPOxTgbHedzJlcPrcJuyHnfx9O7Pb+
bahhAS49i+F0vJHXFyVDR7t3RcrFTufjvZOhtx6vz/F3cJHamSr7BGUulW2r6MDs
1xRJOMP1DPqI/kX/nUYBgN8L3RhmjEK1SzXZ+7OLEIb/8hUlAOEYbDawRi7eL7lm
CoyL/VPnNdwAP57A5Z/WrzUzujZgra32tkclMmoQBc9Q8sNEf6RxKMiMt1w/hn7n
xR7EUDKImUXZBOUxvqDmbsZrUUf89w3WKxu9raxK1XHY9j8cPCNnE8t7XzPSAPT/
3siaCei3BY2HEVq/TEHkxB2Zp5UNQZ3mH4P+WpmD0PatgNORhLmWBLA/xyl2TAO4
AZTOU/u6MBDy6MxtvwiYbuHTGai7rOtpbPDGfONpq5VPCXlg4alCT8UAmxwzlkC9
Eqck7OrgdzykEz6YZu+Mv/rlkJXR07jomnePLVvb81eJaV0JWX4nWI0voS+vQYxH
GRfZFIbVFxat2foKKyilijIjEx/rA7C3LwYcxONLEx40La9nkZy1wNgL6MPhuIvP
tZ9PbgWubfEHna6dogGL/sZiaOXFrOtHn+FLUPfUyzO6A6YmE+VFVXGrUaxvlo0t
qF7t+MO63oWjUm1hbJEgWNLsITXGHrFoy5LAlEMmjO4v5Yd3HATmP9XnqHM8b8zx
ZotByd40SR24jrwnJOJBIiCpby3h8dbRwIxHmb/66Sj8pHhXT1RJcuCH8B+bnmYQ
6PAXO/zWnkeddM4WrOiMi+Ey8/mgDIbpG00tKt8i2NibMSQLkwpl1X7WoKdKDyeQ
obJ+LpEbOIYwXm8FF4eYD6r1HYdRVkMk0ac31HaOEih7OVpZaVKBl1F6GL4WhoeZ
NEPUS9zXWlUpLQf7oXH4HE1eK2ALTgCH4RgfXFw2HKcOEwv1dWjtePVKG8BF4k35
R/6TyOraDk/scx/OHZGesrwEirT+q5XuiNAZiYTl/kY7hIr7BAgWaAem0u9iYZ4L
xyK6Ter4AWWXhfy9g7cxMr4BuXmRiYDf2nw6Cr60UxZsSKKR2c3wKRligpyrfWBJ
SySPTjxeZVTDeLwuh+GHxTqU6Pq9df9gxjOBPJpxRZaxliagisx5lrPqofqA6PpW
VU/jsttmZfYfZdamY0fxh6NXUENeTWmAXuKal5WwmpZd88MBVRd+UbIG3WEPyUBQ
FVMwN1WiNccbAve3UFQd87t85faK1pLT741rFwMzlnaRKkW3ADLHzkNZCeiRiiV6
1Fd7CPYz9UT0gBq6afLLsvSyVtcf6No5WCxv9F06PoQ35QlDeX0qDjpEk1LS0wzQ
wxnCx5jPitbVXLZPxhim/rw2UjLdSOLJ9Arf1z+zf3bm08NhfpOjtMMia4jABe7M
VRMufYK+2FVhBxw8bTnSOoTNjJqNXE1C3HihMLWQabG8NAnXb2ZBWTeWj0bRc7+U
ZBEEa0pnMBQbLzMjsiq21aBCRJpda2xYqqke3WEy0pMzLr0sIgR7uR5Dd0955wZr
+Ad5LFfoMc1N+6/8piA4HnWWb2/pe1piLyT2aNegyx1Hzh8zf+Z7UwobNuACeSe+
gvDTse7TtapxM5RjSq40zNWazBg0Rt5dxeKsiSzxPBsORclXaYq09iuRImveDW8f
axSQvC38KLFe/mMctiJ3MQp/nY82ewDLZn1XztDssuJgdfrctTo+IQS4eKWS45sd
5r5cS/Bko5MBPCKJEPTbHYUq8AFR8qVNV43IOMbhhAsJOk6uyFpaY55XlLsDv9ag
tIe11Ygn3egSCHimrRnUTuEOhg8h12iZeOr6a348tWg3JNAhGuJzAdJXUz6rABSF
uhBUZZULchFdfEnQ9734b9mVukG8YBh8uTkUSVBTzdxBIVEp1y0GTGPQHxWA9EpF
S5jfgZkk+25k2VHKBYE+hVW1GnyyM6HnXhd9lymdVgrGzV3Eah3K0Ki0nYLg6zBC
XBAUejun3t2wvi74sTJwGwM4DN0RcpSJE+O9hoQ0mPRy3AW/mWxhEmJQ0Od+ICnl
qkRGPbkbpigKUBehH2oli+d0XMcTyD/KXItHkEzaNvI83rbK6l+lpbuTVVi48/E6
8Bld3ECLv1AYikJ94KBxdmzxsA1CEHO/DeLF4cepASfdHwhhOFI0n+BgE7fXznj5
Ti6D35fy7n7fYbWYOoLLtyyWTAj8oibNvmWB5JVPuxcY7FQlaUOYZTxQV1HEQPyu
XMiSmYwW8K6ErhDrrgQle310KOF2n1QIaJhDYM6S5PmK9on8tF4BpM206jOrGgX9
iGGWzKeAjJ3gkoXkiTCyrjJL9vfZG1D5RkiPdCzXwB76bJM3CVVLLYZngbE9guC4
sMBZLJspkMvPtjO3SDGk2QJwKipLbPS94sSGxl1+jDtxmlemOdsU0Q8P69InJjpy
sq8e4Y35NTLsr73KxOST3OFLCoucenuDKPIBIc2EEkSMyqnkpS73lVJIzkLmK4Hz
srRhEnH2wpZCBxygS9KRRKr0+FxTgUW7Wm7Sr9JWor258ASJkyoPHow5GEgsldQ8
LfTVDyPJngJ30RxxzzLsL3enzJHUQevoq4H1nRIMCqknPEa8DUkJ7wX6/HrDDMZd
dy0LPcKJzrXrKdX7CqqIK08bKhWiPbcKVE5JDxaiLt3TkkTIjWWYg41SGpHd0d3W
559tQ+YIH4CD7wgaX69AgIPEg3RAzhpaAMSC+YiyvCu7WS7mKivgTkPtV05VnXWH
OEnNKvkdub4EbdnAT7uBZ0qO1KfiE2Q1ZMVfxDBr2VdvO1M3To047adlWf1Nktzm
ERiTeOYG8G12hhPDS9biLM3p8ucI5H3KnZSBUQCOJHVf+j6RYLq0XZHzH0Dq+VNR
8xvSqupcJ5/lxvDVt7mzN/2I2sbCMS4n+LfELH5Wpf3K33on4pn0xvgpwCQVzAt/
Xb2OWW/JgSkPOba75c+TrgE+w+Y3ldusDIFEHSSyHFoi4PdMiSgbQfnQ1ETUXlhk
ymn9ocfsX6mqvKLBE7GYU84eiCwvlP5O8QLBkukN2NdOhJZDMyBeA1661nY9YLQ2
+zhFebiTqgEv38LBlBwo8RDm0oo+dufRSU11gtoNvrVsBWBsJBHdcJbx2xft9oWj
59D4nBRRYdEvJlICYG4QVyJXXlx+kRpk/8du0L2OCbb3DCitz16tyRxJLHiYUvSs
AD9c2T76zvNEPhEi4qOEQVK54vvwFnxJABUjvyxmsaAIbMwfOHNXiGbJPFO74ozm
r4TArnobKWYM91Y3CtKuV+xwhzdMW1EmCWtA/wj2exCW4MtcHgGKtttldYuasVt/
JG88g9kdgbn7QGutzkOsydD6pTH87KBxeKShBVG7Yq+WsajDcEFY3Vg09H1w9N1g
pfSYEYBz37khdMZ9OrTrP7NIXIDoOVWJFO+QRhJSvyC6krCpOqOu6k7LBA3dKzjP
rb+cq51pZGmhnmXUaopkyXMkzUXx3uMAd3U44xCoi+76D1x/F5xNl+HPK1T+KmNY
6LdftnxQnJVUFHsWkxc6pDgmFwCFK20r+5/jLWHZlBinNl8KqU32o1usE9codi4w
74QMkww5OWWu90F/UM5kvtXHl4XJzSZ74nZN8Apa7f2ocVQeGSHnV5SFYryPx1dr
NsKbog1TtLTKt7wr587UH7q6+4Kh6btDOVfMoR0rui56xUA3q9VcylS5vwG3qwKa
24sxJLELHMeMTCousv3chCABp60M+YaTe714KMFQp6HRae5ynPKLz32WjPYTfteC
9BuskVurynhCUKLib0bUUY6Mv4dBxxrdb+T4ju55t04GQLxMsLecJKAKKYFlzlDs
+d5JEloqxmLhXMUN99AD3YvIpxSyALbhNUU7aYWScM1No0WzQtVAhioLOxARkk7i
tXgUpMlwmOqhMC0QYGRjm2yIIWhKCN3Den0Ws7/Mqfh4x+B7DssPQThEwie0wia5
iYJRow6T/AUgnH/pi9sKeC6S4orSG90KPj//HMbF6fRQjdfboElWffnVXlJKNW7Z
L+Wbz88KOvS72DmfiQPEN0ef77Oo4q8qOtTwZ/8njeoadijwCOmga+4Gin4/KWbV
5Gyd71r5nbvv7Uq0M1k6csWLvpUy6vlPl8D15OyWdEXNhVe/go4zkrnNdIupODvn
nxlgiD/dN17RIBWP75ADq2/9mX7ENh/ILZcD3KsHKtcfujRGrEcYrrOWbFSJHbFF
SLwM4AK7sw+zEkA0K+MFg767/3+NYsGEtFjQpQ4quEDYLOW4zBs36rSI2Wi7Nyto
XRSkXUFIb75WJ5oE0NZ0i97PRv5+33IqSsLmjOrQCZZDNHy6bxzQ4K9RG0CEm8H6
rSV0BowiHJXD5KSlOckM1GgBkKjAo68Pyvgk/7cC1NYFYqd7fHOzqcdf/1xA927F
gwn8DW9hv73/Lb18rl3lUnKWyTyU3rZTMiRj3H4UoapWfxc4svx1j6tbYuH/GWTe
8a2pc2A6JlAYptYm9lgeu7OaVUfiuK8K23fmEUvdj8dPTogCv0mpfVdhJxsbPVL2
WZpMuHeW0irjRdFRrHQrllkVq1mw0g0Nz5Djc8Gi1G9nnuO3kDTv4gDwbZd6Tm3J
lEkh7ecVBE4eWq3xKulWiVPKGE6pZZVxxnP0PE+SUba1M1vQhots2LefZ98sFNI+
LUn8g/R0Nq+7nzd+t+Xb0POwIgb1rmU7LAFGvRMjEJBnF2uasz6X+2nZHxK7uXY7
dTafOLkUNsjyZwpZik5ELYMQ+bWWhp4ibwJXkg5VcUMsIITnE2MZIVFMud3tZdZL
+N9caP2WLH0+bDotBhZq+sGzgNZr1Zwj1d64lGYG2zHDBoJZ5Aq2Hl84f0ETbiZ2
MVmvuDWj6Q6DiJDDfGZGL3mpmYfPrMQqxKswKOLQiGUc6saIA9GcU/rUdp0HR6W+
MF/pfVFtgK0RkmyOJt4FA/R7ixRQlwmBNQkgotk/qatk0erbXFH+Mv305K/0G41i
B0/ZkmYdNYsNixBahEP5qoLlr39WSIoed+pHuuyNmiXYFYcLnG2+0uISwQkH+eyt
18sdbm22eV2VVUdXPOmvNG/QQv/K/Jy8NnjoF+FV3zMJsbI97sm6Sgqw4/I11RZ+
Bq7tcYFSluSKMWics/2Yv7P+BIqjngfxsm5MbZHKtIGoU5Nv83R2wGK4mVkHFJI0
seD9LSiCibYJMJi8BswUK7DVxm8zxOWlWJBd9bossVx8gmUwv1puv0BZAUQBsGFT
mXsMMfQaKJOfOujsnunt2WCJv5tMHNbd4aMsl1FA2olxOECL2Hv8sisG9iGiJeO7
rfNTMZPKbUuY3zkydn2bHxfKjZE2ZcBjLQxKUPTPQACVo12l//1XJnMztV9K7ofA
0QJDkHwba8RQhBG8T3lJ3dGmXyo47o87gXnDV50Z7oQGIwQVNUeUYVbw3FnPxbrJ
8s7V7xGMW4W3VNz1SFC+l6DtAwm/38IeIXnrGY0jInWB4Qm8oRff1icwHa01z6vo
E98UqNmQHVhBQ1vxAqlhHrecOb8Oy81tWUHGEvXm7cS/nodB0Z/MkJraWEUN0mI3
+mYwF92Uu8aCCRtnZXj7yEOmtBcYLmG+34l+vrBNmjytgJQEO8xU3sscgW2jyS/7
3fzci2H8J2PDZwtv5PAUgSZNZKrfnOxMf+rIP5G/YuTm9cWHcgz2m0Rq4SKR+C+G
CH3hw+7+gKDez2r0Q4KkOaQZFs0ElU8koO6YXi/nLvyN5E55E/WEQzkUas9GtPHh
nE6xufqTA/tv0MmTmtFaCFj8FAYGshXqpJnZzYacSU6dHStaYPVv249lNG5VOBun
L80lDgh9Xln88sX4R+pbiPzRExetIbAGBW41mXu0tKn58dxnjcJe5Vtu+qmDuEyK
x7dZM0W+LO0RTZjiAECYhkZuutJVHG5s/CPEmwIlg8aqUl3a/Q4GDH6gd4EJ0R21
BqfVD2icuXbfJoyJv8tWy4kDkSHe3tZ47/N4TRTHRHAEwqIz72Lejax/2auCSgT9
MEa+63GERUMw8MYAqdtIio/rsSGzwULNoglyXMgHJksiAhVDonsaWBNPLjW2800L
2nNtEfEGgMFwowIuhUOMKUPLU7MFcf90jfh19tP+lbJKZW0Zra+ceLElmFsSBNSG
UDA0TABHz4WeXWYvrPIFHZW5n8ZnD8DmuoKllUWGX+ij+9B5ThY+hhiBsS852gtu
mhTN673c59a6nbkvmzULXR0s2MCgue61YJquieZqbli45dhllLUFB1Iz52R9c/Bj
LBJiwRwjd+XbUiCy3evehiZj4GlvQkO/nbL4OUmp25HvNChJZQk9WufiB9yLIpK6
IGmOMY3RYK/w3rizym9+LVr6yqZYJb8BXF79LLjsrnm7G4huRCyRxex7QiRLy1PZ
5Pqy5CCWbHuCVqAylJUKxI7gpgw0YWXJgCSeZxASHXOpQg3C6tCjHborc5LMY5tp
5iWuXCkI2bbOUVwtqxhxWwe345jmZKmieUJPr3qy31D6G1A9c+05qWDklvB+5D+V
MZEd+zSMsyDfOJyLJNNKNMR/KJaRMjSLFFIjLKDTqsVSutfKSVqKQTlw63lfcS9r
vgSp0d8+rQ82in6mXv9Gb66X+SgpPsdH7VQ7GwsWbCgugUxqSzkONDt1ec8Rqvx2
zzXb/GFltVIYMb/SH9Mh+FIzP2Fal4LSy6zqSfodPKiwV9Cy9Vp6K12wniYgDfgQ
ZcS++UpeQzLH7l+zi1txirZA1+mCw2ROS73GjrvOh3QXJXpCC0E12KI7rCHDdj3i
95TeFAbEbnnCzH2reyffwgjKF/iCcB+s+1QqZGAib8+5iWUHdnzcLXRZ8iXoBpsd
A8crIxy/mkQcVZAid7wJVAF0k78LqTDOj9NnayUdrUeIyR0XNyMsXS1DjGW3Yriw
/lSVvR44KMAe47paeHG1Fq6bUUpSblSq3OGiaFensZUbdwhuJtx2NnEXA5Dp0J3G
SyhPjX1pP5Q0ey+nrTTJHN4gHsAEP/7q73tL2VEgSYbCrxibuWy1+V5sxGnz8rE2
zcgWQFigWoZA9Tvkk2pbT1tilJK3FH6Vhb5wKng/R8VDFKvlQL/KQhJJcDx8J0tS
60mdNCMmHFjw5RrBA/Huo3hkEzvLvoaffGpFd7GraBA+msYa7OmwGLEAz1xtQUJO
VaqXkWR6zljREWAM1Cz2J9z/jzmDhs3axarH6xlOVzqvT4h9fiUCiURsdoQxqKqN
My3jrzkGZlzA93eQGAED8dOfGzrT3OEigQb73hAkIX1Amq3xsOD1tI6YrvHSejDs
zkDVTX8ZKNlK2NYY8Kt8/bgZgygv8X1AOTUlUKQUfErPv4sXk2lbHvmtqBkxQ8r4
gwDOw5Ns7/hR9b5VJuuSkdOCQJzlMyLYG2pJeJxwOeMFLxw1pudZa9rzbPgxkty7
ecV4ef9ttG28w+mPu5pYZ2lj/sYUA/l02uKImBUY8vF65S+ds/KjAE1QIVpRoFXO
hqxM5qDG5D3Gz5guI0WFmt5ZbQiCTJJ3kC+TjmHmMk5NbMi3Lv/lQ+0FHBjEArZ+
4I6KjfL/xxGHFYmhhKj/C4IoSZWNJiyXpxeYn6Fu+lZ4ZVDQeWvrpRLsxnybxqx4
qByDG9Hi1Yc0Z2PzMVkmGr8hgPg0+ihYoCGTz9fIJRvq1UE2BZj/nIXDg1sR1WGU
8zL1Setxtn3Jnk5A24UsjJt5Q+w++nSUBDeyGU4ega0tnY1fG7BNBPifn1wRVMM3
JYlc7YuW2mVfq0J2cXzMj6rVZEFpegyZhLASpLgFFcgA0Ag44sBACq0p2VkeaMg5
ohnky3XPvnaVuPxPAjHxYnlHVFDhANUn7chrnf2f0mB8T3oONQiu5VPZBW+2A2Fw
QGCAY3nk2qdex7Y59dyHijIbXJ6jp+iCJGj+5HkkRXRKVmC0DzcjkxV/I2sjp72S
E06N0I8wXE2YdmJ0DJjss0ZR5KSOIlbsQGUUz/krXvKpoNB9iuWhXa83M7Eqo7em
nmqgk9AvChq4dcgqQKxalTiozsXulJYULiItf1cx19hgH5FeBkqP0cmvwKzEHKlj
4/1c8dlDGaSv9ykDdlQRzdhyiTj3+GmM4n7a3c5mM31+mVWHWC5FNY2jbhxNn9Lw
HVDyVIi/Z4zMqlOzKy+YY0KyjggRBS337jkX8NFORNSuT4IaykcMBHuox2Fjqg+g
M6m+x6MsxKTmLz7HG6sGWfIY7KNu8cGgR8cCcJJed+lEA/gHQcO/8GvGO7ot9ob5
lt4gNxKp8gaxxcOtk7nFLQ0Y78Ztzu9BZDfq4p1ye0dzO2Xlh7D2HlyQL4tFmxwx
Q/PwrpXZR0eIOc+uQJu6CRBpuWtPz8038H0nfq3wuHE1oe8ktrlYAWXws59IPwrK
xUg9voOMCcGj+WHkMGlmMuxjJUwBAwzw6ia0xsBIP6kHgBf4KZ3slQJp5Qj++e0J
FWC2beDonvdJozYky4xgCEMtXG7HtbVrP3pCwu8jPDIq54970b9a77k+CBIaqijC
3ib3zbYuSZG7YckbWbN4bo/IEx3UbnMJxtyPyLbHOy1GWphYhRe0t7iRMw7ywhsT
5t955MageGmIhZeqbcVH9tQGVCnnDyP2Fq2daXIYsW2KqenUFH+wvlyiyKxk036m
4qS94NLGSz8hnU9PGiFmG5qXT+wxbbLYA003NoWC5ikFR+L9MLuGFbTq7YnoCvRr
7glnuIJDA3jZUb84cgiGbxJCBayYaAW3tet0j6FJonEWo9ik63yViobd4jlCVmAR
N309bTVfLl5eKlycJqJkuzM9OoHbKrjAShLfw8k4iPPy3RlAgNAmaMDulN+evAlh
IoNfalcgfeBhYrmx+ZIQzJA3fJX6wMzBIU67nk3f2VkXJ6D+JwAVS8fpxmT6sKQN
VSOta02W8xlun3x47/Ah9rW/30YAzt7CunFTIJsK8BNF+tFPE/PvfSM4kVMg5kX4
yHo1grp56nX+pn46aqdJ5+9kI6y7XV0E6xtiwufmq8jOjM7O+IvFVIygj/lB3JUA
h9J+06lvc7PoWouWgO8DMOI9hRfX8mrgePy7CFZqdqH0rzb1DYnwxODQWtUfCrJe
JsjBUejxWmRWz7WMukmkFNBvbrd+uWWsfXrzNnUkf09gGyA4Ysr0JbAeJ6+lbLnz
YFrmMpV5xR248WTYl2LDUgs8ywj2hqekODyKjYgbBI3+rMhjEbF4fFBbmGhPqye7
uKxE+UG4j7qSY+Ke51uGJvGIfRSoosWXvBsdVuFuwg8oc7qRHPMEwpiqudpgu/bV
EdgjeFErb5O/wGJWj/vRhflyxo0noZp+TNt8kZoJr6wNnnSxR/NvAvd/hOsU8Tu3
4sGorIEegFMMVKF9fd86amyBRl3q4SfrZLs+72jy1zml4/jU+2pXU/hwUtLvQVTr
hd/QLgm/qGVzbSb1irEVSt7T2JVDPV/lRb8q+JZZx5USRDQO2g2DhIu1oNiv/GZh
GIx3VQLG88Shsm36JrQ/mnfwuChhyvs7+aixOW/AJCvMhGCRzq41PoUxtSYyG1UL
kLrH5XK+gCWW+mhvP7pXiPwNHEa7jzGLxVu4oS3z3/symG59WLgRO3+r4kyw4W3F
2Dbm5LdCo5uZFJ0Sir9LwY2kFSeynb7wnUgUvyKZ9e89VbgGV1evRLhGoyjiD1Gf
GtRhaH1rA9LYUNtBFEKRV5fvper11HUgeK0TNcuZycwyo0vY4EtGYMMQPM/UtRqq
nQFrxejgwp3rSgIpMgOuJ2mvfGQ9bWP5rMGRRLsE3Lw2rB5lxXpyYFixmOq6Fns0
JKg1o9xN4lvqSYBwxbWI2LohvSuwqD1ShJ4WnDzRQKPSZtlyiCt4w6w+i3iyVM5B
ea6Dx0n2deK4OPXWs8eL4cXl7V6ot0egqHA2C+UNJRjenrX6AEsTg3QJElQSs5V4
IQGvyPT1Dfy60969ggGb16EYjv6NctHS/jhdO5VVSu/zCI80MLPaK3dWezlMne+o
fpSkDYU7HcsapWGGFDwx/pte43vKPVIuw9sKe2dHir3gFmMnlDInP3WYlmJS1AD0
p8dyHkDgbbVTtQ4p3JKuvf0dMYVSHy7pzbfRO+zgK0my8KXawdJxe4NocaT2pHtZ
RehWjKoztkJhY+ZENJPdyRujv3bcjEPcGmvcIN7TpdSGtb7T3Z34ehBnPMyovry+
kfhlDBV8JpwjM/Om/8I/2bOJlgI75ntTqt/i2VqiIUIVghvIelN28K4zATs5famK
Y2Fo/e9JR4aGGJaW0F3/WTKpOyL58jAQIK0Wk/MBDHDWf/b8awCgIxUh8IT657NC
e4qj6UAxm924cQuOeCisLtFDstyMPpozZG1enAJAQ89CyMjc1QHSr1ElgpyBby5J
vgLQ3vDVXHrh6dSw7o1M0Kdl9Ccz97qgx9DdiUO/3YMju5fTuzfS7357jRUCnA20
XQh0dbscDUp92gMe8rx0g/JhXHeU3SNOJmDrO7dWiUJyQmsJFZp6PEe3HuBl/tCK
zhVmjjDUI1u5Svlsfk3l1B+O8TJC90STT15XuKEnDSKwNE2RpJ/hYodfV6va1mj7
ieP53zJutl60PtcFPOcmYXe0YCJil9ldTI4IkT444ub9n8F2aeuLjtr0C57yLPAu
fPTp6Dub6VM1RVff68WBcFIKXUVAp3Vfdfw1r38d3U2NDC9tAoXfcR6XDPDf3Fha
gB9Pwh9kgCamua4GY2zIJmmA7CrI72hvZnu7l/WNQPrwyqFJT116BDOmhlqXGkc3
IR8yUxf+xYLlbgndJ+1PawHp7eULEKujIepjuCsr8KbgvRNmBY3id8wI6ps278T/
qTWyYcE/tJGto30yij7kkOXh1udvPWPqP9KPKB0EBgJ2RigcRcstBON2VFcclSaJ
ZEOgcebSWQE7SSAQvuXy5YoPs/Bbw/Y1atHtV6UMw74G2rXLOQbI+E4E1Ic2k6E0
5YRH6UoCyLCB9QDKzzhDEtn0MeuY/hCYu8x2QMnCYtSt2vJGMMpTSfEbc2LArBPX
seD5FIdQaWBOyzcBWF3tb6h0q7yp+0yo7nx9A9vTQvOLUkWO6DFuqnm2T3glMBQY
VwRrA6u/5TT48jkMaBcvjOEr8Zi58nLUBAg8si3fiUFEzGj6YtzRh2MpdnisyuZt
FFe7+ak3Vbv43dVPeUG/ZhtoTbwiOaNHwITKPzWiDRiZ3qc74AmdzM2YkK/hpdh4
Yl2/9MMfyOdHBocSdpJnZBbmOd+QnaYQLlbCBK5WLyPWd1YyO1jxPobOCC+j9hrL
3yHPOGuDLRUqwygPfFxzJ5mJlQvtaiDXl+tACRPzcOIox3HMoiU6sHdHOQdCi767
fAUPLm+V5LK42arZr/UXhV+SV/r2wAkst6PK3yPtZw9VfrpN6yxmEAIznF+wocPL
FjgSHSKf5jtbQMJgyG+a18rzDS6JkKzCAW3vGHBRED+Q9hDRhNLaOHAMtqAx9FwO
WXUCqFYhqf90VkQnTmncc6/K0aay7BgQXpYJZhnDxu+MUsIkKd8oMPfKyk0R+3xs
R9IB5P9jtr1M4bs+b8hei9zSEnGd9IG4JXY/hUC7fyirjh7gL1cbq0lE22nzCyM2
4oyNh0K13KP+OvlnPmGuZDByNhWrp5YX6E4P+zYu+4dPhi+xWIVAdb18px5lBcVR
xNbtniQx6YQzqcp2UEQI9hFGUPJQ+lPLcNL3JSS4uuhfX17vj0IYPaIR7PgePlpa
/8qF/n+Po0Z0l7tm8LC4hQyWDZZX0U2iww0pp6CbiSW6odYKbYOpjzQoyzijwe6u
QV7B4nm6Qp93c2FkpM/teTjEKy1VdI+0LjXWu1qA+0M4EeNynlPKpHdo8BiIygN9
wulX/agll9Fts2jpYtRNP9x+3qLYZkDUGOoX0PjXb7YYE/czYqmUWZTqPs8JV0Bn
IDzNAMxW0ngvudMAra6h3OcOa2lhfXxJSG2tMi8zbmouHKS7Wr5mYMnQPpt8cU/w
tasmTFYUuhscqo0HMigXmHyt2o7cy6g0h10naFaleUHoHf+3OQ4iskE7IIM0pui1
HIJDchGdXytfW8cRXBLuZAKlWizTPFzKt7GOds1kLNtylwrqg8ftMGxPAuupF4qs
wKCsXmZVH4KzHpRu5VgKffIbkXnd4xGm6AHJ55Mw/OwzHN6m4JQdXPOIKboH+lR+
Lun5hkeNfFEbShc5sJ2qvapZR4BVNuWM2CgkZKPezIqC4sLh7rvgnBXYwYUXtJ1h
b6k0wf04y+Ul4awGSHj6YnUeD6mJfpm4gXV0eJnh28XqBwPGmJgPT0w41NOIP/mB
um08ir2vfA8j7kau5dx6e6Td8wXBBxYYM+AeldPUCbXA80G6kVqmrR8yLVlVYZ0z
t3kD2Vst9ov5g1KI0Qr094pXqeOCR9yxT0R95cfQeXJzkLkWLyDOy/rxdgk4otMc
PIcDvvRMLx8Fg89nrGKWMMKyL4hPEt1sj1CI1zB88c7Sau7T9Sk/gZdShhtPXxLm
fOU9r1kc8D7tgd9OVPmwBL9CwkZ1UfmTLuxTOcWrRi8bwq9MCC0feeCDNf7oQzH/
0HxrzdRHwV4qxAU/t1LwIjBIshz440zfePxFQrhowbGnlqE0T0x8qfTSjocK5vk4
MTkCaZPg02jXny7eAZFZw0KJKWCTgivh5zsI+wtmYkUgvn9UNlD/pgtUkK+CiMPa
do/A3QB8GYltM7h7jPmKJq6dqgis5JanWj9ouYEvH/XoPBsYhdb17Y32IePifM84
dw/ZTjuCZVGXHL5YQaBAMBSiq4wuc/YU6QKuEGVKil9mWhrcs4xij+O1Z+TPVez1
tuApqW5H+OxITIOgG4YpnoQKeTj/j+fBfaE9R26/SLR6oQ0nH8r5RW/OcE/iNNKI
nq41fP1xvar5XcL6ZvJcqYCP648nhZ9G9T6mRXGtRND/66pfYI7UISmOWlfiFZTc
PRhbkT2q4APBnW0ZeOpFF2zqxWKyL8888bzLgxRi2LHplpnblGp+Hbg93HREOBNL
eu/dutw3pFlFmvyMFkS+ytLQXJZG/Mjxypcr+TdfJeXCFg2i10pKQqDctYKIP8Ey
rBDOrBlPELLnW9QAanhyCOzZGuEIf+uCTgWZXwd9ShiQsR8pOMwkVbWaRnA9oFj2
AqO6Ey0vO/+uqUWsvp08Ih9UufJWqGubZd/kpFQB2Cg5Fb9zszIJBY0WkwCklYTr
1/qtwRlnRbENgtznjMeY+hjOQr0eQGWgEck9lP6Jc7vOwgGfcH6FoGzeYN7Xf1da
OGN7XTkRPQmV1l/Nq65tvqOmk5R67FAlzh02iSy/lgjsBh83mj7aa45piIqxZRlb
YfuG4TbdHekgrJocC6dz+Tq2GTAYrh0VzJjRSyVCvXQpcAtnCqPG+QRxXu8Nbh6q
wGEXIRAujz8Gkt4th5Pkzw1n2dNd6g+F6HzLVAO7cxWBkFKLGdMDg88HmS4NZju0
oFwlNR3mZbn0XcMjyPXlzSEvLCufoGQqEXKQ5jLJ1uEDcoF55SkysFpk0zis+uCw
PbCaLn7pylm2qNym0pFcLpCbwebs13anG3PruP5+AhpVTcPXA7FLk1WfASHt3sRr
3uPic3EFbNPjvO9AQtjXSVJqnOssJOWfwAv0VwH0d6OShFJsMOvdEaaluBnF0dTv
HoE9iPWWp0mSynd6qtnbVtZzydI9beRbECgyZgYb8bhnkU6sJXPXw3SJWPN7FEMj
m3qQNtFpbJDO6Be/sgsXF/h5D2dmaYVLjr/y/9BaGL1HjPiEC85qbqR6jN6KtMCt
gVaPngK6/SL+Yqi0ZXv5/DmEdo2vRGv6yHq9E+UpiRoqTrAkLQSeC2uDoFzPZARX
XdICOkP1WJXAmGjsO8jomL9BQwojATvF69l6YqzCGV0N1P9HbUkb90lumL7KT2iF
cz7HdmMGMTYn3bVx9JTfDEEV30HFcNHXlphySAIj+QBNZqUSydAEwI7ltSuZ7W6I
xOBsLlpQuQU8SpKLPNDcZsVhygsLxZ3XuwpMxaqWUxuVi7DQnLj5mbaMyVwLuouw
GSIzc0UBftz0NDCXBEfeU0Sb+x+4pzEdN4S0QycDSoXFyK0zz+2YS1W2wG7y6wKl
BUueWkOW4sNzPWsW1Vxo089TjjH/fIEM9V8w0VsvmzjFOfkKFJgp3a5DWw3GwjoT
xMbFufysLYOX2e2hYx/jJS70KrkNgE5ACJoNhJfNYClC6GzvBBhLQ+AEwFJZ9K68
lCvh92gLac0EAyi1HyE9ZM2hCbWgfr4/FKVhanKbo1yhYbVz97q5dzgMDp1oTqje
m96fP147Bd/eoa6r4XwgbaREPjETGDK36KAdJugAKHrXTQs8327m1MfdisIgfyxr
LJkL7vvQnJ8sXjVS1dWeBJpkQmNlZAxMGdMrXxWDkeYeVlLwcB2hBKD7KHATrkZA
8m5GnMjct2ObuMIuNoF2hCPcmGdxTXHls+CGO9rq74KCfDw2t1PRUm4wY+APSLkt
hSiiAwXsHdbvdwdTKtOIveDYZOAvrUnwe6g5rPuRs5WItJsE8KB1riP33OAgS1uH
AUiLto+3s0Q+I4EiNiWQ9eKOFF9S5u+bVK5mBlCXDToFqU2UvlbBqhsbkTaY5eGC
DyOmEkxmEkWIaETtT7ahHSuvlJKGkhLrAYiwVXyBWES/KXYJRwzDFLReyMzM8LoI
vmbRZC1flGxgmAG8B1RUqW7m/+7WwMciDuBLzF1dnMP5VAZ5y3VFBXLciLvO7S6e
bTDtuWxJfunEJETDbPrz+BE3WaBROYBXXIOh79L1CPO9Vg+kYoknFlzWaRB49Hn0
h2VtfdeY9RUMAneXvALuGpq0Ma0dsz/YkLysMTxJzK0noNvibSfGz6huAcCUCPK5
UFb4lQX+iaGBtELtR2FZpidTgNjLeVqpDA5iICUqOIrIswQ9Ti/w45IhjnefBYc4
YR3LW36h6mQgEhaNz5hdWu7vHrsn4j6lOmqsXP5pkMmXZhtJpjvvue3cyy1AGbxF
hgrt3DAEPfxswy8XdW/Kw72IaRJQAjJ619ATcvf2HENaQ76C8O4o9vfnAcek+0/2
49G1sQiqeMBHMI/iD4eV+Qcpp6Gi6BRpYLLFq0Mcm6j+wnwOV0JdKTU03iApGbeX
+99ceSwtLBm7jsQUqcwrFScu4uoqcYrBnmvOmVbHk5Esl2KwPIm5hY+ilHH263pp
asNettfuoq1seNbmLa8EwhIZ4Bg8zw4DQR5+q0fWyYTMnjZpUg8gHhZDDg9hO0M0
5zcP6540tW8CwLZYTlGlsA/4isoMxjrcUepMECJRVosSUjgrvsnn/Y4iAbYRCg6B
nQkckt0wBXbeogBdKJVs7XOLx1uM2CSl+hAwH81IFYezFzKIi4WxTcM9ytuOvR+5
aZ8qCGNoe2a0cB9DPVntwNbwzjXS4o5PvPsglWu/1VLXKQApjDVwGUgOKY5zmQgk
1T7codw+UDvEwef8F9rVwVKDGyQSf7TDem39BibJD80ImTYkeJBKvFAWiXFUWCPW
X6Da2H/8xhSUEB+gCzMZJ1et98wnHPEbg8jnKMNf4KH+NP00OPdPKAMKZ8vm/0SU
eA1uGtU4J6dhtKUuYilSqsdt6D+Jdj2bNGCmgFYrH7zD91t0mIEYPuujfpRoV9xR
JIZnnsVgxJndMlrLI4ZHzXcWUQWKuVnxBE8O6zVcWfh4LF0fNMYxBLf9ehGjqqLj
PjZJcuC9Z64gXuLsu4fezqM+RoDyqOs0dKh0TQG/gS6FGkdy4Sba0E1XxR5oedbG
yDJjK3W8wKrKRg8EuGwco6rnTx2rt5EkxoLoDapxMRfJrdr60EyuYvzuD4qDkNn5
i/ogS/NJYUmlVfmkAyfRU5Nuwob8E+PGI3wFnwecvDBd5iCWtL9AZJ79J5MmIHkC
9/4WWEwgdycxo4FRIsw61XjFd6ATb7qX1QbvYvpSMFYx3EpI9tyBaDn8//GBVvH3
LebIvJRImHQkrYpSpP0+Fr+1Vh3/4k1YgEOd16Dtbb9n73+9oCrJuLEFIAdsq3GV
Q/ZzK084CKNbKV3iiUKwF7DwQp7au2GLE/1NdlmPYt/8rbKHLB7WCkAofOsMkhzi
2RPNszQSmyVaDLuJCLKx8K2xn4K4qjCuilyHqpVZELQQYaILXlcseOvkGLkl/PRJ
XppmnEovWP5Aj0grYfCtLW1tYemY+ybig6Vis1n8isKEqDSxpUI8ZSAP7Psyyk/M
JvGDq/T0iTB+orPYGUv+SVJM1p85pkT2FJGnm6OGjCMKfOqS1EX9+ofbHrpGYmIV
FsAq3Evl6bXczAyv7V1DchHxjbptYlEIyJrUJ97t81tTfO0LWYxMvOAT3hbGuin0
5+Nnda7KhaF7l4bG3QnAfhSIifcUXVfJNWN04x52pEqeTyaIjz0ulpm2IvFALQPw
j7Hb7alr0Sye9ECOhUNK03XmCtU7/rf1Hxfek8cyLvBhD0HzkdVgU8+06VZAQiQw
VPIt3JHZp9g1Bsk/aHVLniZ5I32dGcE1B7Tf1m2rkC+YIIbRgNXygiiZkb5iAhhY
dyuM788HxOHWLSoD4NbKqgs9K9xCOsdjvHmh53z+6MrmwgS1zT6edILzipK1GSGy
un3trOPoUu+/Gt/14xUW4xsIr71uIoLGzOFxJG2S80gteIFXm/dZROpRT2a1XG5b
/0csSAmlLszk/pO0RqyMl+MSvml7MwYQDCncK/QpB0B90lq98CYoxZnyXkUX928A
2bEjFkryQ70ag4Wg0Keb+Fgo7WchrMe9LVVwcWIMkZJKkCGcX3/fK8t9UWpgKEad
3nGgEdJrvFH90YHe4YiZy6E/WajTwtTN1/3+l0rcZ8r302zEJmI/q4NFOqtuQ5f1
8a0ALOX/K41EC75JiC8Pn5TYwzwZAbEz3Llm+AZm1GYoZ2fq138UhFiOm5Zr3xyb
NcZFvsOkJ+SKFWJdjCxqkgGq+pDpaCmTDYIUcPjagaXX2v74GVrdVJGFDdj0vLtt
eUTkk3mjlKYyv2btdNs3wBJwRzqMmu6ec2ds1lNZR7ZIPdWYt9kWQDmas5fa6ALo
0kw/tVTLMsBF2Puwbhu+PjpuQoqiSPXKjuvhMFA2Zsx5/6pgGli67UkpYuf2xRli
eZaxOYPWUNjL9fkrWdRTsuIX3em6oViLXxjrtBxrQRouSqDqKSYNJsEBh1Y0m4Ia
QuL8AddhyXFDjQl4UIvdrUIVKVcmj3kTsfRFH8Xo2PUAyztSxaFTe4pgypYdKmBC
IWyQ/LQoEvFgrIfF3hFb4sC7JUN4E+nNUIdwVs33StcMbsEPPyrrET+hGaa/7PWL
Xars5dn6KNExsSN7np2y0aTVjnq8eP9iU8NfEBlPd/ab8hoNGVUepU7QJq2pl5u6
kI5NtK5zGbRpQ0fq5+cMTXSE2kVCb+PI+Hs3Q7v9NVpx7069F0J98r8Kyy1tkc+x
rbnnyxi37j4ySrdHI7LgVeMJcCt4meFqpTRH2lhUjd2LeG48DswyEwfq3rncanVA
TjSQNPGgra5gyZK/QhGJXmQMrpeTc7y+a/4L8fEk2TenZ2pbubv0fohxQ79rnH59
w9o3rYZKgZ6tUZf/WZQY3JV2ZsTZYpxr5QNZZeZapoKBOB5YSsqHPReofJlR0Heo
Ki+o3HqxgIWgZjsim7iz7D63bbPQy5b9sL/02gzFi04Xpsb+s1lZpca2mSxHkmRY
kTQY1phj0wZ5OLci0HrsMOXVDjhZ1vx1m1d7y1AoKwTYlucPABT+H+HRDLFN//Cl
ewv2Kr+dOY9htAkkA+c07tpxPxaRPLe+nVKjpphsx/qGGCPx5CoKUzZLbNFcUypv
96RIKNvKiW9vmSY+4onEj689mNS0Ee79E6ekYAXHHi39HMEw6kGl3vYP4jJ2ZDI5
TVpJVAgfmHrlaCItkJhxzq/B++tLL/PKW5eV3MeO7shUUaUsc3JDYj197QGWVz04
E/56bTHU/C6RsxboExwlf8CXzVxxJrqaKDlWk/6zInfcGnS28WJ9VatO6QVjGGsk
DTRWLyW2LjbsKcbCuJu/V9QZm4FM8D6LLQ8co/0CdalFwW55TfpSL8afxX9w3Bfk
STBqv1CEG0ScO19bXLqbGk1Gtb+NRtZDSXXPNsGHXpdDgYRLrgkFF1vADXPIaqK2
mUs3mZsAwuHv2zhT0GjdNru1rw0Vy2DVf/H17FzJqSqfuAjbZSoKMeCAbJmSOETC
HbEcOjrVzbKXGjsZ1E65wc9ONWHxF1jGsT4eQg3bd+FE7zJwdX0ByaRpdaw6gSsA
xtjovxzIJYGPpyU0ovetBkuOoifgXAOuc/yc6h3hz5KI/FfBgb9DFqXEpIr/b7qZ
9gOH3DxJtJr9roEbj65j8ZbOfO+GJBb+1v/MxPPKx3uBb9yJ6XIZpp8E3RcUA18S
Qmc7PflkWuppIzUeOe2jMqP1T70202NgD30oSMkKZxeMd2IexBEGQxBkR+4XdIKe
RW5l5uanjWGxxjhxeruFIuYgoAAIpa9vqEiJCBmzeAZ8k+WfE5oU/q5Yo6ZbPoxa
aEvGocfnCQKr7YKo9URZjeCfoCoICwVxQAp791Ef7iI=
`protect END_PROTECTED
