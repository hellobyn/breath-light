`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqQKjYi1uoPYWSwh1m67+Ib8NxqK5lXbGHurhdTavkFUswAN5xxIlcar9ota30ar
5A0cXPQdzHAuzZB5hx7EMPeMInUQCbyw8BCcaqmLx8W0JOAxPQn2rDblc2PMa9h+
0esQddDWGnjI98BRG5QD4+4wWj0ootZTzsYNGer/PPrhfSzXRBiquvlhLmIcQIHb
icw99zh9rWHSwJ1N9rbFK8IqDCM61lkGpAu00/GaOdsAkc33/kTObFq63vz8o3rY
BTdWD+BILUhw+8UJKJlofHki0+CXN29M46THZJhWFcLphuwWoPg4JJbc+p2BQ9w7
zYbPMwnmU/ADwyJi56Yt6jSGUDMduwuNfyQYAPqZ6Ll62tRPB/g2U9thtdgqD/MU
5BdpPs9+7L4ZvsHVB5LeNbuYjiWZxENK3Is4vBNESGrHQ4x4/bYCBoW4PwQwjxHW
7uhO8UH47emJiinlrr5+g6KyhtPcDYXtPKeRNEgkwIj+XtCKEUa5FUeo+pc1v7zm
wKHi5mcBVvuPmmSPPIzmrFYmmOr8gELj+dbqZYZ3LSvxNCFPIuxhcfrgBkjCj8wl
3Nf6VtJDv5cdE7slAJQKZZvGtit388zZ5bQL2OhPk9TMbjLLXJ9Z90qgW3XXYzxT
t2HIfA/YfZ0oCXnAPf/XzG8uCYqVdI6Ja9ajCM2MU0qf8dbjN1cbU4cmtfnVh8J8
IaGpfEnk7FNwl6+ch84P8w/nmngdta5sach42ryDjmj8FlDX+4mtifBfp6mSv8KU
DLgBX020KVt31CBBgIExvWdO5LPJtvtdsMejGov7/mUvhRrvyoa5nRKJjoFHCIqJ
ipdG5/uzNkzAtCOhW5DrhjopR8qyDi2P2vjM/snJAFwNYbKHp5TFVeuJ81XIq+VI
LuBzFSWoCN+Tq3G5rFuU37KTv3EUUrXzxk7/hh7noTDsXD/fjtUZODqa7V2Cco5g
tt2H63ajY4DklxHeFupwG1gkGP/LroIATtLwMnmsEU7hwl5exXVQN20K+2P25G1n
tVWIXdMQxeagJh4F0eDMUxTNGnsu3oyzvoLZwMG36xuMpCe6yWxKaP3TT6H1LJaY
0HQS8ym5DrkQWEf3+Ij2LLL26nDpTvMy9ZIBa4cMhzHNXRiK6+DBH1iB4V9my5FI
y6ocrskh8qLg/OiCAOrRV7uZ3U8Vff8IjroOHFoAcw2I6GgGoVw66hNVT8mtNsvg
2y/1x+y+wj0taWxq3vGrFlOSizdWuTjgr2iJ8ym8I5tFr+QuKsMC7WUHNAdV45AC
UF+QMTTFh7hUjcdpSnFt4tEzaA//KUgGWbKcM9QJpsigVKfYj3U3sKozcUYracl6
YgfMhMEaiOqW+EVVkEVzKnspU9xNBNWnZC2pAKsiuYNS8GTz3fo5aB6BRMsVT8hf
YNCKXkxaMMGV9q59WOUDJzqrJHuJxawTfECox5zpZLkObW74HWBIsUodD1NmQI8A
8fCQMVVoEpl82KYVEhuUOW3+gqCvcNAL00Rc8uKMfw8nmf/g46cX1U0emosrFx7h
X01nfGvyQ34+A1Ja2+ZZjsFwnwNKw0cSLYzMGzJpHhDAsrkO2d861ptzNlbXeGMI
qc9hj31bow+yJ6TNPEBtjM3Q2fS9E8oWJ6zMDidL08ZI+Ksr++lG9nZD4idy4R2z
/Nix/5lPg5EGwH/w5IUz7a2nkolnFpy4Wmxtp4Q/H2uttYuxjfDscL2X/QQLnmNr
1gcSBn7quns7ghG4EXcu8jtM753myo6t8FGc2y6EdQmGV8c5pZmxZdo6H4WkpMKT
znGu1N06Qw+xbIlf2fmP5vjQtR80BXJC5BP2izkRqJBLXXjg5zPAe0DBo5JYxdt9
g93qwJvR9j7yNxyCEzCPn+fyCqFiYx6xpDSr7xlqtOb0oDqooDLdhejXPr/ZxTqS
xwMr3vvBVdD8PyNwwi8Zdq0n+VPoniqj2iB6noSVYjaG5swRdLTb0PtSCoCRRwZY
8OHh8rAwlbFV8xLHPuryWfM8R49dHj86hB6OGL5Nk+ebM6BbsSwlIA1OEzxJDtcO
Z/KRwU6XdhBPJO84iaHzBujfl0ODYLKMaEoX//mAJsbN2kQAFcCM3I+PrGkCHlCf
TiOvphYMBQ7x7niP9ekLITQD6A4r/iEMcaSfZlCvOcjzxnQO1yoMDUjDH8/iorzg
Ls1gOdNG23sJiDPGF38URPM3s2NCKH0T0dXcR7MIbHh2Do17UlcFgQ4PN1458jcW
XL5Wavk+j5zERjU1L1lKGzyD68i6PLrsVOcuZJLZ6PPTkDIyuKDz1Ji+Xyzucyjg
tPcT/7riEEIuHBYadqNG+jWTuY5rNz1fqXcQDy7YiDAiHx463uwSrgiBMDQ7vcTn
hNP3Vg6/h1zaTp/q9Wk1a9i6JWtNyKnUbbs124ldDAtDRtHC+CECXWBikEAGbij4
BDUm1r61/lTqj1U71iSwgcGOkNKujbvJ7DySVntr+nO/yUZQHBkyGqzAptYNDMbX
8pQ0g7AVZCCiAUYbWxlXblRvL7TY8b/nTR69jvbgOymnUoxLn7IWjWlJHjy8kpTv
WwcZsAd+1yMpXyrYoCHeFMkrXEbMHSlyHkd9ydBJNP9PQOF2M6YYEdluVqaNJebD
vpByaGOytqjInN8DACkJiHYBM7vA05Dj9mjCoAl7HOnjjR/XHqX5IgRPRz13/SXs
ADpccltRYZdSey4gahxzSS99htkrRtELaX00mMmm+5yZnS/gTwSufXTjAIuitQMu
6VoWjGI/pXFa3RYmkbfDfsVTl8acO7YlNxy9iH5E1EDvW0g0ChuBrpUx6/TdI7CI
8Wm6cCp/isLEbfw4bBRPXt8vG70BbRqi/rWui+Fw1G9x2pDaINt4Ph4EXR127rt3
jBrBHFis6wjkp/+/GBc/D75Bc21bqBwash0inc1RwuBBNBbezpmo7CsUtujETKSN
omIN4iwnxfbQ68xgUUp9KjvrHzF9oYwpzqpbo7hfrgbZ3iFpQD/XcaXhJFDxIKV/
002NN1W97ig2NopvinvNjuK17RYNpByDJo4ahJ/oxyzJmI2EHOHMtT2j/zhImBwS
wmRvUAaxrfKcuuIqydz7NT7lvKyTAYA7uA0l7rbKCD+A81awl6pAUu0AgsfDodtL
udHyiLk9EqZMpevLkt3HJdbJJ2VN3VlOzuHlgQeXZeLnFIFzsxM67mhoyofPVzFA
WnRntiWYXUYla/z7lMObvbMT9gFIZYBH92MVEF2O5CBpdSUiTO1XD2UBSNb3n5TR
U23nTz0zkvmc+w6g9YfumxFcPbEdGItGDSfRxtCUZZ5ZQu3v0Is4SlokDhBl7Q+S
h+6xw9oLzBq82i8qEekyZGb99MHUgEFO1Pjz8Vw+R/biIdZ9jio533dX2y9EIcva
mSaL84/Q1HRZGwjCLmCUaiGNxsa5B14ku6H3LfCYPiAu9xV7LDfYJaZuJc+K7U/F
QgtSTOVWTRkUqQtr02BttUN1j0T1O967FyXXcOfzvELTx32ldIOmC9M+L78AWDA4
utt6eZZGdaA+uEbUzRFDJ1V1/tXXEKum3FDCvId+ls8nzM5PmjJBdSoo9eCMzzs4
ct+K4x79Uk6C1t75YR8mY4nijBdHIrI9t77lgIq8XGMUMbiavLRl+ZVJT3g4yp64
9JRtmXbi+P+td46922+j5tGkxwa8ntqAVbXidifNlY/vbHXw/cMLTPBwyXmPVQhF
aZv2TH0aKJHzmeYT16L4Z2YV9BofDqyb40Ee8kLkuUQ81SAOQ5lgaQMYbgsZg3Za
++GQbZxG3zHcI1+q93YUOzqnb2et0ZSbdlOkjLDoyz7ESROGY4Id8IQZYmjk2pbv
xWzdSyqTDeJ/l6lOUS7w94MLztBw8xLD3KffTWZHUc+AQ9FVYXw/WOd4Q3feKsEe
24l0I4iJ7NX3du5CB6Xkonplre2n7GcH48cZHFo6ZHRXV02En9S6prvpnnQyzgg/
MLBG16ucEf/290WFD1bFQ6VLAE0wPQp4F8YGUG/SryEbfILSG28AaVpk5wiKpOF+
SsI2V1slsrPD1VuRG4FfSDhnHirysgnKwuxzhAFsfMd/nvMgUHf4wkYX8UJ7VoPk
r9DiOUHAkH76oyRh0zD+KU30VnuCaBS9MwSURhyb7aMTqLFa923Q9oWCUvBV6vmO
0HksFwlJY9SI/3SYdXhZ6IJYK4v4ssgZyqzFVwRUTK+hlGG6BBHjfO+SowWFZRny
OOdTvSF7TRxs54WE99UqACyN8AL4xyaDpwL5Q31S+QkLFRx4EY9kQvpQIxubmgs/
cWdYWc6/Hbcl3CPFLf1iM+rZ0dl0vnNWyu61H+S1GPQL2eBsyxdp2Iw3vkaxNLda
0f1ROv9EABquvuU+erGltmroutErNW+fJhiTZTB0ShgLU1rfripnNWKDM76E36aY
3SAqHJLgqYoSck75Z3N6Cy9YxSYkKK22BNHgkPT097eB4V7eoayyx7b0ngUXOu+u
XsYpto2mEGXwx0tREZhLoVPKb6F0LaNacnp1Ymc2JwQoOFFEly4stTicOmGQiq8y
8ajRa6Re4iJrRhMCFaK5+Hy1U8tUr5qw9A2OCmIy9pHe7LDgq1rqkgAfZwBDlphg
VAg3PdKdkBRD8avPUA4yQAxVIclw5/8h6F5n6LDtHyV49vgFtXE4YOjmjvUbrxY2
Om8u2DP11xshjlOJjGm+Yo01gOAbuIm0gkO+by02JaX5SYFa8LEUrq9m3LtRwPfv
2QP1MOHORBkmJthSeHsJub64FmIrqdJ4gH98HHAKZtIBiMmSmArLurCTT09u5hHe
MEjj34XWVmcoXPRvLQhcJGYwLR8mloSQ8i8qzWXn7pygUg04GSzIdHxMVVNsyrgY
WTgVqW1UyfbfMZ/Z+4cqk9CUmLzgrt0Nn8GPeNQ5k4YZjRnyN2/Yi0PnPFybTZ4W
yP75N7/9WPmKZzP3uTfmZe0aAlkFrYATxPXcviMsxCniyEFT5elOgcB6IwE8gg8f
ggnCi1yFKYZGiYG1Z7N5KNlqD7exJNRUjWf+7a+2Dab0pEIbppmBdv2zpuxBYq30
QQClNKtrOPOgfvf2FijGiORzFd3AnLhZfPa7rPZbPn8C9kYAzFGeGPv/BAV2hLi+
kHkoTSOmQ49Y5T/D+bD3Ckn+3i8bancK9YRsEzabQwyUGo8FjZKLmZxcBhL5DsfS
2cN9YcrCzLZ6MHc3SYdj5rQanYxv4+duYiQnQ1ahN2yPhbffIQPGUv4ICwd3WVUa
6Qw+Ctz3yblRK7Ci8KnWMIC1TNnHMt4btuErXTeZUa7OUnhgOhAZXVIKUJZzGKfC
yerCWYvMhgEd3CfTcO4+gV4M8lA5gGNw34cfkBHUbkdf1SpUgJHfWBSokbM1RvpS
kE2Rb4B1R+MfytoXLlxIUjhM8qNXh5xDChED6t6gzFtDvfBmYop/rT+8KCdiMGkg
tMOvEgBM27hqGuFoBQxqdsEGnmPkA0J+sdUtcA/cEF2E1PMIQvxiVzpHOfYfOJnr
1vLQbrLW67YfXeJfaMWnvqCvfZymXHsZivmNPF3iXPT05aaRiP3G4HUPwCeTWwVd
IXNQcsEuMSiaPt9IxLPbSeSr635n2mS1LOTRNu3jIJi2E6BLd2Yy1svJsj6wYxeH
MKEDDxdHUT8V6C6psFyd1HMizOx+Htb0soBDv8gojb9OEVC5ioP2t3BVkAfRoIjR
TL7qFf6vDkOcHVOqlV5Jd0y/zcK3wrLAqdONP5XAxrj0x/3cs/F9Uyu4eBCHCBs3
KovyqMKQV4FrFDbykZA5YhhDIHCJHv6sZo4VQ8J4vKF+Xf4eFrI+VdUv0t5MEaII
dwZtWsYa1P0u8re2+CMU8CuKANUozN/svHPVyTNXK825uQOO5YU2Q8D7tHj2VomJ
ockhInPBRiGPirf1qHmk5nEw6qiPpa5oAHWyGF0NK9enlaUJf8/Uv1tIJgsrtWij
D3LqLXHXXJLiTHLPTds1w8g7h7zhK5o7BFK/HXdSVmFJH53YMbiug8Ggw35m/H0v
0JKeKgcVJGFJa8tpZZAhmpGdMT+OEVMOAboc3fXgqZvT2gEh0Fo5mBOpgPKItDhg
kk1YCq5mwPrkb50Ffg13YasUndiRwta/R34ly1GUwXD/GB5hX7A46pozSDC3e1Kd
qrcHlGmgEsT1w+bmjtAERG9vyuFoMa4kPl1S8aWb5IwzljLoNxczpTWLKewEupuZ
Il6v6gnNhqSsbC4lR8t1lhEx4iTmyMtD5icH09plxHPB0eaKUIeDV9iror6Dh64P
t3dKLKoUFOznV06scfqbO2i6RLfvH7fm2V45mmgQ/qyuti/MMQrfnqPM2Has2PC7
ZrjbopNK3fzmzRqnkTbDXXwV+TjHmkWDhVehPJr0ilEAjOWnKxnS9x5OoSaOwy5T
dHAhKhtMav9tx8jFT8ZVOTF7kExvQaU7SkNeWxvWDL8RMH1wa94zuApYSw+v9+uF
VKR5Zh05FgJNQgQ/ctu1A1WUCstQY0sMDzdaT25CqA1ZtLTSmnAIXmWTuFp9rQUg
Ov91/5aCk5nxn8J5vT5azQC2zQPBwffm9GfiQgZUzE8qifyOLsNSaxzIpQ2K/fQ8
4MuRrWRGWHlpiVhAI80iETZBkgzYgVo6L4yZ/mDxQWYiuptmAusgc9cIwWmx9ZPj
uUozqQa3jrEIBDeYtJotXDgA8SDpEr3ZdirlJ8K+a6cyaScNgr4dC77X+jmKma23
rrpxBGelq+22YCQDAhuXf6idLOXrMv2YmYQwo5IjKKEWeaUvfi8OAI3B31w7wFrd
qnc2EllvglYvavwTZ6dIXKOt4wLMiy0bMSRT8ESsKtcIJeHs9m7jOukLiR0p0djK
WOBbGJnrZDmF4Wpg7Y0c11Xao6kVexqGhO6snLGqIK2wvoKy38ZRUCWKsvDR0b/T
ndTyYuGISNy9o8c4kzRIuoBDkwXrsBEjOdfEcFK+WUXpzBrj3bVkvAGX8uKde0Vj
ZOrjz9Ot2JCwyCcTvZ9tsYQItfKtMLJvrbA05Vx0hHiRfjpUk+Zl01vD6tw2Fa71
7faeHMYJlaz3QZD/ZPrgLjtUnAZSb3UidDWCa2WDfJMQc77rI54uE+hMxv4z2o7z
qrRe5GLYVZCfF/LbJPVPnoLH1nedS7Je24ffKesI32p8HIAqPObvBs5yRZbOiccu
RS/s7sOcfDBlLfluqLsPBrrXL/z2rzD1KJv1wGhDv0UBwx8AiJYlZpgACOQHCdrq
q/GfOB2dghnb26lJ6QByqz2/0WXuwBV2hsW4asvke+I4SmqY+fh+Qv4T/eT86QJ5
ATkiu8pgMEdU36W+rE7EQNn4sgoEGBd79mxkjsiRld+4ggg2MjMaF3CvirvDXAoD
ZJ1GZZFtKFOD33GkLomj3nSHt8IWEjZOBtxN1TQhwvV4dn7IOZlo2sXjaY/BLGxc
2kOHvylnKd6gCJ0IC4vb7gsxlf67gsOLdW+NlKU+RKEjbo0Ct0B5nh3v0h8crFj7
Xka0a86fb2LC5gusAkG7ztbIiImrRv+zYHPgXfMgwUZtpiAUh/0Xshc4yrau6TSA
9D2xXVFmBIjeWWkSP7m7sZDLU+qDdKT8gH6EnokP7z9C3N6mvT29NIZwnRGJO9hX
Vx1HVzM2X2/Kw17RoyR8zQQfSHR6wg2TSZ/Qgd3AZifqQPe6BH8TLCq1gZmmZxN2
nlBWiE5kSaGWLqqlSLunw3hTJ3p5rqinbIbVzQjuZly2iL4DMxTCkY4+oczS54eW
IrZHSx5mz0RxA5hjF3GowYNj9jbI57aS9XU6o8h2FW0ryi7jbGbthgswwbEU2q25
a/Ji5fPWx592akhGiQrRqHBUbCoIA+MSQ5Az9B6y0iQ7LIYock4pACSg+mcr/eDh
L+vZq29Fa8tTxfG5PsykKLjG03wXsZjk300pn6fyoPK2azmCPu21BZB98+DRDvB3
ZVHJvpWGez+Fk42dmZHi2ykvworZP34qGBTf1Gby8G+5m/2v/cUHMG0lxZ9O2khN
5svuNxDrGddxYBVR7kbgFcTwLrPdRV5ot3ecRCQN4v89ICMZhPtLwTw1ipoXADOZ
VN/ZDOtuRN1QNOh4+2fjrJex9YJeLax/0ZA6N52br6QJSyQatzyCNwWt1eH/b95a
`protect END_PROTECTED
