`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5bOV0TW/QOtCKqAWRrVP9mttkKcziaBuaMX/Pjd5yi5rB4XWVHUl6eK6hHkt8dV1
tZgYE07vOLYPjUAP1mL0rwSR5kmTDxo9Oppq8AaIGkPX5bRetQXpgXx8G/Z3+yor
hA21JapGAX7q8Y1PyQsImbre7oM/z6qBXth+hbb2Djnw5Hkj61MEyzDI68Uf62aR
cUV9ll3HznD62XJi/dWJOdkvoC/yy9uf+7Q6vIb2OUt3hqZ/xA2ZckY9uNCVuCY1
DWc3q7/VMsl6ZV8mnd9lKqRGRawps3MjC7h0HD6HL5+BqymldqrKcPLGa9xBSWjx
3+X3XPJqk/p08Vt+ZoWolcCQf4s5uy0XLYQg7Aey3axPF8hJgiEV06Y6F26WfKCB
DQDH3LqBBdA6gTphXOnql+jQwzP0OO4rAqhbK0Kp5CZhOjwqY4MQ8SbNMdZ2VI73
NwkmwQobKApqeJcExIlGACISFobm+glm7BRj5DXOa8NbIRQrrX3qbLnrj3CXgJt1
OirkvBKpS4Eo5lSin2+zUe3JKerbgQ8lXLH04sI5DKbLInVeg8qS/ubtkv/tNMR+
2vrQmYBTrBLUdOzIu0l8UBbAu43vxDJnzoI7a10AzTExImmag27KYcs4r5dLbupU
UJVtd4PuRmKydUS5wrlAE4kpRBxfUsDmZO1RyzobX0OzDtgcVN1e751NkFW7ov44
xj7rTjlv1tqK6vK5V49AKIMVRRplsWeT+8SwoiZ7uemvjCfiiYr8tYesOqW5NLGn
2zj2w7KLKd+fIQ/KDfPK4YMNDfgnwtPsu60RtAtLUZo/2wW/FnafWf+SNbG+AEJT
dRb2q0SA1Y16cmjTxd6Kiw==
`protect END_PROTECTED
