`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY2WymApfAigrGDuJ8jCMlvFNEcSFepP3XhuU9hTO8z8S/HXN+VVT7ymuHow4vpG
RiNU3/Hn2JgvCbDCtdwDORyNHj1Kte/3haBiNjA3hZJaKymyvPvcjbwxe+bvYy2B
YABgo2NwL5j/F7vMGtn+yIhAbDMy1dguR0znJlovVaSDzQALc1c6aDzr7E9ccQbD
e5YxN83o+AZ4VJPLoEvZNEcof7pw3bTqkjbb8Zz6enRTLEoHEVvq+HTxdHFykXZJ
B8nlAmQLsbk2WigntPUfHQjKHggaEhzVvASaRgVqP5rokOChMLCCPiC4xajizlAp
scudTTwsgn39RpPNKbsrEzoOwVRQb3dNaijsSbBErQJy6hJdYfBXCC+T/5O/R/zq
C6+SpQoPYB7CMGKetHBWq/a82uuKbxxqoERy3KT679RYre0ZW7HS7PcIthJ1ZYDP
dWnz5z/vQ5dA5EdTywV07xh3IyV0ZtImYLE0X8wwJOtrnbK99ws6/DzvoqqdTBdP
75wDp/7Tu7zhjzQuAmmemu3XJDIrBqWF7OG2YIbwCTWrCBz7Y/xBxKGtP7HZqpt5
Rn2wWbdJJBMkrGw8aPRzVPDrpyNYrj4nXtvSI6Qe58z00aj4UEJKnOEzmuSN+8e7
oQzyANqWdXIQCd84CcSypPc5B9w4xzRVUxlmJfy3Lj4lEWCEBvIwdVUAHE70cDrS
4WbHEvLkhln93lfVeJlJFN96d4v+berTZq4CzuMyns3Ithg6rXUpSV39jn5eK61r
gRgGLwCk/Qal9TAD8Ke/SoSM9Wq1PGv7n5a4HPgllbNbX351VYS2cGo3RUaGhwU7
E4Fv+5VTZro6hxQkZ0uuCrxzejepJpMN1T10+pJn5RCliXSGx479ixguRiLV5V7t
FPvgTTFAolvwm6zVS6646/Q7BrCKWXcJSyhnNdv5Bl2wWG+Mr1zzFmLF4kZGAJWM
YeUtTVvoHkOQxgSjoOhgXcTxilCknpr/PzMnAA8TpTTYyX2ENxfN/rf12JnkhpNm
H6nHpE2G0nAYfjVez8CJ3H8+f/EhUpqnHgl/nk+sbuKVjJxY7pAqj4Atjfn2uI5A
MhmMdOdV289a+d68/XejqmGFcDR8Sw3AytqOSL6J3GBabixTT0r4lzwZLGp1bC7k
fK+Po06bRaQDGjwqf9FpYwcuaXX4IkEsBnv6Nq/4DiFdL874PsOwy1Y9OZX8sTVj
enrpqD07pHvDvEwQz6ffOZQuIfzLQ0APJTLzO+zfBiGBA08u88PscjxjX0K1ZpK+
QifEW14Kae7SfpD4o4eRQfxB/oWsU8i1njp3q6DJK+fuhR2bt69hpzxgqdm9RSD6
zYY+EeQ1yqGbUoRt929J/71NnWUAD++WMDcrkutsjesKyoFoYZDIbTGdwxiz0qS1
JxvBHcRp1TNZU6ZWxEc2mGbf1lBtZn6svA2QCTyRyxO953BUo2MuO27I0vCPxa2T
e6R13BkqYWqbEOK9OKxRPYRo4/jAf9G/l0fj9rg3WcMpsDXXqqn+XR2s30//H/Dg
k9uINAyl89/zfJJkYXioo+txsldHvhHpfomUEk2uKFes7GGx9RKxt/X5XmlIyxzC
AjA31K/MDbF1IEPPRlyVIzYmKFlR5ADrDqed7sBC6MExt9OLgoIA0DMFeQONhRs2
U1lkYyUursgCOQSUemde2E/GNZVj08afw+m+xueRHpVxDaS2+IWSy//83Cb1bCFj
2RufMTWFqOwqVt61TTbUT8rrw8x9LqVZGafoqPRd7b8TdLn7ex1JcgtdCT1yxpcc
qMMaA/ElwVQ6EdKH0ZoOUhdAIPQ209rjZW6++S60uM1h7aIJrQ3S2MMKQo2ixOH5
Sr0oj+38agnn0fxdqw957ujJLioShqQppfFsfL2OEh99kZuHaShEPxl57fKdFgv2
pj5HhcCZgmsEKkHqfNCv7jRaQCWBKyYVzrlPflEwNSN7qYuKuDfsKlq4hByIWHM2
dt+wHCmf4QY79OlF+WxVRXg6l/1gm64bXMS1RStu9X3aiK762uCeRjcgpT7aNcy+
PN2zuGaAnsfhAI4JzIsGHiCDXfBM8DeWtxD8CChQ+KjQVYCL+MTTlYJb3ln0YgD7
R2+JBjSTDJT4W7sop/fhKebZpkc7jgisQ/70VrEqlBSRxtURKls7ulVQ7hsib+H8
NrdCNn7XoeJI6Qwk8+/PXvf6fMJO8Nj7Ar29qPMYJe2xUb843sDbTWgsvXTIVQmr
OjCx0caA3/vjZjAoyiXTAAAnAJfAo4FqFzhgP/hGkRKZCuSKXU2pw8Ow6AZrychq
LPWsQsHJKQthjm0DJr1NWnSNRJLdiCtnYjlE6J7RH/BqNwbtVYco2lij2wWZYKB5
/Rfqgz8Zs75xy826oekK3fYLjwlmpBNzeW/H+x4SeIqnM2EJmTmpQM+HEKP4innM
Y81VYAF8qq2e5uPjxxeJoBBdTE5EBH1gqhfeMNgJhPBJQJqdnkqKR1QFKnotLZfX
ZUWHipSFqZMu1zC/dWzMvlM+WLOvDT+83cUCLvowD59AtEf/ryKOw8Tb2q4zx0Ij
CcoNBb1EqAC4dJua7mCpw+Y61cnFot16y+XYg5cxeJmHm4gPjI9DiVAStbWd2P+R
bj7YjKv7gOQQM1Hv+Qo1w4qxw9MqV5AtizklTQVDM7VEdeliTpOU7xOZF4uPuS6m
qeMMzVB/tSWTXg9AwL0HLMJCHuG50f8drZxabj6mm1T6K/2IFFBpeWyiUWTHrJb9
AnL2W/MVSvRs5yA4t2jrz0GAxKFrMJu+Mb2AIq7+4QNFTGlgPO4j75WSE7R6YD4A
vhKACV3dJLElqV9uhjoiHhRj+JNTBYCL4z5KlOy/ry8I7iCxnTUCf8/0bpbAjI0S
WLRcqPUN0r/sTr1KJeNxeN3E/I/6X22Le6UPChRGPdbWUSQrIujQii/RKwjjqkW3
anj4OUnvLv+2ASG2JvejnQ==
`protect END_PROTECTED
