`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1vwK6stQKuwtqi9vxdlw69mayIhRtRrpB5/S9IrAlvjzt3F6hmlC82obDEcT7qN
o1NsH86lOuaqLlMg1lsJQCm89j5/8Gel3GBgY5MWxq2HfBDQUzlhcjoKh22+YZ6U
rLOcOmc5/c9jpie166p3WeUv/KGrVgHTjWq2AjLDiX+11lxenmdwJEOXy9mjqP4H
Yj/ZCop7DBgjXQic8bVQHFp59+s5pF3GC664s1aZcAe17/Uiso1GNyrimWWhwDph
DeMIVPSiu08KYbaDScZE6Wi8ZmAVX0ecSCzqVYEsUXEBPMqVXBBRjH0ZH2PSrEkl
oR6U6quDXsx6vHfVKQICexoB4Q+VX9Vb9bY7gSq5AlZBcazrppTNWFeoc6w3r90f
X3mZciRcPE+uvf9bo710Ef1SbCq8EXWBOjSIOwwEegbpr1txe84RbCyBRlkO0y05
lKpIBtAigOd+2kufWVIJNktmBWkjUa6WV9Weo7fzv9v4FKSuMTAxH19+s+kXAJED
X7M6megFdfEdtYTYQHKZAg==
`protect END_PROTECTED
