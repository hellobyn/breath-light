`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
It+DMAlJn6WSqHxXyF6TzfyVLC1g/TQq7VsE+5YDb8E7p+EiQx55OAbVFOnE65QU
6vNOQ3mUOlwbvGPUCfmhVXprDIq0Bjtpn9i3oYLsKL4qEVFFH+6k+UtFWqkNSpFM
wE5Gx5kdzu27+HYE01Re8Kx+E3+gCcNPeba/MNR9/a2M5GzLjkhYhzWNMs/99VWE
/1GoKJ8D5ZswyaGY+4z9BbI3k6wYPgS94iWloAl77UJ/iMK8F3I4eQg8F8aJo4KE
TQrtZCjqBgPT+bt+6PKmgdU9LgHJ1DF8cTmBYwQMdXK6B5beAbhHx/Xx3kIu4QT4
8JA+NAzkRchdMYS4HgzkB3O8faXbtVY/iX/vDOx+UJ0jh34F2L7E8p+CDqaftAJh
YjR44yiOqDgyChzkgVdfUYzYGj/UpVfWduj1YU3qAKObMARFT8Tb4PvEshExzwl6
UDunmKdbBZSwRG47zIIAl6jbriKrlcp3qzm8Z1v+TyMT6WcHNCAFNHQrPfpTYXHy
Xwa6RIHGNyl+n+k1rU+rZnmxPP1ySVGThx/fm43fThnTsOhLlbKAQMSYvE2AbGJR
AGPpWomjPw4q2Wlt09UyDkQncW5VK4RBriSEGJ7oTpCnfWIcX+OipSDNttJJ59LZ
11J6ayZn1HG01EIFlwLnpu1UdszISrkA90Yo92/t3zmztnGHfP0NYS71Oa+stT1x
+PqS7nIyjXINARG6+ggl+0ieGxOnMEPKIAf626GY76YJv4cOFc3ZiuvffG1mWtec
tzq4YBzAmk5FkI+bbIffFK4e/QXBYEGz3QEzFc7R9gH+bGSegjM5MiNUO9iqjVph
S729tSmK7jOLXEQKyrZ5TN0FXgLl70oq46lX6fG20rG/hZX2cOMO3Sz6Bii1cfc3
3z59qwu0czChgfXe3B+Q0X5g8BAWjK0hS1JtFvqQiZk2sZiWnfPpic0bQX0JT83+
LYa6OMCZtiAnmri/I0KfgwafoQzDb1aXSU83qZcDluNzAD3s+e+cbLObdXE2kPLc
kFdNc/dMRkTsIF75UlSBBNyseIywkmWZDkxfk9p5rm+xLRjxJU8xaBz9yW/FsqyY
B0245hc6NGbyJ9RXmrUNrAAJWKm1O3m7+iphO2Fkt+eypt/M2BqNJYcoAQnlTD4X
T0HywlQJh+HqPfyttqvkLxaxU0+DF447l4OEQYz4OTyJkfXDjnEFzSGXdZm9CRMA
wur3VQE7YUFss/KM6AWlkgZvBZIXfTL5DXKVORKij+h7Xv7wa4/CP/mXwbZ9oScW
lZCv+5q2ZqeawNILVdEtspTSnZzW/E56DOIgJF1yAswkqmj7Jb0hwjmz/r/y7ICT
yXtc7Xs7eU1EYxRNTnzq2lg4aqlR8qdRfbibV3+7Wg6nCeqo+A5GXu23zLlhqnwo
jJ6/vmCI5tPB8TpqtA1u+rQwq3bte7ZSNzSlg8TkxzsUK2XoWIfNx+sf3eis+sli
HqJoTowZMMfgYzqklbcndcgviqUm8SjX3vPGvPuMyfWhNKAB6LD35GeK1hW5B1dM
Q6I4pov2RhbVn/0aWuPb4wT5fPpCiedzxkHvpN1IyHkWkPvhmJVgXSMBf7hKljAS
xa4DJaNnpqZ5E8aZ9+eIDfKE6CaSjRUauVbuDDOabmp3IWQczpWlf2rIO4L2/r6u
dC9FCSQnkXmvzHxteNeRRqYfUWi7jH3jjYaoeEn6KqgrM11UvY2Bqsirf5VjaCCj
VLBIcXldRUUSJk4367PLw80nEeB26tFLChjMaxqT/41vOeusH1Z9AR47RzfOlZKO
Kt+EnMU1tF7tnyGl25fRMzV4iWkoCVX3lHN0ePpikNqyiaDUaz9xledLFRGKtVC3
y3QaPrT2lSsdzAycrLmy0gpO6bijV7YTUF/q1+90kfuyQKCim/ADvaJ4R/5CHbG+
kBGSATiut/AKa/B5z0sUrTFQGXjfo4pofH9M2ZxTbmT8apJtq0380JL1URjsopC8
cTb6GzZmItYxjf1xU67HA0i7TqYsUCb/XMBgpzAfWcCc+E62FfNk63uCkohD9IrP
6bJs8DH0a7+uEqKDQWCpAEFIc3idWc37fiVzQiMa4o/WP0/KYFgAQcIqPpUPq8aR
hFi6iru09IGWHq/7XQOECD1tz6R2FJShtN8aKpKp+prvdI4X9ldOgc3gc9I1cfA9
s16kT/AYPbR/TidQWfy0Tt3i019CDC3CZ/APBi5Hjk67cwSTKXznG7jHQZlFbvPV
sarnxb+eERfk1Cr+76ajQ4lLz1ubNphCQ+toJyAZwqrc6SlXTcFv/5Zukz+tQ3ki
8Msf89s0bKRW2/gVuhlkU0lbwFwHqpwEaLHfD/Joxh25LPKoy2qDvJES0Eq0RgMb
4P/9ir/auVHGyq49ssIzTkfwlLhoANf47pG6X8+12d9+5gRMxH6iHWB284Rpb59L
`protect END_PROTECTED
