`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyWyHxWzVpFG5E5//JXnMQBLFRmiFtb6Be4cBn3nL/JOXv6TNT2ORrJiJkDp78Dn
36Jp77Bw58IsybmUbdcCk6un4C3Bl2FunSwX2FY8//OQ3HRmXEWikmG4tcUPLMVP
s80j7F15FiZVKA1rk+/EOcq7BeG+izJz6DPZWkUzmU/0UbCPq9yiFN84oH63AoxW
k+GGWGeBuq1XHpswhbgJ3PHKhmYBQ82jD5vjkdQ/GRtjHm9AbhPM4KKTdNXXRlnO
uB5QYTHM4Gr4l120Fi/2Oqdwm8BGwGC1FAs4riDjcs0Cx8X9SFgdBD23153GhZBl
A/8fbdlKgysCW4XBolZBY9QcwJ1+OOoeCnh/1bgE737tv9acHrrIiBj1iEVax+Oq
QEOFbIWmhmbSTeOJJx/PZLcyJD1uc0wv6hzQztzJ29FKZog+JzE58kQ87jxSb883
X5xw/cYwADaNmckiXSR+XiopjMNYFE/XiHKBRzd8yMrX1WI042lDlBdLtNgovPiM
8SUXyQNZ0M9oNw2MhAjxALscBf4EjIlQNihNwxY1sa5kpEfnU7ntbRULKTs+RSwJ
akjf65uKZu0QeeF3yyj54T54kN7Nj8iB+c81LuNVfxASoNNWCa6P5e2I5oGv5pjZ
tiMi1UBn2nDvcqFExuglhZ/VbYaVT5Bl7tyI9+GA4w4bZmvFWdyLJiSPdqw13/av
r2xvj/cZnoMLPUDvNabQn9Jm9wK61BE8hOfPQcD7x9yiczeULguFxXVcHf40bMSL
OhLOl+Ko8hBn7ZDpYXLUmA4CvepUQd7EXCtDdhOzpYz2Nt+gQrpCrAr/Ec5DMXTZ
w27aQnOWqPMTAaGS6FOEBGzC/IKX4hPzDMscb2NJQtDzsITdE8jUY3xHshxt/v3m
5xtISHzT8N9s76tJCTuGlW7LtJvDvf9k+Ovh81t7mHOApLxtnzdYm1bITDmOYXA3
XoWXkvci3T0S3JWFSagZpwVwB3oU6hBYhCtsF/qe3S1yIHIM5Vv+7YVi4A8w0X4r
uRBKIad8FqbDWxC1tU/KxOMCj+F8xdKuLFdOtNcTX4oznMwB3SPYSXfe9KDJOfRG
mgokj20WhEKZjj8nmGMJlFV2VE1hX70cdC10Auq9lOurmevpBWz9eAzNaRRyNV8p
F8g4h+iUxBr7N9hfLTbQj50uaZ17sv41IYJY5ywH3j6Q5i57nIz+HdRHREmAoboQ
Xssvlpe1lpWsHPjoJPCPM4QPvybjXtGU/XJq6FN6+HhrZOXxqAgtEo6qXBVTVDlk
G1tt4ygkRVTLErveZN/u41FgKKIQ6UjxwWzBtpgvqeXer6AsDJCZgfBZ4XGcHmYd
V/WAb4Ywq8JsSQ9oIGUg+1vqTt8q68NjkMfoL9JjEcQJkiu7iRYaDQ+c0vVQnST2
DW+/3+UoWRcJZUlbV6Ut2L0zVZONkcHDGlTUWWM1HTMjbgNJF/JyFS6sFp0H+rXB
5B9Hr0dmJ6OLs5Jb1nMIPIPRTS9/4FZfz8u9ZWtKReVHjaUdAWf60Zo8gaCY+2Ob
hVzbRC5b7gELLhpz08n01FUt4zhig7nw7v0imzca8fodAUIsPBrYSlX/gO0Iy0AG
yinzqshFcnRQULCfYR3WDE7YpSUr7zbzWPm54pooRdfrErn/MUFTIfxIeywDGV9r
zkL+tC/WzyfDMU4s4rhRUPgrBX0ShELCgPDbcjwtE48nwbLk0+Y6RZsCYpTpwr68
yzZDi6cVkl1eXLPk7/r0OfWkbSDijF0kmmFvg3oAXIjUTrm9OJ8gmoTiuARw18AP
kzUFv9lwMFjcwl64/Oa7TkFR3d3jKiHrszbhVjeo9/M7+MYcyLjJQBPAkXSq4OEj
52ni2SFIruyYt/ZIxU9spHMObmZEMXCO6JpMRxrzf/jL/uW8nvOZGCj+D42O1rp1
dXKkx7oinDr72RQu18JqATzGD6ObrzAJjXxf5/1G29rTtQO07qMYJrsML68fj81o
cFQm535/+7+zXGdtMw6RsDZTfW1zf6/B2fDTMqff3b/hSpEaSnCoyc5X/nWsjFRc
c1+pjikf/hazzF7xB/ehc4ZBzNTg4Z2LZU4RkCQafRSDO2XiPDdIpBCLKWVG/Czv
ETkFPKIaisNhebrBfCFYjSt3KvSb29lTVGhuzq1lcjSnzUVmAtOR5kOSoUX3bLbu
lujZDWivOR+EP6jKeBhPHDNJkdPHH57C3gkeVR3GVpjst/19fhXsrw9B6Bmp7/mE
eH69HzNQ4eQN4YXI1WIC+kKoCS2fK6w5YsoBoxv7xXBdH1TG5oRC8PQWAtbUe8+R
NRJ3a8Jvr9DShgoWPOQrTYwIPJjzjX1Wyk0fBoQdxOf34Gvj2m7WYLGLIzwsb41t
F9DqCA2wf4BY+KSxAAe28P8Vari2BuElLz+IUHxqCK35yC90okB5pSBUMysgyWIZ
sGrKfgs4dqazln5NDQDhvEQrqa9Scdds4LMdcpfs2QaMcDDyKjWliB8e9Rf6MzIK
UuKDyFnWsaKnpxZwOazyDfmiL2a1OFkA4eeRHUqpOwsZlvUhFfrm2Tf6qO6Yoxgk
Bz/hyxce9vwse0obkYS5PuyOkAvJ8n/zaCDydws1VJfOdezIQaI5Yqskw0iVNQ/K
9p6C2cG4vR55W8Y/b37+bsEHFwKWvFH2tbMyX3sS0FPLHK4KiCyAlDzKKXkkymOP
goX1RvLAkq/cnrxsDSD4zLwPrK/OBUT2J987Pzz0kyEsnBl6PHFi9z9IWs7/n0V/
phQNi+KCTQV/MkAkBkjH/4UF9Zm5tN2eDsyBoO6sdzS+TgMpLbMOqRMfjJ+YIPii
5m73yh315PYH4Ej2fWtEM6FUNhsoZQimvjBaLR/Hq33tpZHVTKI9Kf7Nl6+cqF6E
Adqt41uH86hxNJAYF9nU+pXsTbYFKGFhyD5tXikcm0qBt/JDvH347xO76LMuC07/
gY9cZCXroyPNC6K2gVDfqGhdnFroP/GKDdqIe+fV8jEHrzlQln+o4MyRYarqXbCc
cVC2N8/kHp82yXJLt/sOjR8582W2J5bO8cdKWwI8XMHc4dEYGJdZyYfbaNggjBgF
49DU18fN3dipHyHE1ncEIr173dKE92Pepep2T8lzvUR0hoBcAvKX3IxWL5T4uRGn
+Wg2vXF7nhgDRsU/c9zRCV5jVttz44UTD1uQ+c2K7rCUsXNPBMLIvMyOdE2lndHv
yehlEP7dMdPf8rYeIMO59gAJtyQCXcZEqNOc+DPuEqR4DZpl92mrHZ4YsKh3grux
2tIkDw1+wbjEZqaXJP4HbgOpdSxWl8aZ36015D4if9mRnJL9RvXwPi61GtKZi86d
N6e6dQSUEMWC0nSCM6iAGFyOtclTs0qP4c5YzYzPzUH06KrL9F3jRzVnVXTQcAt9
V4pih3nBaM59uMjPf9DvbTmoGndXUnLmFGJqMUHLOcdeAL6mAPOUOdVHFuAfLp95
F31VnsUZAf4v+jjWE1VhRR4qBHfajdP5qYhLFEg1t/x6/PLEQor1fma21BHX4UJ8
ygNuFLO+ORaTK7Tj+hXChc/XEGowRZ2WC8zqfoQIgdfONbfeYmb0cyOQ4BrsjJlq
ztpsySoj5gU9hY4JzCpcbsKOaaWbBrmDMaq6W8lKaBKnrayg/bNbJ8hVGF+P3Oz/
2rIckZbb4UbO0nZZoGxOt856AUhEuGSREseLkSD3xTuR5ACbuH2jgQmgusMyeDUm
vajtgDD/q5nDgLT8YIsJUk/+sGifFE034CElKatp6Higtsx4K374WXTU5U4yAPgt
v9aw9kDtrKwo3/AU9S+01aExg/b5lzEI8TfhwOtAYbYSn7xSI0DWcgda5GTCqhPY
hDNZtOrCmKqoAsI5BzQ5p4HEz9mMigEK9QvBpBUuJa6iTipZZ1kK5vY3Ey8g/HKe
tNIpUkV/gMxhUlu3idl13tzgR6A9lSvLwvza3v88LNpYbyRuHX8YBk0d1X8FwsF9
4f4Hb19RCEon/h0bMTUYKEEOh1aWsPe9uwA28kJD/9c=
`protect END_PROTECTED
