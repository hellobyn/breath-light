`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+msLh81TZY1VhL1Bk6cexzvuD2hWTXP6A/lh3g6OdLYKTYZo3xDQ0zQS8A63dIUE
K4lfyJzdp+YR6gN9q3MEDcABReFvFgVb01LJLjtS6IC6X6BeYFt21z1WHzX5u/gT
Nky+rdCdtbupDd7hEyve/vtJ5AmHOmsWZJ1NlFMaL6zRZejcEcMp8DxOQaVigyTl
uuBYtMJd4dEHdXbZBDYuGbLA+rR467RtDH4InfOmI7HBqoxiREZ/qjNHZkuf1IFz
LLDrj6cUCWSRLs8G/Y5q7A6XOxqzIEEOpR7Nwl3vKgBmZKZk5px04c5yj22zeM2U
a2kWlUqPSsZoRDzY+16v7859gQJqeQhlrBpmjHe8MLAm0b25HHWbJS7KXNHlz3L2
cXhKjxNjIxfncNKjnBKMVDPzfB8tG5XxzjYECm1cxhcOzC4b1CTOcdAAmrMOPeVv
e8teo3HDlV1rcrQDL073iMO7zPD99hI35XuWmbVN5eoUWxd/KI2VLbZA6o948KIE
HmJYvt9af3n/seMR5QgKWiak+TuSk4nEQzAr5LDEyPE+xTJNTAIjY6YgxEuJ/fK8
3AgTGFC+MxnsBlrW/mkZx3M49CPYUxQQAkk+bNn8fsa4JMh7/GbpTb45TtzOemBj
h1Q6nB7gY9WItDRbHAnMnO41c/dvFGmBARAm0PleQ3EIvWhgpvy6JRpSQNPBJ59X
sh2jQHL9kZAEXN6nSgUXMw19O42NB6zpIDeIevU6oBjYwH5Pq4AFFbQv+XRoaEKI
wIcvOuGgMSHjYpLU/x4JYDQ7gtEEnOlDvtneb4IIxuEwzaJ1Gz2c+ZBOWhIRtdM2
hwmcFl2Uf/36i43Gds6l73n1EGSXx9sDUWSW7I0Av9hpvGMr6yoHlJWP6N84ox8A
8OWNI411d7wLxSv5gf5+zp1oLqro0cf+G5FUkffoZ5hiBviMhPPW99ooeJxIcJAQ
ds9yHRCjz4QsE8zTEr8qjoc3ebG+4sBzxfiZfFK2WP4RT/008x1IGqMza+bb3RUr
bI+IC0lf+MoUNuC9lMHPDAAPihfs1b+04ZBlEcmhtnE5YOZ3htxyYU520mZienUg
0rv3ue7KCNdEOqlkmsxifWFohnARrIGs2/1GIrNIWIIOr47aLX1kzTld3T7+5Fws
SU5G/EDrhRDF9QNPq+ZTxv+pwOXHyT/9+08VSlQWBSSMmnLPoVj+AJ8xqXAnIh4s
KCy9OyunLmY8tHG5DzELEqLUiBCuarv5wTtu6RAel2vOwyED+3lq2Mvvgq8wTWMs
9p8/rBgsjGd7RJAOfPcERP+1Q/txNRAbb4gjG1Mci3S+crTNf1N2b4UeYsTMBtEg
Hj1KL3/tjFa5cKbem+Y7EkR84OhSlVuiWc9fCz0w1lGSqFt/8wL6zs227oqiurwB
zH+CJOZYBs2Fe7woBMiEJ+ZEWsmYrrWwDHXNn1to/W0M6tdDAJBq3DsbTwFVBDhh
9O0SgKXF923DnIgbIHF/vUCul3Gq6Dqwv2a9xrqYTV1BfdfYTCZUKyt5RSoBY65E
Lz1emsgzL6vykB+bgmcaJDfQxx7ZmKbsKSPMzHFL41wvBf2Zmb7KgR1IAoFsjhTg
3Ol9L9JXjYgZ6GrUwlR7ZXca0mbOhThxuh4K/yziebME1V4v/hyWjIv+366JP55k
ojzUbnHupXc2Hu4xtV45BDZMM0rY/4vyC6j6fF4NKuaQxIYQJsJg9YhUfuXxOP2k
0s7sBDTh1TwWxG/5yj0RwgrlOeKeT22Ok5O5PwQBRZQUYN9HjeuDQNoFKXtdoddc
yS7+hU7oJ7ssfOHlTztipPQSN9WQYeJaVBdxw9S8jSs2Ra8P28fPdg2vTKq/vMQ/
PLd+X4cv8eMffo8ppxW0WSYAk6TznLN0vpzoCCKXM9zOSQUOjr8uQE0/mOqrXlzk
2+stIQsifWGay9oyexqal51ZlwgA0jrqEUbZ0GC88dlx9xCkCQSmpDjM4c/Mgkl9
lGhZwuVUCB2ED9CoEVISOl2Gd2jiueewXfMCdvQR1dfvMYI2dOUUGRr570s7ncyT
EegojYMxMiyGPTRwa19FM8FpLXdnZomfR1hFiSfbq2Eq5YDu2815Ipd0KWvb93+l
4AeDx3l4u8zNggYdlRwmr+y+V6hnqXwesPCbwdkc74zdGuKKo33eVvF8wVKKU3Qo
Ioa6MlLPwC+NXGDkp7wpWeVKdAECKI21WDhk1+/FrzmODyiXHAz7AlJf+Nv4yFhU
39PJqKaFHbi1rkfOJL4/2U/HWoAh5EYAhyXOGlXg78M1uzCvYJ2SACq2OHkQ2Wtx
7YYU/xVRKXGAQGPYQStM3ZQNSLRi+nkd/683uU9u5M+5uuDij3FWo2hu0IV/yYwh
ZKG/g52VAt0FP/TuqKmjOWeqvzHcjtn5FG8m8bPqHjRdaw2psOEaCV5OJXsVC+Fx
P/IwJKuQCvupsmekLC1mEKGa1xLczDfq31hfp6BUH09RwOmx/XGCtPWcwhN9b03b
h7vBqfWofXCpNiOE2LAqIbqeRW//yMiGeCMvWKbCyYLcAu/u4E9FxujghLEfGSbb
VdMbPj45/3yd0GhdytFW+Q0yMPrxu5giJ1X5kFRxfHzZaiCOh0YcLwx3qCXBuV9K
DPkpYG3OSEBBe/Db7zifXsrTlt4bIUJ+ZNzMeO0e2CKHu2gB7MoLQkWT+pTZGb4S
2EydCpWmmIG/U/a+P9e8c0ACTBaaZwgH518bpxOiBR2wQqTj2WUodRbnqUI2VmuH
xa70cR2RoClBEupshhREQYQf/t8haDkmZL4AXKHPJ20jzODB+JNjJv5lyu5Fq3GZ
xtNgDKQ0hWQFoYBLGosYT/miIYmwB3IoCWxe4vDIXdDNhVYACnDi31wPdjn77gSA
/+QwiVMq7ckCylrodxaOCkoJ3RBx4tI7naUm23D1zI7vcFimqfSbSKYitC6nIa+2
gQc9UCeA4iutjH3qDW/C8CoRebhrBHwVFVN6KIXDksY88wa9qfC74RybPpS/FiMa
BwOVbZDEuOj3Dhsv60DZ9zniQJXamKS7GLtbF4+3qkB1dIxM982NZmhodB4z8DGl
+qHrXimhVBAVxoHnphEV4VRhPpqed3d+ebUZyX3hRwsgP+V73Vh250EATqzfkSXj
JgWkFzCi+NflTaevO4RwN03vPLeKl2KdgCHbOu68oGQGjnFywHT4ia2hB9ZJWkeC
5FH8kdrFtfUjLOE4VOIHddxknvXQN5fJfiXAXujIkUj7xOX/UgIRGtysFxyenoaz
R8HV/diU/Abpm3E4adcavG8w7kueJ4ICU5QlhSqAN5k6mq1rLCiIvSJzRiQWnjmu
uEts8KULp643tPYxPvmTWfqqESlE1qBx/KDX1P1mzjHrdOCi/BsX8B1WK9ttDSWs
nuQaPDRpkM0LcrR/26wx5jl8tPc4hUToweyZl5F5/XwC2A7jvqJAx5HxnA556fCk
ZzRaFFlEHB1S1HvM0vt086auMMh9Os9YSYnDzCncvAh1Re19X3mLp7C/Ew7GlG7J
akRakF8UswEidiqZqfIPlTzkjf2Y9ybtX+f4DgGx9BdMlndhMaeQQYPveKTeMilW
MbwlqUFblqQi7m7dI6gCb/CvMd+XwqicBoMabTuCOegVnGpD0qidblwvodCu9xiB
pD5hLYuLKJtMZZcAumEtIdDaoTnMYfHUJEhCKuxyOIc=
`protect END_PROTECTED
