`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3sJPRX+INkBG0Yn7umUjt9Rw8GCCeWdke91sGNH5XBJ4Y/nVNXrcORKCLV+yNW3
pLiD44ULZYBvWNG7bPr5g4kFiRCtlxKSRqkkqZ1/CddCK3XUzi0D4eHl4n4BbTab
jwsP6NoSiR8HUxN1j28i75meq9dhh3hdjyITJC1RRfNryKhO0DriLvcAPC6ya5Sw
chFTdSRsBrfmXaH/5xJ8uvEfiHDeRSjivzzpeKuygnK6ULADzORSvGdl/QNUaSvj
ONMNQLXX2qfDV/caev+u9xQgYGKzuH0EZ3cWpwcoQLVlCI38g/EGsHKunvSsDd3k
mmm9IjI0PpnBAXxT5UyPfZIJOZawp5rH+YqNNB4gPiSeJ3QThgvy/QXlemBx9ZMC
25fPGwq1Ys0Y+aeNd3jPbFML2RzL3q4yBSFxGDKwvqNUDCi2L5OJ76UpnMkxzUYz
4T5lGUxuC0k/sp7DVsN4XwWaOx4RNtCyKuWX7zbY3GS0y2z1PMudE4CU6Tll7i9t
9KdiupWWLxcOxEV5AWx5ksZB0kL64aEIx3XpjfhvM4v0/4NblcMkAKmA81nB6sDF
xzpbEOHKgTSiwuoRr5N/Dm5yh859Bb6Mi+ZvXOZrfx68E4acvyCglDz4mtTBdN63
8kIyTd02RNWBbAfsZLg+8q6gDKaxdHtXnj8wal85/tli3QErU19pn/V1eYFsaFMr
cALwmFhThWK2CCbZNzcDIzrgmiDgqutJg+NB24bMkBw0q3m/BGDVOVZyv+Evv+2I
p9Tm3ZFL37oNHbkACv8JgDK0qQGf+DxLfAUn6txB9kZcFmZ3c/5Q3X+b2l1+QEie
ulMuzmBE/Xt+Dr+9MpPWdgRtQy3XHGBFHWBchOdpS2n8PzzUE7Lhx059iTTPM3SE
OGuZIcYrZ3Vc5OVCX8LhkdeAnDUcSNr3ci7p1Wp08AL5v0G440fJ1bQMTohAXfLN
ZgY/4LkVbUdYnib3aN74gp9DPlY1gIXkjWuyj8fb4zOrw2nbVCsGH+kpmwvVcsC6
LYDqUeja3N/yvTnnWnDMlzjVVqiBIqQsc+i4nMFPfEOfRPdogtcxmCPYZY6dRh7s
8kATcnxTzvM0lDDCJ1A4n08RVvVOpLjNHXHfVSmgQ/VjueE8XXNTb93hSatpkUIC
tlBdUU1ckq5pH7E9FrPAYFd5BUAHWCPQ0tVIxA45B0+afq/xGhBcKt15mtG9iC28
4DftJf9d8hRj42Jb1Ws8ph2ZesX2ygcTRxW+sh2VozQpWTabIBsjLRJvQB2+UxfC
geBFX1NvllHUgsLVlSGftd1XY1iyxXyPwY1TS1Xghq0BGdKLG4aE9mhdANYduDyB
MKEEjIQP4UDMWJzoowxSYoqLZHAV1OSic/Efhe+6Dw88azZwrBGWySz4dmQTqggP
MOV+5F/a+TPIiAe9vVTu+5VHHPZtVAP0a/c20Jj5Y8pH2eJu8b3/VMzAfkxqBcer
pizB9GGTPq3dGdmfUoa4lCBKCyDo5GAWm3LCVLO4CeB4neUXBrxAS3yos1VCl/iq
2ZoRyTKD4dxt8Ciif9utyTaJJ4A5CxUkJgjEpfKvfVEttXmDVFH4AX5mznUq82EP
RBbF6zDEHWhu/2cIV8jl0PpsCfkH0sY7Ji5I9JzW/YnT849krDfFNC1sJ16kpU3e
NUNmypWfRGhytF5aMEEgOt3HG+4EESyHD5hutiqMmclKkB23JxhZRmy4+pVhmJow
6WE9MxPzYKX622BtYinhjnMOtrwU2IdMwyCYm36uAw6fukYDMYq1i7DAVaNWM+Lk
dMV3xjTwLm33LxeYbm0iJgy8p+G6SSQf216PxYC4LOAseGX/O35fvCnNegyxYC4H
+lDDG11uX4/RHcMdOSV/PlEYMCpGHuXXUOYuWFY1vsg4pGT/sOAt4M0oP8NYeRrV
Iv//drkztzT0OlWzDhMrMFi+cNjDiWlb/TwJp5DlB7x8o6Q1hqcRB/kBStD0Po8d
DUVxIA0jVxon2lfY+FN9OeT/o18X5A4W2DLdULEV9E0SVXSKHxB1qDj1kOLR09FJ
I4LCuHUNdHPL3WITvVrInVvSoULN2Lcx2Lv+p+00urItaYsqpa4mCRr04OSmjS1P
iNtztd9oz8M7bV3IM16BiE2cEKmtWe9wZsGGpk8f7/w4H9i7+FBM/QMexyVzyPwS
fRXZbg9tCZY0+MhjJW3K5ozV2SpFPRCfkjO5FVc1ue3aip/G78qqedPTEHAzRbqx
+MCD7lqj86kghjrJsxlfJ948ZOcAnvalKp/DoRP9tjW9/F6BuI/j7MSBNtHlH6ti
VXQcIe+ljzvkZUMw4Qq7RBcKhSUX0GOCimV9VJPr49EsfCHsfIVlUauZ1bs2Zu9w
PFKPTslC3X4QAotp7bDfo6+qsMA1q4eJfvKa1gjms+GKqJrIDIUcweE3xNu2LwNL
TuQfdBaId1LKOHOp9zI4Ocl6Eui8uIPMzb/By5Wrzfmk0qXpl9NnL0KmXm+vhPRt
b596UG0EEv5Q1SeZF+aA9A==
`protect END_PROTECTED
