`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThNU/XB7h2SR5z6mS8xzUK6ycssrF8Qyd23MX3MXsQLRpfZSIBZWRnYb0Sbh0Vx2
qNFVJW7S48cccKAC1wBii3gS1aatK+j9M4TAuGiXzN0oITT7DwGAD8g6yDC9ktMw
RnP1AsRhI5YNlDRN/h34AD/IOvJeveL2L3hu1LzNlnSKnQoe0zC4hCbczAzzlF8f
ToRoPBFu9K4KEcmbXhmTJ5ufsTf6j/jx3u0hptj69vR3atGTsHqCGkYXeumcjNFv
VdOUblWKfqYZSYUVP5i2GNTUFBVkJ0fsXtIOHiQAHOE+bb5td/dNF7MWr4KRlcQb
gH8tQ6dbjbbowV43g2NDHc+hUqNYH025pQ8hZhDQXC0AbJImVbUu4cpf14ud4jCg
8GnY38uyVY8OaJqQNfP0rc/YZdIzQH7gKjtyF5rs02pm6D2TLiii2qvuNOhs61gG
NfDeJHyYOOfAkDkz6h88QXVSs3dtnMDgt5SkTem+eMQxJ0Pj1GAE4mogKkXE2/rU
iP87mrZ4hXIDQhFLmOryaGgIXMxcHlAJmBNeZ34ILteytgppLZWLcWdrHmDGI9ob
/siXeoX9pGbH4Arg4L1iP8tY7AidQz8SN0r/3z00cKMELxNks04CoLQojMHuIaJB
ztFsLR1LTlfjMw8iwNhtmYVmpeN2Q517anrYvzVRBux8zI68A3MNYrlcvqk98BM5
yUyo92eK7G5FFdHuZPpJUXMk+e95bDGaOqV/Aom10KsB6D6u3n+rtSdjeqsCv0Lw
eGK0SLe7WGZMyRsmTXB4B+kqm+ywferJuLcKADQMPx9T9TIusoaFhN1m2L2GpyB5
O+XQGLoNn3wPzf19do2qBaJ3HeaSdE8+azUmnxp05BoGwALM8pa/DcgSnRtQdzep
xYfO6Izm16Iefbi2rSz2no0GPPBvXifvbQLmI1iyMr7tT23rhZmPsN2eJDmQ5sKW
S4l2u7qp4XGdt37Da4pCwwlJkwZg6PORp7q022grJG6Aa2n7ANZEbYS60ljgtONU
b3e/pbHQea7lBIhGC14Jkl+8pgdfGAYudrv5Lekhbqxi6ROw0+j0xN+SJ78i3Cb6
ziFfmO9U2iZyoxXPFyE6/YhN2wlU/xOsrZqAjHVno5vd0wnt4IETKdtD9HWPwt+k
c0eUdeKqkiwE1Akcdky+O8mjK9yAHEVF0wX1V91tzeLTUfaP8oOlbUoLUAwJZ+K4
WeKw7i8MpENG5My4sXn9mN5uGq5d/shvFDwpikUVJD8blPElZeHPAt9r7Lk3aVFB
meM3xBSuFIecxpBBzOHu/cmgUVra5m3Kzj0UjREpZRcV89Td75B945c3zntg/s5t
j4H7bX+N8pLYSucwYCjpKreZPoQUImUEnMOOc1E8F7w9O9onzz2IWx2KiWnr4q4k
Mq6os/NzDCxLgiSGSViBw0hTNoQ24OklhpAoF6usm1XUCKbXmuUt+Lf2g8D8+b3v
mIFqlJ6WfnjdVh4ikD/b4B3m9NBbZpqXKBqKSQzs9Hs2BrJ9rAc4hpAp0V8bY6lE
O/4k+YVUXl4nsyb1LHhsEPDBl1E7B1U23SJyaE4hvOVfYZ73p2nGfKVzIJK1OJuk
0mlXs7jJXQWFD9/9NqdgbmhVX/+iPQ6Aaz2W6ikStaRifYaK9DEYKC7npltlZRAI
tJUBWlaY+3A8JkuiUl3PBWvU92kecut8WmirNgi7vctI+3EO02LcWLHOA/Mw3bvl
kGL8QmrsnryBpWbn7zvSVYKqzwdqJxOnXwTk2eQuhs5oEcqgzqwJdNgrigb0xjLj
`protect END_PROTECTED
