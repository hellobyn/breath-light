`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yqB7qB2pRSguxz0s4pe3jcq1+Sikw7lPbtMO7QjJE32586ADkDrEZjN2Rqyesb3E
NNrM5laPSGAWJLRSY33WSivx6D6WTRbv3N6avGL6ax83GBU64owC2kufQgd+MITB
CpPpqp8Wzd4OP7H+XH2khmH4ALa37LNfWTP+nFkFTyIOawRV1JC7uqnUnW3xki8X
5lI25opYUJnQmvnxbCRTlcyNPyKxnriEhRkYAtvFNIGHB6aHxbodx60gP5dwWVqt
MijE9IjXbIooEG1rGHpb+8X0QyOg7/0FK/PyyE5CaMm5CkX/7aTey1/o7kzCMkTh
iiocCeEZ25SolOC7A1jZayntou5BqgGYpu1ri6pdEmNv4GMz/t4N0olOifAX0+BH
P2QsfCylvR8Ou5nPKd3gSKrtugM5QVHluUH/X6RVb0zVTjrZn17/Tk+oL0FmvpuG
8Cy8Dou26FwuDgKcAZu/hA5eUEhG0xqEbmkND/WTLpBXRXgNGy0kfCnYp2lJ7X2n
cGUSdqkCd3O4hrdUQwvzVCX4pRY3h58+wqMqggVE5/LB/4pB83Be8bCfMz+4euXA
EqEXFUoZGC9YlLuFG6xH3XINDPYPcLccXzsEoA1bSBGK8goSf23vITcNADwV7WP9
0K4/xe7ncK9fJhDO4iRZ/t0LtDnknOunAyz58zYzGhe43pC5WXLZJpP7B3ZCMr4Y
ZsTVupdGceryofMnBNDq6u/BQPIedjw8nDJG6nZl2c2Rr90SHhCIaaASsBGYYNMu
2c30vHUz6+f3iMXX+07hTl9YL7A3hBtCHo6ChG/7CzgJvgb/GjQLE2sW4wKOl5Ff
4WsoBBHmfr/m6gw2iCcEbw==
`protect END_PROTECTED
