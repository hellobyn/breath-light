`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlFCjCWDSAcJfImhG03WeYMuvlpf5yfVWy7IZJ08q+a0BvafwaQNGhNzPz2XRqz0
4F83iHeYUiiQFWEaijuncdxWWsx+/RkPnYYRrB0sGXdNIWzt5G9CEEYlMOjW4Eud
Y2HIVOpN6XtdsQFmT14b7eBxPzfJVrw09sgnDIrYhMaPsYNyzusysW4LSL2oBTbf
`protect END_PROTECTED
