`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s94QnbY/wzG47r8UpmCTG2IcBnjk2TghaQz63a0KAoeryTxFmo0uBMlWkppPj9wY
jA2Ug80vmct1lJ9EEZFHsmrpRLkfw59aqRYLaZHROvrKS4pZRFPQztjO0J+OUZtj
H86kzlydVj9HFWPr85Nfu+lUT53NvtxBbGNimgOm6j+uDczwmojzE9cKcrw98rZE
J6+qhZCkrp1W+QHrU3dcK1ac5ci86mT30LY3uLZEq6SzOqsU6KIy/7c9CTF4KECZ
u4dB1kOW923axQdvjlbEqxsfgoWuayVAM10aLMyHIgBQXkVP2TPx2IUC3erz9K0u
7Zf/mZfmZc5N6b/ljbvuzBNqOHAuIHaVlFgDP9/33QAT4JvYbdaimP0gi8xL3Dk/
u0uAErKdzh/NPVKC4wDcU8bA5TOqSNtAaw1mVEMLg36wR5JuRDHsLBMHaQXKlJjk
`protect END_PROTECTED
