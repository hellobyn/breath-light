`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5eDWzkma8Yb15/iJZBtSDkDvNvoSXkx6QY39/03cMIGtyug7p7nk5WtXlgHb/vK
gc3MFudsCyHZ331kgDHth3GwHnvCPaQ3QfnLTRT08gJqeQn/lb41AY2TZft9IocX
rCmxYw9vWSTWBjzY7xGRy7xH3GiRaUDSC6ThtREX+0lXy66pKZ6s2RCBgJo6+mHX
CGAE8keQ2yVB+hNrCPZOkJ62CH8t6snq4K6zP8zntJk6jsBS5dQuT52dawCDJGnR
4dlJHqpNux2PF+ipYfMhoM3QpbPkh8edWFNwf51uTla0R2TrffPVHAGJFsAxaViN
/Aun1zjzXyazRCJzPT5Lk/5v9CoNjU2m0DP/M4JFZufBiVflIj6P8usORGbtl3cC
v/1ZMvSAe0k0sJ+F+88Q6qDEgIjR57E5r8+gpJVv1ciFSCpsoIYTSille7N9N1DW
QWkr9J6oRfL68eqHjGipbngnzwzICQ9Zr5YdFtP94vCYI/kcUngEK52oraY0YtB0
3eRzXpR29+hdrW+pO2bls3BdssyY4Q8yLmWPG8w/tM6OUrvzQ8zN00YqVBkQ9oVN
mokYSYSPN0eU8iQ9dkXo6Bf1pJRRPtxbxaevGXSwCj0hCobtSww9DD1ZvW5zz9Os
F3F44fyYwd/AP/YSjOEw78ztZEU8ImfhmDCo0TrfkfZ0HuonRkgSTn3VPVDEVYrt
vKKOHpX+o3Wh4ng52JPB94G6O4tIADcrsnJzBjb3pBj4G2FMdJB/kfQnyUscdcKG
iPAimEymsmScHP57plLwBzXqkJ60qN9BonXfKb0mGeSHk0P/vBEkDwO31G3jFuUu
53/4wypCOZnwBdWbFAysI+zwhSRtLyLaKYdS9Dd3tCv+Gvzu7iFcEnjVHqMlaRE5
i5TgF7JjJX0ZGy9e1sRvHuDra3QH1PU1/SdczyVwZ7Fv+q7N5FEmZEQwoElQsGtb
atTGdXcbYWvvGTUlkkVvD4kgdiBFYLKTLbA9QXvdSquOk8PKcD2JIjFYNKPp27iY
K9rlRhf5VepMW4fmTeJdAHxwZQIKkKPjE3cpfV7G+Qu5Xtr2qHeNjMeo9HNdIqnJ
nQq09SGUwNIz7rgyRIE5E0wZ1j4Lr5TfsKhydhBDn/w7pNMlQtFsa91J9XzQ9sGi
sMnpaPsJExB1t/ICGoi90e3TiluFdLvNf/YhrNPJkcFPmhcxW8FrQfOBwEERdkQu
f6b6d5vyEzvhHrbDSW+UDJdwAiRr84dAu7JdKDm2RSs36O5FKfS53Nxdk73sDthl
5dFPtYwekoWI93iYMIL0bSIvZruXI69Qfte4jWXPoIQ0LmY/gl6Q73OGEvg16czN
Qz+uaTxUIMWssZzzHmbLToXQ49qtgl9KJgscmsFyPp/KTeoGQGQkJnMbUoacj8HS
SDbROHIF3cP5MfGIBks+28Ev8mFcuvqXVT0jFGpJXhztAX8wp9I41rdKkSL+AuPP
Pthv6mVF5b1JIygTDPRS2Hp86FxybO5hxTOOht5ZpZ0a5vvhj9vQXMI2a3hchu6J
5kKHLrk8NcDiagIogPrZDjscgEbgR7YcGGzFqPWV1QmuXbi769DZgukkEzUxIaTj
hkGs5Js3WB0mFr/AJ6c+5h1dq71PMPDG6s2uJXiRMRfr1PzC3cug1M2jPbzS7E9H
RuxshvGJj53fxX6QjFvXMuG3e3AWVmKiSV7kKB6tTq3syH5xyXxL457Rtp/f0Zo5
BHAmSbi/u7mgKeoOy61P4OESL8um0j9ZRBh3341yIVM=
`protect END_PROTECTED
