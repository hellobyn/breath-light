`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGQaGKuYBNjoI3FU4QdffeatIw+oROg6L0JBKOv2OEwod1eN87+QbatJOwKpS59b
dXx8t/sbmmKouQHUq8jjtERcQZu7jdQfWnYzW+ZPydTih8Wb5c4C6NyuhCEFyZti
hicZbypANZLptVAgDOF33Rk+LFGbuT6L5wPzbsDsPU97thGPzPyqgboSchi1WUYM
niFQwyriL/hVE4J4FmfjgFBLVYGcdvq6TMis3SuUdPwydl9JUnXF8OFupS7isylJ
zD4RubVjvXn6MaDlyqJRQEMQ248iprvB6fjtsgO07kdwOBIPF/7i1KXmA/49vczy
3UmEbN2DrmO5sfqZx1aX/X7jFdZ0c5ej/Gxo+5fDXvBsAdKpbrfftCCMnjCTjF3B
9vi9SchvrF86VJD7JLlM9I3JpHnx0Q777xEc1xMFtYfGjHxvZZpxEE5dY/O3lx9o
O3Zir+eiObU9GfMN6eUrrYehhxa3THyjsV26pat73QHMHQMkdTUZ1uBkLRC4VcsK
M8MDYJvm1iAhCwNNWNy8nLevfqIpFPjr0iHgg5zfm2tFWRlpLMAou3xAcYXVC31B
RkSJTsMX71LzbwBrx6Kxau2twfEx0Ejoe6LJi2QCTWwctli0qhUEIv1fYb8Kxdg9
yqK4bMUuAspFMcANEwaZg66XayHQa5WDpSpd+aI7ueWKzhd2Agyz2WE2wgKkYLJa
B/Wd9P7ChYUwq66QOflUbKTBPL/gLPhHO0clY+fsEbAf+ZKUIM6t3p1pHLz4DM79
Gz2IqXNdWRufFQ67Y3RBC+P/F4dLXFFUUMROjfKKM3gNBwSOrYBuAoPUtziyf5FZ
1LySUG8IsLC21KH7kNiPJw==
`protect END_PROTECTED
