`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
REQr7SRZehQtHRWqqtDOrhRKBT3wFXg1PbYyq1Wl9z1VSE98htJnEGUKySJ7hclS
+LuANoQls2kRZBCBKSH6lwt6f27JZ4INvmvYGvSmjqm8faefKnsViaOJuHPnHUSH
mNM7eRvRrc80UovSgeazCn4WEYHQuyVPFFLebS3/eJ06g1QJs++mlritrkeKgNyJ
a+37WFeknvumbuf/t5acKniqHArvUJ6rlD7cVjlhWVax9v1++7FifRqreEL6TBTK
b46Jxv3cru92Klann6WmorwPh0kviUU1h3t9FWGlQ8iUBg5jhdL7A1tt52gdd7Zm
rNjWrvGhaNpwPHCFtyC3C317+t+8r8QITUWQnVLYeYT/TySiBs+VL82pjtBdkA0T
mfmb2/jOmrAulgVACLqjCy7xSVHaS5k97lfnnTMbRypgo2TUz5vC9PrxlNp/e5y/
ruqQWehMpIOwoU4aQEVUZ4/mMkOiDDxFswUZiCcOlakMgPGOU+elQDJj/IDY21QR
DBcOQ3umUHPMu2R1i3Ru9ZCOPoiwE538FC9oQsS5RE7AOCmFe2yJZWzqaqREXFha
3tSaq6+6yHrbrSRkGcu8sptjmVdGwXV64M1otpE6c0V8m4qfgswlITNoxTtaG/0m
/NbVfHc8v7KA/kS8PHPY3/QYW98cKFlxPWYQSjVaEjSzyEOh2eA0bXQfXZFJ8i2e
E6lJFgOY82quapwwZR/OxXSJvG2eBRRgZtA6vujyM3yPL/cudDLzIohkK1E9SglJ
+ohl2kb1g+KZwYAQ0Bil0MFj8ld8pV5P2Zs3fVUW5PRuGXPUcEtzg9Y0AUrHsWdu
wgOmKvs5KQ2+Ys16RPqbItvCBaSzg1Hya+ykVyasMfx9+FqwHALW1UtPE2W5WfMm
qgyzNFxaqjP8q72T/hoJWxkAH/FOQd4oRSKTvDQM1xuuSvjWd/cPINbxF8Hq1exV
UPDqCA8jch6RxqIa85RUu7MHMYnH0HLveaWTMDzKI6nXqAx8V4NY7NZJ+1m35ccZ
yoM8/OP4wrx+FEWryrY+hg==
`protect END_PROTECTED
