`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2ixGvjkCrXxSZ3qRhqwnDcaD9pGZdAfw++1ry4KElW/EC800baYppaw51ZOSDAL
MOWP5XHmVBEQdsr+0f3307/BhsYKnO1jua8BWTocqQvoLbNE2OqrKFlr4IqKV5aH
ZQHbBaAaxR0Vjv6kbXm3kzULoseiPFKiNeG5hE6vUZD14w8+Ahz5BjjuILX20Gs4
2PuXCHVv6W38EEao11OXYsaCJdcrOCPXqYGX9dF59gEpGOuKzROHqG4E/y61wuKq
ohuXSuo9jYBR8jH4T/OUVb2NBEp3dlollokiy+PitYKgrdGHHRhAT0CTjXhbrNU0
KkJXHmgitgPN3sCWpDzW50Y23Eh3jV1TERprj6GZBfcM8Qie7uaiPKiS4PIiskia
imkRVvya/IIRzRE0IOzE6YmOj/d3szcj16Yfsk/psCMLQmfi8NvGHVRByz6VYZfz
suZL4jhfPfELFfCsQ9BqvPSVIYL8PJNYo2y1qrZ5r0Lv9KguShKBNHCMzRuk3EN5
9efx6iHk27vBQxUiCTEnJ5/5D7MD35uOgKnkwljQ9/e5EiCB4RiN/ZjFjCIsu7dZ
j2F8NVnFA4RDQBlJPbBReYLaDtBxSzHBc0gS0o1XUH4TyNb4x2mvCKuq90ccXz0C
WDARJ9GwWsm+T0aJfmIyKQOtljRlrUI5u0Fei2AMgVmuiZiizr1G9xpYgREKorzA
G99K2mKj+vLRNBDK9l2cIOSfrLFEZs/eZAoM2clRzOah1iAjDtKQl6iiLRlNApXv
lLCmYZ2mrm/4uyU/NCozSTlaungcupyfbix8hLnuaWTQs8Mzs/MdimsBWE1by57F
PJSMgxz14Z7cgVhCldSkGQoUHdnJ+9wywLf7oFAh99ayR1HM9Kl1JjQIrfxxYeE4
/cZWob57i7rsGN3gV/w+fUyFWwl55iJpx3/rHcmLmUWCQ3kyOvCs4kW9CyBLUHt1
qhBk0JsPHEcJvTJF83K87111C86ekKue5yCYtFTtwHSsFoQDTLwwuxR9x4b20WPz
seA2IpbGTx72YwPdiqJ9fIWEvuWW2TBTH1ATJwH9RHHPWD3P5pM8wWL+JRGZK/n1
anH0yYojAtm7zI+IQ7Wp/KZ4u3AVYKNPwbvTEhViDQ1N3TeaVntGj4w8OodBQgM+
Iz4mP9YRlcZLFeC1yUsh+zVkHJRMqhu0+T12FO3zHZ3rMs7ylTORDYxKroR/DUOK
fnisGIxNaaEf+J1dU5rawfnKIUdYCa17a/Y3hu4cW0FTil1nzMsFu8wdIDKtHtLh
F3iUBrBb4DLjvyG3UXvzzspwARjyDy8WLXo6F6Z+vPywNNZ1xNyiFjJBF/9XHwVw
hwUHNgFkCwLEtQcDWVEkn0FIe3vQlJV0vSwIkwrD62dl2acpAPe2MxS/zTHS+jy0
LrKjgxvd0l8rDJj3MUOXO6C5dQH8bqodB+jqljbjLvFsU4X/YfNDMclVgrPmhw8H
1AC8swccq32c9iaYhL5eD+OMUAjNAS89YAbiUCv5WD9qJeSBeItI30j2B2VJVnSD
hXzivUFrFgWn9BgjPho4UEWaZk9e4bY6WC6xUqTIxkCYsxV2d4iqS1S1Zx0GKPb/
WMqeMxwf5ib7WWaLazC8vm6mYat6AXI6TMmLGEZP7PCB5Kxr4hKp+KjlP/l5YgOd
x7GZwniXkN5RnQDZkV6bIR/Y024uxPox54x9eTTSLQPt93Hq1rdb5W45n40vG6Xk
UOLZB0B1GLE48NWTj0+c9RGPRDa+oHuV1mQxdW4Myg2TRgCfwPKzmx+Ra5EWIFvS
6gXunom+zZIFdNIessju9hOHXkIhMesQHS96UdkFCwZajPlWQBT44zTSJznLPGo3
36f5QfxCAs8cbDnImtf4psJ1M827gBwYuR/hCxLwFpz3wd5Omd+58El5Vq4hqYns
9T+Tf9ftelciErWqlHEsTfhRmJWhTPJEs2ZbqpiziskjWc4BkwF18okGBORuLFR+
3e4Aa6K2JHcOEztCBXm7RCiamx+IsDT6YQSJf4nmAOs0ttAmPFx+OCSTSgtlf7Tl
TSJBg0rrgzWw/f6l55b8qN3iOur3O9V87Jp8AnGRwf2YPLzHj/s/B7XS9KIeGXSc
m3dg2pK9Uzx7Y92quf/H50jA3Mjt+i6YeXfwp/YS1Rk0jJsS/GL3mg09zr7ytxFU
JMjopvk/1Uia4t6nFmNshxy7OrNQ6QvzoQfbOWc0WsamvpJYlG5Irky1l2DePhZ2
ppEsHiAi2ENAQjEmUCkF35N+2YsCBAq7Gk/24FBZlwanq7suxvmkfMKN9kL73UGY
W5UaxQ2lqKz/8DQkAyrCVAx/aE0EbuhOUMOPdbHfJEoQ36wusfcTxwE9W50+6nls
WIOtJ3/o3VbsIEyM45nZ0Jnu0po4ICmrEp7QWcDui9u6P1ADJhzIfWLeip+hYnh/
QFGQJSM5paGzU1WKwDU3YeaetJIvgbAuF9H83L+M/fbratyLcOqwjWnBsmj2jt8Q
NS4aKZVVyjRXPpdCbhaLlDtb1w3MlK1CCPDlTDFHi6aC0LOMDMZrLaBalLSKpJUi
5W6CSJcm58Ig3GUuwtCHzFE9YakXTwSSKLQUleHC+ULfaI8kN8BGc0f8Ovft/3wK
HQlYjSk3bjxPAHP4jx3xm9blaY8H392tfvdzAg6OSaH+GCA9Fl/XRv20OPLsPA1N
t8kGLKwJs3Q8LAFMSMY2EMgI2Rv/tHdxhspxwHpTwD6//G6OgDg+zxkN5U7eU9M8
0TxQ1FYtO5fm40w5lZI+VLw3JIVbvGuhabMF/9zR5jCeVriTLGBdCJjlwGIbkjoZ
85s8UkVF06GCHRFscab5oSupHE8VOQkkpx30mjVh8E4hOPXVdf+yHH0DyVexU/ql
5YuMgfuYuViecJSS4lZvsgCXFjZfN5VutoVwZrIbt8PkUVyv4aWG27nDb9hUnpgo
+nTa0AlQ/b2irDbgH0MJBZFeDBMt9Ru7E+8sjZ0doOeaQO05db9KZOWGLrf5rKNz
cESHEjkwjqBPjds+vHqtqh2iol1+NOBoIh03d55dy/nE2G1i6hmX5iuzbFDV5EeS
5rzcnMAW55WFXYVRJyVkLR3YbHkpQEQ+EjfrOBvhTe/KXerggib1gWozdR0O8ghl
y6Hp78jHO4HBHrzU6Z5zO7bLwfFRMfXe/gzNximC4YdJojCQPhxkPoVHxyd/JVza
Lz/kmpZ0YA3pNiNCR5uq1LMmHNlI4OfjaLFjrFEyY113XMnu4ifN/eSH7qS6K9QC
4HnVVkyAA6yn0oIY93dbF8MNXwZFbvg2qu9u7qlOfCQ34Eim6SnllQi6TYtZdcsG
uk04yk2UvqMv6+TP1NfWLMGVAZ3DTboW8ArCaJVP5hd8IFKUNVRn+5qydcW0qSgy
lMMge/NDcA11CjnOqePozM6BYQs0M322v8K9bDzEMhEVIYuv6X/CjGSmqN/CZqYu
7pjIQKhAV42AO3EHyY9NunwV7cI6LV5w3tx83P0h2nR5iXJX2du9ChaTK11EZRy3
iCGaEvsU7WQGfO1aSkxEzbOj+q/DfoEUNWRZobQftEdZuz4flqdwIe2Q5ijzs6zQ
Z4X5d+g4IMLp0YAc75q368yluIs/zVBnteDAwHY/SvVt1zuAD3w8l7vf7rpWIJEk
`protect END_PROTECTED
