`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsH8gOfyGFZuAWMy0VdXSUY5BX3Fgv/ced3YqHxjc8Y8tkr0zxYpXgflZcQd+iL7
kojuVq1ZFQSJKQfFaIUn7Tnh7ymhCFvxH6F6IZuAyD0u3aU5N0PhQX2xS5J1uB90
1Q+38XECrkasyinftpOGiVjqhUczP42l4BgmaBuI9sjjLO7a744iDzPyILRHv2IU
AS8Ku4+Jbf9965tFhdP2XFemdlsfWx8it5d0U6KewKrUqbM2+L0pFgx/HOlqsjKG
yBF5ZAtlz3ACDs4IxXnkPkvenal22XwOjkHvxUCMxn0WDf6HdwKo5xwK4tslRRUN
8aWBXuDdPxLldQ45qWOw23AMM4tU8Cyt8Dt5/GHyoYIFJIWI5R5p8H4pqrOWyEQi
c3N7DNXLSe8+NZvObnjYlcXu1nOrBel51s3/m2icPRnh7ejfSHX26yJnQroLkpI0
31NJpLdxmpSmClsXaqEt6Lp6OQ8vzz+jfWu2eOON4Vyf0yDi8Tm2GsRV8RvyJBwP
IDJACntF4r4mTgYSZHMj0XUKbNKaxq29WbfRF+yD3VxqC+TOZl/6RTAotHrtAS75
rCdJuG3mVKxe6MysDIQPry1vVxgDEJYKWq65ybv2NgCrbxfL1ufRKD44jX3iggf6
RXAaa7daB+llyULbeslPXcKbOBKf++JOetskKmek2g+9wj1eHL1UF1HQZB98m384
QBL7/IxboJP/V+70OK9Jhv/xot11mG2QOqrrdEMaW83pfcYvU1L2pIAUaEKvFtp6
qk7Jh0ZZTx5LX7oaDR1efPVEhDHh1O6/4MI0sEMTVXnKLo4zBlCFFo+/jT9K2CI7
/7lDHNpQkIOn8V3gEZnVm7ubmQBojwHUZxeODWz7AlSikrzXybzS7RCfMr0uqCbU
FVgh7JQyzNLF6Etm4ltIeI6kXZWI4Z29/rd7mI9AWZX8efJo81Eor2y9/I4sdxKx
DHWPiyD68T+AztGjY0GUcnFHoV7h0z7fu0MQp8p9YNUvxUxIpueOh6/825Nr62dS
OA6Eyya8zNh/ZU061FgbbWzEGZcZ7TYJlASTeRLzfWs1fNhUkwHuenZj/l6MjPdr
n59S05PNtcFqk0/RcsoTk+1ezhiTRlYiZLl7zZNvK0D07yNoShI3bCQ83u/juuxy
P5wUfr6YKQJvRoiBNdR10hFx8ZEZvjey9raoNBf5PWtDEabGao2pyigtOqbYJCXx
86pmRug89r4y5FCkpW9IOG2d1vpVJjEUy1ilQKu7IrM=
`protect END_PROTECTED
