`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBsG3WoFsUnewEbkjRTHQinxLkCn+F+KXI4qJ/pgeL1uf062VK2HbJVzr0dE3RoG
ncOgW0UxxCtcrYQYFjE/XN/L/EzJjmZyI5vM8X4xVqshSvV3/GrunxSNenMSXJqa
gNiJdTgUTPtpnm7f3STv1A04zqJ4yjo6xCRYYQ5I/+EE+G5dKkP7sHKGVXZJpT2o
ZYIufWGRAgR4KNhKnTh04ap50Vovb1nB9JFQkIdq6bJrEdZwAj3Iv6xsOogr8ItB
/4UqUBoP1E0tH8dS66xNRxdSlHZonIe4Wh7GjJ+UsTdfA+zEpFckfzrqqitTx6gz
iScvNFyKYQw7FHIPPiLl3fxEY77NmeAM96jHTwHUyUI=
`protect END_PROTECTED
