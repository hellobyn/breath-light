`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZGXmyFSCIBNp3JZewQTDFxjv4J9THTGsS4IPk1YZCXJOKO2NRJgfFp4XVDZRocfx
iP4oW988cnp0hfHX6VFD+EK0jlJX1+yo/tlVq95mtgsFaj5jfIPz/zDe/se3ix34
5RbWvRbga+Moc9aI4JQobJ0gYBRPuvgD8okcz3kSH9TcZlI9oeUSiwE2Y8Q6yZcY
1F9+rjk8uqdwNmAwcIT4aZKtDw5k5TqwQo/3ZwHUNWMx+X7+P1Muns37vXMQah/j
jzXqbcNdNbZO/LZbMnZEb+tttuiqJP4kGc3xFvsI2o4wVKl/wjfYziKCiI9WrBo1
ka6vjQWyGziIkRDpEEomOygwJpo7seffkls/YQi24QeymTTgyHcS1RUhqDduIWuT
l735qOCAt8j6JGQq9IFyTQBG8mS0TwPzrVcerx9DTm+zhiPR7dtBAzpGtea+SteV
pUeixeNhkmQ8/Ercbw22FejAfSHvThZiccBLid/wD34JNfEPIqeP8DoF7BVFPRSR
pVtAyDQjXQAQzSpDNX0W0fEkPSjiOEZpWNGeFKRugktVT5RBlO6tbWB0UwW85F1C
7TwPFB6yMSXIS3JEI6ZXKiKL20hyUAnr8iRYfqpdOiIOq4Ih2qGovsuAjVeiKA+6
63ivGHN1wzSmEt/Ag0V+D4Mlr6MlO+KGlWpbIvNheXGAHUNKgYePRl3QB7anxqNL
XjFvRHo9PCqmkfwwPEEVp57HOjZbXRWuFyuLd69P03LLeGn5Wi07bp+9eS6mDmAQ
ViRgEM5cM8inku52PGkSEKqfAiMgxdVdieNzV44cZ42fslILxbX17ldwHbhrGGRz
S1hAN7dEEqSfLPVrTS7adba+6EOFAZI3HdmHKQ9TshxDwYwRI7csSsvtRqdUCZg/
2dSynLZx3YUOqF7JkPlOw/UVMRKVx2zocJCin6ibSwXx1t7I5PZ8zYO8/nYdzW5X
NqysCuVgMgKZ1B434Qyg/fUnfSde3M0XzRa9uB/vnzi9ygoYXoJAk+4o7NM4tpHv
jIe9B0TFd8iB+uIieNRD9UjhsMmbFgBuOhWCrjSnpuzaM5gk+VEA217q7yrZnzYS
pGximhrudgomBObRXm/TcF8pC7raIx/9rGzrWxsxd+z3Nv0/Tbv7f/l82Y5u+s2B
b3aaEDPqxL43yuoQo4OGDjZyiKrIyPIQ32H8nh8DqAGtUtd9B6J65/2egLRnmPmZ
86ZIxt5k+8WTWAByA9b/3tKfWASPJfXfX7Mr9Zm9KVsAb8wkMj+egRreJO0kOzZP
np9kfpy+0ks2S8lhlE5Ni05cOuUN5rGrMdM5AZPTLooXVgKiEcA0w49eZXQoLtGB
UjxSdxZr5FLUF2+fwIKxQ2kkibopSMMMsEua/tlLLYKlB3mH1j5qM/JeQu5O9tiq
Z4kBhwd2KPltKFDmqVoBMRatNpcdagPo7EzLdSUXdV1BW/kxddR1XgAUV1oHOnrJ
hZ49sQsB6fpr3qicVTNeTPAItCNoG30NU6TpPJ+fr8o0PrM3CkQlMZ1Bd941OvVo
FOSa4JJ/oGjGzRzjJCOrPw==
`protect END_PROTECTED
