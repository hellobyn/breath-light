`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hY5ndQZRcqz8/g+TFyj8fUw0VD4XbdF9RrpxZEJW7Hdlx2G+n6GagZ0BCnuysLbu
e7NSmCb6+xUBhsrqatSA49CdeZocBGY7iJeBHqMNoYxV1fi40S51ryZSOrdIN+Xv
N/sTHLlokmVgemkZTf99YHk7Szhk+lGTtgV+T9zmgaiheu6PLDjlqDRk3N3VlhI2
JXeamuQJrTOT6cKp+N4Gmce8LQ5b22nl/ObSHFmvQNoJFrSnUnKM9x8x0QFrTfiE
eK6dAkTToRtfOGCzC0bUue9At0TjDklJ86Zl5zXNEoo9xSpZ3YRFNhJk6WDp8B35
I18slXIfrDOZfa5L+swbvd0kBbP/BYr8YpSS/P02JKhF4bN1vRZi1LBP4AqTgRfO
VgeBMpbyjoAtvxRwtsdCPU/n599BOpyxDf8UV4e0+fVJrldTUqSM5uagIHBx7X2A
a2xr6oQW9+YYit178Qk5ycOn110zFNptqjQ+8e0mPrstctEQXsAoKs7kV3NCzGpO
9T+HhCaQtTrz/tlvZ3Fes5MkAAanUkIM5qUORCMfMDbNkxZ4PEEGk0FdRvK5AQMQ
cN3uHFir1RpvDlX7Q1cRjuZX/6iqT6Bsj50RBEXiK5BUADIwRCQzZjoTLcBN/tfg
A321OIbJkPlQ3NdLb7FIs2WWr6c+nIEXlwg1BhasRjhSo+LVHVnmpvn87MvR2cB7
ge9J0/R41wXN87QuOW42d0QLKMacEORR08VDgheNUWCzXw7AUDHNlZtC1Bnb0KgX
tFwvc8ksXOkhh9UCikurLf1LiozqTruSYbGXKoc83NTJ2uj/qyFDzXngmvaguasU
WztPQ2cCneLv2IX5geuyjLyzgkuZLB95ji0EYhmp3c8C7aVp2SUnZmiDZaREwY0s
hDJJPMrtFkxuFxGSH++T2xRR/ScaH92zFaiAB2BW0gtqy6kO6/gk1xQsnHKffam4
bZmpsx8FeJ51vBlgMUsIOxdEMcbi/m+GMBx4SBtBCHyd4iisYoiiJ++JkLligoj9
ok79McF0Q8Db/9JXyve/QxvSGdL+syveMaVkOkan4XFOuYZ5dEcS4tkcQPO63sAF
1WpOW4O0LIeM48ifCg+sEXJtKfgrCN/BPGU3K+gVUUxcYMXRf3IPpJXfnRV2E7Ui
IyEHsYrs75+Aihy24D6CnwfdkQ68WhRxJ2Xoj7HpBhogX48zsWLnUWWDu9n3Q51Q
5aN2aqUcZaCltjJJ+cYXLry8Rs7Q3Nnx3pZsdcZpZhCmk31mjGGv/DSDYE4ZpFTB
hayY3Cf9dQOegzZBa7O2NnJGKviVNacv+ok4pa1GkC5gjcAhs0eKGkD0jnfy8kLT
UchLjnHfYvHqzfLewY8xLmt56AAuC+7dQiLh1uQ/qYJbyoK5lei96JAFmazmepca
6QX4JWKTbLq+No3ZCpZsbLRAC2m35IkLDtOUsKh4sNDuUgavXvZYxgmldIQ5ryg8
lZX7zoDgNe8Guc8JztW+o7rMc2KQMkJiFvWOgQMG+so0UhxDyn9GqLm+ijHH+C/s
MhWqumMAooThertZDU8na9PYSTeVqfqzIJaNdNPMZwa2m0d6zXm7rabp3bDlbTgz
+OGYtDOQUitvoaNtOmz+gY7vr++BPl469b8IS0R4SvFWWtcnqilJCwO8PXQ12+WH
flROhI4iza3eCUBk6+flV3UM6y6mnug9Ar8DUHyRJ0g9gaBM7dECGz0vdbveMkV5
t4gv6lRav6BC73F3B98Jcxa2aSE8rebl3A/xHJ8mAbX5pL6nqK/8hb2p7HAY+cjW
uiNI2mz6+IjzrRTh2HiQj6/BZ9S/PN49tszEinqiwXAXZvh/25NowhLgap5K6Ri6
vHqMyT7BfzjENprRv2u4ZuGyoqqIRoUxuKrTVp0ir12EIqK11ooyIboPBNKA3RYv
908ns/SUmgMQz+5UFcMUDroUkhtGJZ380EnRzjOGbTEVl+/uIRy/gqvSxR1p+E2x
IZKfFaY0JjJSkd3ew9tinM5DIjW8maP9v/+q4zGq9QhUeQZknBE/9ji8iY2TKowr
i9Dn1WX10GgW9cw65NqoT6/hmJ6RkKYwpUSnAR9FTP/Bth24Bp2e2pREU81zFeIR
RsAVy/DsKWPTvjwE7OlzC+sMCm1cmQrEJf4F3KHCKBYN5C9CdteduXFBm8t4IJyP
3ROn2D2Uj/FfTzNbJg82DBiBAd53TldFAfg/gclXZD6XRSD+xuv5RnK1xT94e/hr
CIaFnJ+vDNtU9dc/D2e/f7HAjssm5YPc/4u8ugprPSVH9g2MfSt0rA+vbNw9U+nz
0gAxXPZpCSjfQB2Gk5Ii7IQZblOBMB7Tj3Rn6yGWhDGaVdGLNTlmv7lwSLMK8rmO
gLUDCIHdsefvgq3OSHAM4cW66Xq0Hg1VKzKQQ+TQVpYtCNSDcxqPmGfHQnwS9k20
/PA4fjo0K3HQyahc3Muh2JdDYTmcvkBURbwfI9Ep6mQVqp5nKbNsm5FafY6lANv/
+3ySB18K8zZIKijJVAPqzPzTZ4tZgWyJ52CJaDDAP6CYXYQhS6nGf+F2WPygs/w1
KXbvpEixcvSmJPTlyqVFcdsyLs/d72s/sGro357wGX7m9g2A/QuzUINCIt17tO61
QdtNMX/3UVWPnkoNWDxD6ldOVhuQiYJUA3cHMMTq+wbfbogi8xdW5gpxV0I7KCBt
tAYY4te9Ak1LLbRU0nSPt/3p7Ez5iMg6qe54weyTcnSeMfb+fgk3Q+ME80HPL+4B
5v04g0P4WahymCMo3yMF9x6DIvB4Y2jOKss88CRiY+peZOiUeU5VfPNQi6Q81D6s
kbd+zgtJ6DitgjBlrIU+UTkb3NSk2JbB0HJ1NNqfw0iilAHtRYXG0pVxXkpXb2PS
gATB/VlxmCKV1/ZeVi70xrf3eIKh+kWZwTr09fNaw5pwvo4nkxoDtFux7hJ4wV4Z
WoHgHsc1eV7+vqnxmaHQushumltdSHOCASBl2IMspXelLc0S+F2Sz+FeprbIVRJU
4h0FTMKlTGSGEMATwVJRCico4oGYCX2paAmPXPxIynY1AK1lxZlsBY3gcvmF722z
0LCA4CFKjjsvxFSssVdoJS8i1a+9KjmaBEa6JciDFOOwdTZZLkplfbpZBQsXmelQ
FwtRuLEOkNygCDVZVc3725QcNR5xOSvIsdpsmKzbl2pTw3sjMsdi6YXEqMX0i5vK
KXGIUgKshPx95r9Otp+5SW9YNpBUkVwngNfHucK42WKD880iO78q0gzHY1C9PQHi
ZI7eBvm6TMop3G7V6jmVwQUO45dY7+QbEL7c9gQFqVuzsawGGI2oIlymcjC+/R8+
U85hrxmP8qBm+4ngk73mpx3CMz7WhqAHF8JYoT4LpryulJH3cGmanu8CQn9Lw7Sz
Zj7sept8KjP9+YnYMw7x7YKNuUP9DY0Fo13O3yCNcoLGiJP2t0gG/vuqUyHNnEO+
Ob6g5XdTNYXdJzWyGcNEj9FoYGX4SUyYNXGCDfDCtIGM4Xp7i3SdN2oORBHNtJ2s
xvRY56B8PqaqBMVKkyC0TW5tBT++iH7lUZ62OXsLuly8U58NsEcZfmCNaWwoBLpF
hjPWWQ0ZDv44kIge5t340fU6kXpQ0PkqJcoh7LzMD5aOWrhd8dmzSDELAqfGThwz
E/6IixJlhP12+nnHC3LCDK5lCHWgwnmq8JNfstOxsK0gkdhn0tPeq7sDmH4YwLKb
s4x6Ihh/F/RQIZQOeLMQQZkA9GzE0Bksp22ZcNwpnTgTadalnILj5wS3bw+KVhsL
re5xQA5/FPN7Si1Ve4LyW3VNmxst+3Na9VtqIvNuGhVPYzC41kpnUCOjHSxNAi8O
COoxh1nk8wutphdJLdkEj6poD7pj812dj5Wq5QhDlI6M1vpQyVGT8B+voGh2374H
drZDzIdBcxJNheQwl5cu2uBN1AS+pYj7MjbfVEVMJHURU4EUy4t0cLzPdfTGw74D
dRMSceffJQbDTGeX59k8llujWRskySpsz2yQsWPvixfQgA4HVPl1BvRKi1fv4eDq
OoIBFcKA08CtwSpa+/UW7i0BeHrKkac8RXsS4twekx10mjQZGuhiaN8gvRmuKEfo
kLyxgPXXWv+5yLJQORnOLXqBjb37d/4eOCXBF4zYmZ/DtF98XCRjm8GBzTNDPygD
xs04aRIhcJxR77sH2vCmmrKBRmTZosRpgQgd8P5+vnCy6f6V7Onn+UwryCeXkmE1
6QPHY2H/upXVX9h/pPXwvnCEudgjwAdz1yqzU/HpTl71DAF4cRRDB/9tX74FQatc
+N+B7Eg4cN8ZE06IpIkNvfw3TFi5hK8GT/6Ce6FSab3BcnWFXIC62R5A2UABlarC
gry6c5S1OXZKeud197ANoE9TsNoXJUnaTZExUR7hzsBI6OgHWj8/f8g/Qsqe7TsP
jECPV7Aq5IxusltLXrAL7U08JhQSeREVfmz5Xz7Tx8cfAEbKJ11tkOzIZ2zLwwRi
e55gMUXV7IRX5hsAT35D1uIIK2AZ6AWaGmg6LXEHSwg22IkP8HLXVCb6weCf/2e5
S5icTs/8zaMg9td3Z3reqJe6SQ7Ky6++tIZdvVdC+ocLgrgHhUZgLCvm5YSprGgn
f1QNt4m/dHLOhA3HH7gLzzZiMJnnjmS8zWilqu/l7fjYfjjdBUT64JGqpcWiF3Za
UxaQHdSFOSbr7U5c0UmrDjMuVu6CpSYGV/iA3kVFnYjs2NTDmNnlSOi3lv12lmBU
wGrShgDA9aZkrJ8P3Pg0pYn5HCrDtqvdNtE3jibqUxFWF8m0VCvOVJtIchI11tFw
aZFmow99RTeC+eeL2fHn84ee/04iGAGlmX73vF+uEFv/+/NtrMOZGKyNFQGeqTem
7Ixse3LZ+XEhRCFFpV3PrSGBp37pnpbmm56uxVk4usKSglloVcMLo+6nDXabAWxZ
nkeTC2KeHb88zNl2BS8k7NjUj17FopXKnHC+WbghuN4UfdDSYmSF0a60qLBPAx1u
XNhbY012H/HdCdisY1qpGXL4iF9ZIa7eilNZS1ohfKc2+/0/alPPhQbmZ/aY/Hfn
CQyIwavKydb9vBW/4kV2sJctdyklilmEaPtCd1pHX9STogRNy73cKkh667QefmYp
/uYH5RTcmfHH1L6HsynUGTRauFHTvhihEM7N1VBRgbs52oLrw6K4KPvQNk20OQXw
397W74jUbwHnsiM897BXVgwkKDEhYKhgLhqlq4XOMa3Lsu9lDpDrOZfc3kJ1996Z
TUp7GIRG5BYvGREd6LvBtHJTcc0V7mb4tJBkYiKpMgXdw2/ikKDyo5FOWqpDbNxk
/s3O8rJbxsNk4UtkUKeHJ6xjbe9k4F5E8Zhzdfa14vyEC+a97tDhWSnxT9auF7Sr
E3c8BiQ5z+DiBtP8X7QEx3XNzXQtTH+eDITYRzP0BasjK4U4d8Ir8tVNJu8E83vZ
kNxf263fk7tP6rtsJUaA1OuZc7D0mEbS1fVEd2AseV+p+5xy7KW+Mnm42JZjqdSc
y6i5YUr5YEGrZ/kkdixJHJaYSfGP7VAoGxhLPxqkmsMEbIjnFVVYQdnkN8yE+W5d
xbWVEluwu5MaP62zZG2/vo9kwO01MPnpjf58HZ2Sc/Urx6Sbz0fEqWt1qEeX5Spr
/idM2rHiuH+F/x5YlljnpXjNZtyoVZ9BF2M9DRq1X7Uk3IYn4nvql1QwTfAIwMDl
4mApaoPD9WhdyoUvVX4keruaeUKwaji3McUU9k+bL/jyQFtfc4K7h1dgBX3aC6yt
I0Fq9o9zbE/LY4udrUSDIEnlroPZL7TB8c/5MUB5mTe+t6JpdUsMEn3d/uQfA7YO
Qu58XH11VDhgijnvdPr7h131A25mXtUkgOVHbzqB/CsobzYbMq7WJH5A+S1Sw5y1
+dRWOK2dXNWXQq/ofF2y9WhmsQ7mw+9XDm8ARLHX34OkIe0nIzrHj6cJpchsCeVC
mXG7jvVxOptTmja0a8+yz4h3dlvD+vvv8zg1SQ1KGiu1/8g5Spvp+jMGBRgn8Lk1
mj3aNnuIo1tiF4if54fT7jA7mAg+Sew4r6ZXgbgBeGBYbFENMztKizx3JWNNgXkP
B/QgpuLlZx+697bb3CSttIubSB6W54gixuXD6u6c+1Exqq1oIYrHhZmQR3l09kCP
72rRJL02SGjvmylHeoj/TIEgY3TPBPB2OvLSGO0oI6XZw950VD5GXNQL95vkkYFD
xDk23C0MXGOnVGeTWW6bKlFhM4YDvcdUBdrFtzt7029sLgDESNBMF7I5aKte4h12
ZxOwq6M+YrF5sMsh3TfeJmuSp9e3LosDHSPorY8t4VulC3JUCF4mM/3mLNUMa2OG
RRn/wxXzTk3yZDHH791JrgwzzHgcjk4ZAr6d9O0TKGpJgKPOEuY9u5Yuc5XJ6QFb
KUDP5pbIuhDdcnc6s+JRIDAb+B4e9/OcNSoyiB4OMCIfqR/lfzPmUihGc1P8DKO9
mXbk8MDco8Ooy4R/MDDsAKQCG6nnn0YcL0/W6L860i13c41NMMZSLZIH1U349Cmj
M/xiqqKfZ1klpNxFoFSNTwMoHXJ5u37tBAx+QRPJZIH1FDFHbjQuMbp9B2q5f6y9
9reI2K8WGNN7GbspjGYKU2Bcu+fAylOHErocCMU4BSdu/PrAf56yCkZG9D4kpz/4
ybLDJCjel4H88zWqHx5PWxZyETonw/OKjhE1rR3tU8XSluLycKARw387THJirYvc
3wFrsQxzvYX2tB2o0bCFSYbcFMtDcOrU7g5aYNvwgZUFZVopVGMMdZRPR5PMxIAj
nY7gwR2Qxkt0SQH5uotpPn5LTrNHA2GuiMoolqvDymeAOQqM206tn9nOsD7So2h/
3foK3FLkYEmdPCQZb3E4xpPdfMYZk0iUodj7YJzTRIBYdPPnkF1tHgn8CTBZAhUz
LabZKi0FDsD1+iFpR8jC+aizIgypNtbShOkrrLca5poEQJ+3FTuWRGQcAB2idT4H
7+cu9foEQLZ57YBhPkPds2JknJxj79SnBFKWVDXVKmd5B5c8bVFd7rRID1/cYgGW
nnnVft4tOOmvu/j2krtPTVq17gyw/sNYqKVZcyF7luuTBdN7YYxcPUTCeUcfAMEG
WjLb0AqolZTG+H5/D5JdBh3Gx85XnlFXK78a893BzzD/SbI5zvNbbMz3OBZpoEeu
wWjpe+vckkW1wZZWpEByWeDmwZtiD+GMm8KcYxo5qNAGmc1AJobMOMwAbvRzs4TI
du6tJF8/YucbU9No5s81Lf7GuI1EHMgc+4iYqT59+LK/CXxDd/1xYWTXhWATS6k3
H2KjxvWIYp3Y9NSE5ZE7pjnjXZvSAYzQvCES08W1eNYO/hIvFAG3sulv63qwKuLd
E4mQnr+Yj3ZBiN4jzlQu1H2hraWfyMjZL7jgN1e5PuoOxmCpkMYESZik/ku3oUO/
guzhi8CRhqrHIFGkuaLXDzcKx4aN7Ye0JAmA4oWh9QQV/i+M9qnU89M4MoocE1U+
SFZkpwcMBT0cJkcwPeb0gkizuOPQhXoGwt2bsd/ltXDdeekswFHhqJ/Gq9OhmzoG
7XD53V8iSU6HqNQPEcDarxqKJ38dhS9Oy02qhhk9HpA+yxlpoikGlvUFar1gPr6K
TgPawBlZinwd6IvBCxLZQCN4DOzhMagS9MLHHm94J37z1zDrH8P6RaRAu0hIDC1G
UKZPS2WtWQyuiAWYKGcudqflZDwjeT5DZO8NIXivluCdCPQNl9xXWm68pf4+qVA3
SUFdVLRGQKD5Nl0TN9DWnw==
`protect END_PROTECTED
