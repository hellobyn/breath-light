`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7P4yJvK8iNi+WNBKw7Qzh07q2Pq6sEmLyIvIKNPA8VhR2QTNi6dt6ZRpex6NrX5
aLh40EjFiwxZjMoy6Fw5vgi9pb3Ll6sKQxZYr35JsKe/t9gn7uW5lsqMUx3IIUx4
wLJVAq5Lq9gvek8Bn/b9bSNKLTF0MwdvvUyO46B4LCS5V0BiFASwYWTXDN/MQwzO
MvL8OuDkWFLfxT+akmpDxHQkKabBcQyweQTkWIaoTROa4PiQ73G1FDcoD9nImnKl
ttYQfWt/vKAwzVh2ZfVTFxkbAsiqkIWd2yDgipXKebtmGAb4pXu2uNGjsK2szU3p
4ogaCkxRIF+TjEl7dK0RIukMbkj4Un5+85Cd2HGJBzJSqzagbQi/REGB2Osadqzg
lD/1VEFyjWYQvXC3YPnm1KTrjmyAL/n27mBfTi9utw6K0mF7Dh6cmjkwSxviGHDF
5ciWpoASRjsY2NBT5rgYRYjuGn9jz3IurFe4shej6DFZsLIhsJlSl1O6cO+Rhaf0
hIsfyv09X3p/htPVgGvVS+KFaOzJyDVj9YAVrNy7KF63NHjzkXgbu45GCFi/kmKc
bpw47VL/w6oann1Y1r7EanGUcgfLOnEfRAPk0GHOlBmaP8oWV3YjG+pusgCmDpHJ
zfktOl+4IIrZTVDOOfub6a3pdHTAbgFSNUETtnmmcVa25ecMu3sKIO9Cq0fwrA4P
5+aEyItJ87/R2CbEWO0unpPhsZxUvqanW7fBES7vq2YpMvyZugoN9TS9N67vBj9T
xX3z72Hu2JGfgpx1iVaIZQ==
`protect END_PROTECTED
