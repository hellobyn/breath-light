`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nVamm85weetsCYqQly9tJxwlu8PVJqoOCbGkowjLNqfKZAH2jf3nlyIpRXPvrcW
HuSxq9o8F+JoGGQeQ1r86AFHKJaMVJaOAQWs+ngEXjjcTU94lhsH5mg/VNSRz46t
1GDE3DPUtdMKOFLKOfdsbqWbawnqUJjUzHHzWfDC306zeFzW8M2sz9QjFtgXwZDM
stJ1lWmjz4w+pz+2bH3zGiCys5/xAsQYteT/Zlo2k9ru50Rf+g+0OZM6+owyaRqA
6SFVF3a5U0Lj3+4FEu/0aLEIzD7ooc9VQ1BMdEgrhkuts4luz4rNA3rKsBnDm0oV
h0efO9KYjQ0QIsV9D0qSckLK1k5o5qmZASElDjoMhVhwUy1na6eOAeVphUGRZuDL
uC2ZOUIhdBwq3YUiccv7fmBveCTgPv3PuWTGxJCGGuvI8pXKVMML3aZrS4ICn3gZ
S4jRd3Y5vfbD9MKE3tng6UpURXh9TS8NZ2M52/gVMr5qoDF3UybFQZK4QCShwraU
vdx22lS/MmVbitP8JrhRF1/JG+B4KZIYhTN979n+ffUoXeOPMVBGpdiG1O1vzs6a
UqBrc1SWvPZ3ml9A30+F8GEmeHN7BNrwndy+UfajxUdtU7Z73UY8xsCAPyh9tLcG
0W3RHsdPkC37tQZXS9Au8zJEi79z+nPo9GlskLUTSnZBBlBWYtRwf2GqyYtcgv54
XczKVhg3Es29bRqMT7bM/qt08yWW4kGFmk0mLr3J1wJkWwGi3ErsZQ0ljslu8dyl
NuExRXn3+waR3fOFU52nWVjwH2pqH8FR9HKDWKGC6LoNVR96Ajr6qQ4NRpztchDx
QVDFJNxghlRx8j7AGN3cO7feIwVbWJXHBI9kawXyECPfAHwpKfxdh0K1WEJWGjnK
Ro4IrniY8OUHq+RQfW1t7JZTzFRgB02nM4U8hEBr1ZZFQLV3aHPVmeRCiHnJMqO+
B2kEnyj9stKjwdApyw8Tm8OmIQqiWhm0o2tc/3/blBAUjJjZV2oYWbAVeJJeV+U5
dgFAiUfOxJBNuihu/NMXel8hQ1PmFBErfyyMOMA10Arw3WjnLGuqO0ONIFJGGaBb
tIHSdQ8ho0alaA9fekq9C0+h1fFAnTPXRDRz09TaZtJ4ShCdM1iIo8rdIvSUgKke
5GlzoX+rIKbfqnQux5iwo9uri020nli0YTuMvMA9OXEWnDo6WZv9BLcm/Sf+bVaB
+nm/6mWJ6q3L93ac17+4NLeTSUub8dLrWwxf+9WNdGzE8c75HajnJMk/RNNsXXBy
RfkNzV/yQIGwoypEbisZ3r3GZh9QQTsYo1B5Ar+0IHFBB14jeUTtvFyrCrR4/OBM
2562FgAI7dILwHsdGbRjO8728TDxBdvqqOJA82k8AOjb07PgBbu6gtJGC/BH7Ge3
5ha1MZFw+i/gpW8oTCeL4r8UgyDs/sWSBNCzQaEM1yrFVSqdVMT2P9mPycVPTSHz
yhNosCyvJZyaV1F244wDihm29PmnvsLHDgstEW9Ay90=
`protect END_PROTECTED
