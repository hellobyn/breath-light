`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jnm+dbf8icWxGG9bD7VggCntzKOvA2lhVX4mYPOtipS2dURdFUwwnxor51Pueho1
4L7x1xrXkDxD/B0ttt0EaY8ZP6POkl1ylPtp2i+KlORJamMZhH7RYeOIOCeGjyEm
C6gml2TM8xfPNZrXa1HqtsXJH92/kALL5fuAva+HGLNXUK6II+jyJ6xYuMccgVID
Q6K0RoahdFrr2rc641tZWqAj/yDL3mLpQxCHMyor1FHnhBAjQXqls8Rg1NII1jWb
sru4KDoHU/LiM/3HfZ7LiDUAMJ5WHRa0KJ0LkbeZKbX5YvmlPda/3Hw5biKieBcF
7GBwSYu7QBXoGkjHCacfCJl7857P+LWsvdp9d2oI+07vLudtkKuzkVKQEvkabFgO
Xe0UC8za6eFPzdCVCkeTc6C2rWSEDSJYgM2WKHmBcKAks2o8hL2loZMe/qOSJ6Ca
PoCF53+s01PW5AmQ+mQS8DS8z3CRgcXppkld0b2TPA0D1u1Q2nj6B8xgIrv2mgRI
B5acE0BvJ1BlMy1q4A9Mlvvh0MXsyeKFNHvfzfqxzN7RVa2wJfxpuRBB4N3h8URC
9R9VBBFC9BgJwsd+4iBQF5AtRuUHU2PfamIUns5i9ITELkV0UcxEjqNFuFjkPKWi
49vNluM2UIsg/5b6tJwB4pLX0dMNBNO0bWAv6qbTArdXHOBz3Qk269PgW9WmIlBO
2VIq3YmklegW/VMP1ztwpzV35G7YONqPcvuxNfk+WNeSAGl86StdpDg2zbDDTLOz
LaAadG/AD2XLVTm25qKuCa6fLSfDKQzwlOXmnVugnMqEL9oboshLnMkoiX6jJjRH
KaTQ9zsjXD8fi7PxnMywnEHStyxCgNiL/JOKe/wR7ru4Irzmy2ouVCwnV57CkFa7
lxlu8Zcn8459xcVzTo4MoeXmTayoJMbaSGfJ4jhAD9XbKtkrfWAo//5/PWl6Sj8j
SXFYngM6Ctg8aiodv3U0br1CyE+5jZ0kavm/WotDzy8bikhl/ezk/ADSv9NXn+5O
B6Cpmb3acdCdSwJnClT9yWeW1Wc7bnwo/0VpLZuqFIBeOQjlk/e/XZr0jtyX8A8o
xw1kENSh/R19+h9tT0ORtX/Lc7S1Z6WVj8qRHTbipm/twWzG4Fwf+akpLTndN4sR
qZNWxwNddGYH1dX2fopir1bm2yzOw6Ssoj5OdPtVpgojRg/WA76HBrneAI2GnuyI
hpgSMvDfxz/fE2zX9uM73nLjsD3SqELJEQqmPc9J/2ocyH0vZfBkSFQfsC842B4G
BLEVoko/LnQZK5h36HaVJJTnN+k+W8t2JYyXBEkrZSLYsYKIyUBKQtsrxAYqM2OR
Kui33we/h4GEvQNa4b6P2/fiPTAzD9EbgV0B7+yBl5RE0jNQw5am/aLHUyqLSekc
8JnBs4+muynsnRckW0Fo6e+idk5xyy44+WvN6RFeHaxQ9d5QuQPW5a+jkxsZ/Zrt
tzZmbrZnynawSXiDdbd4FaRZRzmlFYyMOarJzKsIsLfHQ+S8bg2pos939TlrbOp6
Z3Vtbem9HLHRM1YrJOblu+v2A2Z0QAFu42hOYOkHgxwghaXDeaJg19qoAUtpXIVv
vvPOAwNddlAToodKFo+qQtQvQTYyGfPD7eI6cMgvE9DXf2NcAqKD93Mh8LheS5y0
rQLD9WSN87tn3b3oYb6HgO9Ph242JLV7BWKQ0zRK2Ty8rLLHGo8eu/CD0zofXPUS
D3b9FvoQhr5ClP+SMWC7JOvwEIHmRbfvA9UEXONRFCy+a1C7azCiw9bKdEPgOORF
sQhq9u9c2Zvso041DuPlv/WxpE2YjJIRlCSCBbZZgknTY5w0kQBttVkeT7ofXdyr
T7e2V4u3MhC1DOBxOBT1KVHSBjdifwpVkVjqHoLbzpvnAw3h+6xj0PO8UDnv6+bH
QLYiC6SNj+WDKLFmRnmI6qPNcsg60QqXSbPztpWNjNspj2IoL00yjFdiUsJnT/pb
/rZwbzAV+X5/Po/z1p8EH+c24mGZi/TaspIrIKT8/ketazc585spbNHUCBWiY8+L
pgZ4VhtWPCuOq1oDia7OD3gZ6n4tWLpHlKbEXwvQIsL1EJIJqV+jc/TAsv1HXm1J
XS9k9zO+SLe/jDf4LZm9vlNhBewGrsz4ianT14Mjhu4coBkq+ZsSy7+E3SxBvzWi
WR0PaXLYGdsH1F+46JwL1dLKA4uUN1ThLSVwEouQl9jPMcJqWsRlPEGy5Zum7eRr
bZIBgJzYEduH9+mg4dYEofLP1zmwqKifWpTfSlPW7vg=
`protect END_PROTECTED
