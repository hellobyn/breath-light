`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvd1scWkURJuihwFEOpNTruCsQkrTK4+hme54Tji7BITslLoWdyf14IrVxkN3wdx
uVVsPxlOH0Kha58rviwwLkltlUcg9eR0kuqUOttLlPxwW1VrOY+s/Xe9eeyIoWt8
A98Tt6HV0SFsx7pAoYpXT/2AVh9aO1pHZy4zR5o+zuCQMpxfOOlaxs4mlYjCeGI6
ygPFRTeoh35YFAieedG8XU03mnSAJlwBq6D+8ZGzRhlPhODjbj3Spff67WDcKwFL
Fa5kMl8kbss79IkLnsdnx+B/FH00aRnwMqSN+RNud3cBGAKfeFjiG8q/bYy2buLO
Flo8YUojS573fwqvSwWbfRoABVCy43l6f1Og67sIH3mSAf1brnDpohM2qg4wDaUi
fSL/bdYUqu4hHRK/ia9pzejCcKlgN/7OkUoz/ioj8DAfzXjjfnhS7IZGXKRS4Esh
uVCRJMKVq6h/zbVYCemv3DDTrTfblBeVzsBSsvwg3iIzfJRaHy54XZ1A4n8MIg1K
62xFDoXxdaNznNpUjdVopZQPqUTpOD51ounGU5a/w4ZqyUWfvOE9Wm/gspP7eWM7
JXhEPbDU/2On+uBwyWGujOnTq6AHp47+fSMdo4Onl+7sj4TavxdgD+3pk/AlHo+t
XHlWBSPXvUJElM8nmlbQGdykJ+HxEdvrdDfPkwnVfFSZbjVz5U1eoSmhKo/LoKek
grQppKGd3FHMIFqGxrGpef3CkVtOjKR4J5t31jMPr+6tBPrhoOra+Gi2eGQHJ4/O
wYDYfyxDCbG4QuSUge8p6uVX9Tp7Wa2K/Xy3tjUC2JhvV6/b5LZe9gCP1HNhyvyz
IaJBwKG+gEHxVuQxRqAouoC3FIDlNqvz3URLBkjgUzcLQP4C0bOjpnBuZcYtWDED
nDpkZ/upnj3TWUyNsOqda8em2q2TTZH778LeEmuGVFpJbGpQXl2VFgfeocu4Qm2Z
xf3gMYklZroiuIsIWvhV0GuhtG+RNAKFk3weBcpPcSRqa/413nijGa8RY4ZX9YrF
UF9l2X1R3O2rEQ6E0YD36Fl0R/XLRk4M1ptYkOG9Lko1JPFx1JFoc6IHdcDOKZHF
TjLoYRxijK8MFjXZb9EActd3InKj0JzUpkPdOh4Zqo1DTKH5qyrAcAhzlgb9QdA4
M5maQpHURbhGmnl6Nb2B2PCDXD/5Bb4uRmTKXEGRznqWWom3UaEseSQXWPc205eN
sOigeG0d4N49xz8X+FMKpbl+On0aTnzNI3Hh4xL4i8tk+iHVnCC/vCl9w1vKpxTR
`protect END_PROTECTED
