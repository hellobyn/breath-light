`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXmOnG8LC21H0R2tOZxFLBg80srfIsxoWsEqpMTZx5yIse0m2tzBzKRO2zdhDIYy
xEi3fkOZrpkZSZLpxcpENOul0eGw9fjWTnyv73LY5ZtpCGQEAKrk4o1227QoUusD
WwGiwvOyfdyGMNcDnAmlENJwv+kOc+tZCs+52DpHsy8v/GTVWEZrSBdwyKoeXpH0
QQUs8ootaOqgBjaYTdocdMvUv9Cp3qFzbmPgrOwvNO7Uge+SX+lm0KaCeY8JLOnW
i+9uNm8TM9IoW/hml51U+riiWy/zgnmCiZUWLKlP8eH64CID9G7Ffp+4sP8UpT1C
Ylh+jEYulcoIIQnnS71MBECMkVw1s1J/mvZayOUGkxgnT7qj4tMJLM1xtCS4IVOY
31BTV19JIqeCz39TlmBReBTYM38hi46ee3w/f0rgnVx5F7ahprBzuVnXXkIdpu0Q
OXWOxP4swZwAUTlzJJnq75GAnQSLY2vxKk5kNMObxvwe1D2UcryuJEA3h8q41jUq
RWRrwQPc5dQIIZWXNt1en3f17ak0TGvkkRM40qOGsSV4BNJfbn+/Zth0qGovodAV
Dj0ApKp0uGStw/kbW4PLN3q0lhrsmUpsGyNOvHKZUQBa+Vd2UNW+n0ybTx7+j2gC
u4dXli+PNbi3YZfHzfeMjotBnvlYjHR4UepBBnb2OEyRJgETjcYg5iDUAGhLBdE3
ZLnJud8rexegSt5R1CrmnjHiATMXVglpSQX8MKNiY8VWDTgg1a0FlYqc3sJEpI5L
GvoYNKjYk6vZ0lGNqNxPUw==
`protect END_PROTECTED
