`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OT3QqatkUkiFfZJMf9azgN3/yrl2ox+bnn1/miGTyo6v+5HSwGHW67P9/B2X/Hi2
y25pik1yfknhn5oZURMyqYcusFhzDd8j6yrwfJIHEPjtVzWO8MBp7z+9u9cH8xEv
PRFX1/ZkmiSCfOJ9KBAMCjgtD0wG494t9gmotUEOU8DondMfUbPrh75gFPGyYCoD
FI4NdxdXelSOEvIzIDGcLZWkil5NFtwO2Jv16Itir0kpHAORU58hpwhCkpKuvbNJ
mAShDjPAkulx0ok/qH+kWoT8Z4SzfBhGugrRrBCbOD0asR6yAhqfiLVQo/oXo547
N7Wu4eYf2d8IKjgR4itWVnLwCS7uAAoZ8/UD7nQstWlQyF5gk4PxwdTO5DyCI/yP
1PcJMh17kTM7iwLMv9wEjY3QLlUKBn04Ub1mv6/jPXWITHP6vK4eJpS0KkykDowN
FXYHldvQP4ifMYOEtpBUAApSM+kQQmocL9QU1zfCqcuQwoAJVEeb/xx0C3wFL3gE
aJLh4KijxlrY+W5sbmKtrT47PGfsatojP6xEsxXntjsKcWfdZfyJzHiIKvYpSCnK
VKQgXbR5DTfmzNHGP/EcMbziwrpXy7bzPZJ4l6RvHQkbbzUZuZG1Sz2cY0HrXSi0
MHKu3tBhaBoZhW4ox+7Xu0pjpry3BxBRKJp3JBoWoPBRx7ZsiaFO+DLQqhywnp5x
se38pYnPXDrrwNptgJ/BhChxM5RRWqEYCSLv0efTXwvnITBZ6ahWqqdkjcjT8gik
6HsiuPVv3y+fomKWr8trnMizsqZ7hL9z8dHK3+oaVqVgcBTTwK9n1jIUPFConcLb
qZPtAD3PhYYGKqsi7HBwSSlxxMZ53JLV6omzWC6ady5DY46YirCmCW1Kr80WHjvP
FbJVrmaQ1qGrH154aWwr1Q/QCP80y6aXPtXoCMREFuQb1/uOY7hkkZCERsUZOSAY
`protect END_PROTECTED
