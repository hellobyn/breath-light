`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3UJU5AdbQPxMkMnGKNwVOAdqxfmNtDQCyZh4BYk1vzrc+2hKUL46m5cyLuDcA+x
wA4681UFRaObQBoagom2BOyNLB2QBpM0pvGga8GrJWejsRuZTX0E7Teddl05XmvW
SyMnunaAl495RUHEnPFQ9Ejhlz+x6ekENCe18PTw5cDHazKt4mJTmkgiml6MuiAk
Wj8FAOGa6J/e9Q/zh/XeS/06ZMJHpNp+qQLOIndyrnJ3g5t+me1zwiuDzjt0tTwX
aatvHXA/LUojco7NlbDivfu8X+OHykdKpNdeYY0h7aI+/8IQ+tFtohWXSjTPb6y7
rhDa/M/xXzjy/mRucuvFnGgOipLcnMtLEqg9ss8ApgPvkuVA0C1erE440GATfC+D
/Ozwob8geQrlJodUsuy7khxnS0SqSukHE+hwjcrULBpYC+Q9quiD5hati2KoAbft
Tihw2nDsUD7pCfPmurMR54JWAtF/jX66kvj6loS134TwX/jzfkwWOJF18Ztys7mQ
HF7jyFNoIf51P2b8qWrBC6SkJVY495bGbx17c+1evYR5KqRGmavgbPXf2/qunlbM
i03d2WtchAxj0qqBT0L8JAObu2ELXdfu4JeYTKZ7fDCaTEvBcpc93AyyEc2KIRcq
v6p2TUpn636LQQUrGjoZ6rpcNKUyeeasgS40Wmfak+QbONGImmj810iQpmWq+THK
MOO0+aayNaoGSAbbSCM3Tgj4iqxJx2Do8l4KMVo6uePMcUwDsdcqLgZKm6LnMv3g
/WcvdW7kGnVHvsMLWb5wgvbU/ZudDKcBGnSWnkzdohMJH0JhSM7fosxTUjX+9EfA
W2BJlz4X+tPNcaqmO7rlpfIMpVvJ+4MQPVp2fiFkn/8=
`protect END_PROTECTED
