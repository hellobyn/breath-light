`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teht+ERX0DyQliRMvxNXn+T8xptKLpCGqJ1cCowRCL1Xf2OvEACGHJKbzdsZ2YDE
bhoY0UMaTPqinY66sqXq4QsLqGELZgDAFbxmUEHoUf75gQZBpBc42X17ZmzxacdG
7hyVAvZH6UBhGz8vSVJigB9at4ZgUt8lgL/2H+vrgEk2vla16AEmahgyM6v3Zgsc
LdRjr01KS68Rp2c9wjpduID0HQ5wK0PNYNvP8mlqGoSbfqLZ0mEIXE/zWdU/bMgj
nTs139q56Gpltf5TY2ZLO5EUCBSp4mIezj3HvqgFmxsPlNA3IjsYhXuvjlBR0h4B
5K9iSX3xiNajdfLiKjRroGHoOo8i6jz0yw2bp2PZ7mk=
`protect END_PROTECTED
