`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBYRL/+8YiaFSHbkdBpkpcE3yR2o0oSwhcGLOyyoPDcQxAEF+mP1SdMd3CNa/z6r
T9lEtsuUY3eGdK1HyNLyYhs2+5CmW2SpzZFSlAcTD2pgWrwn831XUUJ6tBGZbeyv
Go2x8lSmxYbZGB9GzojuZez0iEe1c6DTLRJyWMrCIpPdsgaSz/M2JkdmZ7tddW5C
PGSa80NlZ/xZk/zauvnmSmtADC/MXV/5LiEuFUftwNkYAT8O+FxP8yS2jR6mueAd
QAaIfXV9rRireIVZtrID66c37hJH6YjobgLfaKcTbEJLm/7iXMVc/Y6u1AKBlQkX
nGfqNuPdMnZli11zWshfZUDktq8O0asmEWABGzxJkJBYbdl3HLPOH3/Qx1sdxH2w
DNpY3v4XGEPpzehYUM867pbWJg4N6xtEvynX4ioXaO3Cg99059EYJ5N/eqeigKDf
7cPtzs5Xf3G4cwXMcjDl0qJmsRBEvq9FW2br0M2kHV/Uru6paHpxdX3wF7y58Tul
wmuuuLSGVcmn24q8jEh2DhX3cDfaO8BKijTgbrRuP3dsctU4ZZcdaYoMk3/2ZpOZ
954+lEugNrtzixQVWlqzsDiGftrqyG+dt0efTt7GOcbYSU50kAQ6LlCyK9Q179YL
c0TOqIM9Mt25+vyPbr8Jrt35KuMXgdD6sd1sCC/WaFaS1InFgxUxa/ltH99Zjos3
fTa+C1Xsfm6EVNKqOs8bigmr9Ihzs5ODJa0QmHoBL9ioQEbzoYhrL3Lbix08W6Wo
mGkchcI2292wVpRBwK91zQtM1DNozmaEoa2aie01e3GaxJA4N7G11vBLUEt4x8uh
W9+aKo73GPDv5OvV6hHBEEL+Vs5PXl2YCLX2BESoVPNFbOdHtzCOV7p2wxFmsGOQ
gLqIGLjGqF/Y5/A3clqsKzB+xTcl9kxJyK3HQkmKTsX79ppmLK8Zk2elGCeWqrsX
RPsTgIPj0tRYxIwZul01qwevYaJqriVVJqeSNo893pAbmRp6yw29+tPKAcg6T+sL
lZbkkDGko4S4M1Wf1qefo2Di8B7iMbadp5QwPyvskxwuhoUdSkGRCP6JFWvWnZl0
9S9NSGsr2krpN+3s0DNUtcd9as+qbWnz41JUFzLvsjnhwb7MoaG8EB7NFXUWwz5w
xcKTkGoOmToYQrUx/N9b/yBUX21k7olQNv4kDqshNWbN/2mnCRxSlGjMPqFiGhrj
pzS/l62uMKq3iQEh5hjT4URjiXdP+cAa3zXqVOObpgFWagG2C/9v4Drk3tM8sCUq
b+7jzRgBMX+zs/JNpEXbNsRpL94K3toEwPiRxayRE0tp3Efp6uT0THBgQ1Ui27px
vyxzRkEdVy14dqNGEh8Xb/0gKKzUM+dO+Qyc8melEZUTkRL/VKDcALhrPody6X1F
qQvOYskLHEQZ+bRDuTQlqrla9LL+q9yi9AX/Kqn2zK7L6KJj3CfJqH0yY1uT7zVy
enahsOizD/0+VWLN5ui7ueraPb08nIbqDHplr6BAzyiWVLWe51Fvga8TyddXF9rs
XiyqjE6UW4j9ZSAPWE5R2IiGPbSUr5qemtoh4sunWiTVXdXUIbVJZfWhwKtOYYAY
9fjebscZJvh0OppM2kCADgFA7AQduGvY+lOxL3R38IxLwsKA8NdvsJnUEnYqOnui
j/7ksz0wzw7FFCXRbKViw8LvzU0cvpzz5oXx70vr0Pf/P124sj2vTrOruLmsXEIT
var0xjEiEALozO9bkzfujpXQiXaqZ1eRv9niqMokd5piOQsf1MFrUc+ZwUxc2hWJ
nQGOwa1Om0mztoQiTKyZ+Oqukzo5UzJySbDTz5tFYqBmksVvcA6RRmxYz8pb06Sj
rL2mqVjLFjlpRygoSOGYsA1ZnPEmV85HF10zkRLMr2QDqSdJtt3hezaN8bLhzk9Q
aTyjr8cAFpAmcel0L5dc6ltY/E8YHs+ufohZ9/ipIiH75dSzQjIpeheeyIiRrU+K
H1qr16fY+jyYEIAxDjr51CXkmLMPEhDApFQs9QkP/tvlEqGxXNdA4fomaewwZqku
rvnMFhVXUD467KW5CA9QKA==
`protect END_PROTECTED
