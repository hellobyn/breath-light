`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20vTkzhgivVIFjLa1zkC42i80ISHtU4pboBp6QFdHBUF9jKma0rPyrbU0ZVcXKOL
iYXxfzTBn/jdHoSC8SCxuFeBGNmSY0xn6t6f+PobapJ2uO4r5v8MYeHggZYw+DKw
FtxAHCFrE7dR04QdE/X/+UeNen/KlbyA3kdzij79QSwGUU1zJMRVEiJtkctbyzd4
0JGWa1LYCNtZhj3XNKrgwsGfaOUxNjjINVn4YXryLE8bZKWHfRxPfAVgbYCC2pxa
0oXYdFPacX9oQZsMHxDVzSkKt4GPdpommZdaqeILLLzkZa6IwJPRGHGArtLLDW2Q
5Toafhx5DFzlLxsLvBK9ogX+nCYtgHwXFB+57IKqarTdi3EA/roY8uZ481veECtP
5I6hFVQi7GqzNy67GssgVzAmJDjWduvT1a8QoIWUC7GLNurajnXeJabHFMEh80Z2
s0QgiGfd6/yqf65szpyMsPY5y5Ofw2O70vmdc6b2JWsyvhrMLGWtqMFW7tjjs3D5
Y07udCntLfXyZGlhG+e2nXTieqpalGdygttoAzEYY3uDdzYfoI//JAjosl1JB6ww
hdy2XNmbESMPhVzD/Hnr4qSzOEIs2RxO/qmABCLrbByEdauzGL5ThGbkR26RhxJY
MbuXLWg3kfnHR5b7gPwL3A==
`protect END_PROTECTED
