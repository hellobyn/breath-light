`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkOV9RDqijbKZqxJVLC8HHEE2a2BwvPSS9LDWhojU68NzUV9zcbPwWqMPJIVLRK6
eQBHRqYcgCSLsZBIjqBm4gbhTWxx2FpGKV4S/XRQ+9/Sp9ckt3nyryLALuToHT3n
Ls2KSkUEGIlyS9ZXm9xYTHwRNJlgkDBekjPLgdiz/R0esbt0a4T4CQmW7bOnG65o
2suX5H0VHDERMZe/N0oKDSAkKGREtFLgmu+rDa8q4+D0dM9d7XPtnJkQT9TanICu
BC+NomNfELAe8wKLY85sl9YFcsawECmG6mNFBuvI9hZA2tN2oSxgKzaxx6FCp4as
1QqZwiRGUscKj6+8FArNgg1B9/2HONU8TRFXv1i+oYSyNylD4Xg6Hl4MxIyQaNgK
g6FuEoRnIzyQOq9s7kvwRgINdd0tO3P3C5LSisVCcPQBomUwZoY6vJgeJmvurEgu
YrlPdVIBOBT+LGdwIHX+wwoAI20g5AgOv1sjNREusjnK3HkXvhB6a7v9bci2ljIT
adf6nXnpMpKu6bkZzV95KmZUJSNxLsR3OOstJ3FO1ajHOBa8NM5d+mdRsolvrNIA
+X9ccx5vipWA4PfQhCtkydGS9uNkAVS13XsU40QWs2kNhCfvtW1mHkh64Muom8s4
qK+rLAVGkMJ5vU4bfGUzGzLyP9y+F7EJ6PFHmvaiSQUQa6Ym5GlussybF+dkk7T1
9deYZ5SWfi0p/ISjj4bGoIj0ezWBTYIX9Jg9FbrxLN3g7VizliIeSe025pFjZv4Y
2qzq5YNMX2Y2KHDD7RpLatWiQxM6kqjmjuISVD86Wf6UPGUBhl9o1Kb4sfTTcW6P
4lrD3/wgiohdqhsynDLzDPKJhqxXwlZhPqz0yz3RONda72mP+uZImwyx8WBAfeD5
`protect END_PROTECTED
