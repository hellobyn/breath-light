`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zfu5l8zpgFi6XhR7rbZ2VgVz5gPCeoODfzV3szIwvRNfSNxNaOrxWhkUbprXOQwf
AoX7VInnSiK/gSMmplbxarY3g3wyL5HP3W6aMLzFJSkCVyXRDmZThBqC0NH54trP
Vc3LsTa0RGMnhwJlJcIaTg6rQYqqQQAUgQriCg4CyfCqYWSBjWTDn4BglcAbHpKq
Ql8zcxymjRtAjtra46paggdWhgoKE4EyGYyTOn2mRQ3QKlUPVNz5Cdkn+jr1+PxA
pHRzAIM9WKW7PZavXIFBQpFAgcTSNtQTzsiljCCutq8S06UlVVuaPixPON51JERw
bHxjwvO69OkcmuubOzd9+b6/ixoFmM/JZKZLjaxVQ6VWV8eI8/pqFaldRnoKxNiZ
5FkO6E1vHsgWS0MOYb8eqx5BnEXY8E5maUSBLR2MSkF3uImChtRam3MdmmYl08x+
msZazEfiUYxpPM09b7vjPbE5eGQ8VJ8r9xkvNIvYGoyqsP0ONj5bDEZkjTQdQxL9
CRd1mVb1OSmMh56auycBFkLp7Rx/EisaO2cqOCt3aCeqC683R+NKK/ri/6ngJlWb
2ZO1dd4zlrLywvruJAwdjps4/u6Qp6o7VNkUEjbnfEVNNPQqTCgr8/+D65i8cjf2
TgAHCmkrRObwrPaASTEJFsYclDEaQnb6JB7nm/kEdFJ6y0IIDlhMekmTmWEFCiUR
6jAkmyDNe8DMO2nAswkjm9SrKm3v7EoMvTis/sfNftsIAvWmwmZ7zJAQlVF9LAFt
PCPUVMbXOsPOS5VBpQVR6a9cd6Oq7yHF4LXMwMLBqSjI1+bcTDrQuUdFWZF0DSzn
2iDbXT+LHLbwfBp/kcXYcJh+I0rwauW8SDcAQeNeOfOmwhc2I8NCF4LiAWkmF8oj
Ud6NVeBY/r6qJZAL/2sEoHFM/TXtsgYVLbm3g6PPdH2DvTN6och/yW7/KEod/Wz3
Pw9SQRPxWQrs2mtJLhZ92lQItmyRavOTLQxlsbgARmFOgb8+TDtn3BsinTdHKH18
llYFW5vMsdTXAyLGfaFiW18upJ7FA9I971OaZnBxXBTNp1BFtwpk16gZ801Oh5n7
KmiRoabl/tiJUt/Zhd/f38xfLpTc8hu2FdWWMBEigw+dKonjC+M0SypIFiVObVIp
n7FDbrhewlWKW7cnZxNUQJb91xnJgzFud0TTTZJt8avFRN5epplCSH2Etp06i1nM
wbesz3JLLmNsLefmVWYBlnvriz8i9HBGYU/Yklady6B/HL0uuQq5dgPR3UVk9Yof
ZQYntaLr6enqi6TD71A+EyPzfXNIjqr7IV6tyEOV4hziXyCV1svgA7r/eWAFjkYh
otp/+jdo8X4gwEel2fhmPmx70HpZ1kkTvbQ6SNM/2FDNZTBk9FCR/eTBnL9OdydM
wMQcVKdDMAn4ViOpvqfGWCzkR0kjI+4kOyeoaGaXZ/x8Wr9GdwQHW+Pbdl1uCH/J
tEVWEjDfmDGF1SWGjZbIHXDJjz2lXOLlskKT1CnG263CmtgVanHFOqJNw/N1jKqD
cRbvGBhouHFwznyMLJCek43DaBw1xyaayb3GopN8nKkLBrO8lZldnBMpR/XAv1+U
zjRCtHi+V5s2A2d2atHD+qpM+NVPOYVO75jlt4vlLhIH36URTTOvLbzF5sDDxPRT
gRkEA5snjefwJiq169krDJo4GrdKgGrmkR6eOlZ9QE9qy32HQI4rGyKT/YxuWXb/
MeDFwR5eyoBtArpka7a/Q2527JS0vnVcVJhaTWu0+4fAAFo787BLbInsnvtllZvL
lR6lp2uIEdWKLjAR6Nj3caR/rwtx43kaOtlgBwI3R9vge+/DrYHwGISnbxzBdxiu
mS+uWTkVO50wcSC0jPsnDO8UPmMGA5nvJX5hf0fd1SJN+etjOrHU+Qgsb2/NaR8g
ulytS3z5Vzsf89yfLVFUpSwVCF6Jj3UEzc69GbfTa2mTuzISNCo2s8miPI1+8Ale
8atOU5jivYUE2HnHoTe0C4LdzOsw0yR3LJjy4KnmDTjZetwAsUGZ3/G5VCX8dsas
3ElD/XFghmybzwRC8oU1+eI7JCdTVTaYxfk0gwvS5gfNR/Q3MGxUijsq8Lj/aaqL
d2dDQ5S8Dd80UgMLJzXT+RWlXCRoZZ5vr7XBBr4gNy9o3UJaJdUWgHp7zdbpR18v
xNNIR9LcX9fmxSPE/kTjN68HNbcbe8bAu41q5+2zAnswubuXvP0CJk1YWSTLvhPw
yAnyOwzPH4LyLMuM1+omH2jQ4R1fQ7E9iVh85baFGwUYnQbOcKIfh2XCWzGhh4eM
iIN5K8FiKXmCUh5fbwYEZcOPs1zkLYdYh1nIdEtFxZSZ/zu4KtMd1Iec9d82Q19k
GgjIuEA2BzE9vDJrAR2D33Ag08dMq+SNBv4rN8k/XoLX+i8l604J4m9Deq+5isYg
/BePt7FnRxOp+EdznaI5/o1qPMqsfd391w7Glu0khxpWmf5/jokOl8tuqlTGEjWn
eqhynt+7gePJONMN/pnh9rZrulJ1zz/zFpOd0PPiYnY3AyQj1b2Q5gpQaooJXkyt
5FzSOtBfU5/fRnSC+wSaDDyEGVtUxR6jg6Jxp/cWAVo53kyJtdos85LLnm5eVzeH
prMovJhKD2fLJzpVhbxTSnRJ/hpaka7BqJuczrrcmeMTj8eTi4dOfk74E0J+X12x
r/wW95H5bAmyFfVFhy1StxT3fTZAlxD01gPU9wBuPn6ikL0q3lP26rx8XYYLr5yE
zx50/wmx6ctPrP+zs5Rq0CF27FEQD8ybKkKyplTs29erHYOnDrAtNaKIdJ4xOC0b
ANln3WDT/N/o26KH1iKsBpVD8FkVuFyxkErZZ2DISz8=
`protect END_PROTECTED
