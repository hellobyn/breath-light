`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MATytcS6KvdzBHvtYEK2ySsrRitClKkg2i7VlNGPoclsR8WRNzvG+cyt71oBZ8xT
ZmISqMsRfNVGiK8qaFSK3Oit6fuD8QcUSRTxe9JuCqaXAwHDAZrB8Vl17aGc4jxB
rCMsPcwp+hRaRttoHUubfoScKgyh1VjnivgwOBLB2hBUkd9YI/pzvJHUja6dfSpf
9/3dRIKd6uFWyL086aeFlQzgHRUqb49PF07ok98NrEp8gLuDxA57R6v7blVQ+5Zt
0hHbAaOWk4mQPqnFfKqXjezdbWXTohBM4CM94VlrW0I9tZDly5yyFKXbHpCIUnQo
xq1zbhAy0LsyKYlGc4on7Mll86Q7Cu7tfzDtmS1OO2QeKEZldJgVWU4PbSKAhAAh
n6fMZTInaiG67sRX+K3JabWTRtIF1nT7ZXiiph+1cIbKtQL8JhwmZp+poRlopnMd
`protect END_PROTECTED
