`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ofy86B64WEw5mfxQtYdz9b03hVRSz4lrxPMTO9cBT6J5uOFksMhhVFpaGKlRKFY
RARjMxxmfp1bx7mVqjJsmIm0fGRakmjfhHCc0fsHBKB2w1+DIRMWt1LYKV0j4sWq
0tD2RkDkmiVJ7SWxwrd3fvBYvWxmUnUP74J4QKkiac7UF6wmWgCYPlwYg0mIyob3
0Ns88JU/SrMORMbVq/UoeypruJwjdgYX6kxyyzOSpd5D5l9Xv4wUdKGl6K+RyF4P
OyFZd7RrZdc2HU5Ed5DoHdZ8/4b7A/iJbBM4pETjsfIIVICaacvKcdUNtLCJ1nI8
OMYUjeLwOoo93N4FSzZEi0A/GGokkVhcEl7ECvUgQzhVobrYurYZRVaELFdN2Fl0
tzW/Z8aIQy70bs8CpuVicZMXfx5zBjQ5da4VVVD7hsMF4AZT42os9RPmSpkDZjoA
IMR16qYoS3NfJpxYmvhiZjqCOJJUj+o+F7Dle5ISKMm79RWkmerecz3aEnU5fEQQ
hy5iOkhnY3lbLcly8i0KpuNdF5GVjUo/4ARFpYmYzI44Zx0tVvDUg0E9PG637YuF
oWRZq5PI2tEdwfKqnrdSawjDa5PRyQgv3pjpYM7OmD2yDGcHPf36o7hlDmIpwRSN
z1nl9/mhmJIN2Jmtbu4nDiQCTr9r0ZXXk7CLLVwNunIEY8pHE8G9OkeD1cpY2enG
iuPEXlgzU9zl95bI3fCix0OmTdvCko355r3/f/D7VQigfBZ0NVtZCnA5i25PzHEy
fJCGzW5TvqSRo8FbwF5qTTacFgHSK4XTk+uxcebqC6nlabacxAsStem1oRRXeYkq
/ZSwvhNNpKKCZj3arlxigFubkebOGWevnvPHkKFYczzboeGoUPGkF0B+TDT89jkd
OniSDhVLfnHM5MsAaCx8+QKmlpmLDgBcnoPgbKLrJtvkBSqjtG6D70yzwW9CApgz
gLwt8vg9cPbJPwtRxk87Qfu5fkIh6c3gBKCK8mhH9Ezbm/C8eoNsVaHRJ0TxxDMR
k/Qo5ZKQFYv0a+dYwY32yk8nhzIiIAid1zTMJsVUPeav93jUO2VTtBGYCLd2ThkH
7oIzlh3e5VLCtZ55p/wCIdQkLCqxbdUn5HJqGK67s6pi+oYERETfyGK7oua9iM61
T/B0NMn76BFfNV2Tz0ZFG4+gn8ECQkFI+rDK7j5gqZaFmhQpkFQPG+gMk2E6dkcf
TfQIVRi8jSKV7fNaZZPhnqGauvEy+9NCjmzXSivWmziYanwM5zx858jnCq1Ln6y2
JbthfOFQ5A9qJiqqXCU1sGE6mvQY3a75FBHyLc7Hp9M/1Nfjo4mi1rjfDHhj6EwP
kn8YznmKBwdS1KgsQWzN+ppTFu8KbU+QfinFPxjHNqXNnKlqS/k//BUu23UtsAVs
MSaz9HiyZM/XVuPK2edzHq9YY0vAQ7i/ThNVJq5MtYkjbbmdiG+qDV/rly04raAp
yVubpm1/OZpm4rRmudCtujspXzqDgTheqf1aJLiKWm6jJX9apJKTAAKgqIglQgFO
og2D6X1zVtgkfUlkGWlDoxF6PknP5/zs6l8VnxwudAQrU/DmH+6TEvmx2nBAdozg
EcTeZ2ljQHdUOA+IOqk2+4GIW8F48nIRv22zRmTg22tgHnN3WJgDf2b+dJ9lsqJ2
ft4VIkqioZ0piOchieaPbxRXhipxiz4tlvzK/LCn0OARRZokaUt98GDnR1UwWnmg
FRdmQ126BkJ/0LywoMjIvAzZTmlObi+E2Axwrm0gtKJJK4YDCNPNQF2YYWM1X8vB
mC1tm4H29pfVCiMCdXBn6GKCiAW7qu2QxucgZX2CvIoXro3jRF3+LWKVIPi7AmOr
qqWj4ov8b6OAKzHyRbs5Wdh1CgKS5iNQJzxQQm18rgWAcL7k0FLFT4mr6u6CYD1i
k+nkVYSV0bUM7OIXZVMy83EP8GxYVcdGk+Yu4OwsaAGO3m08MjcdenlBb8SEiXEJ
rMCabxEkHvTk4w1MoshqDBNjzjuQUtZ38AeTwWKAv9+tf/29Eg4cchWiZNxDSDMa
/u0QGIdNr845WGeG9UKnNRbQrdf/vB1c6gdwH9l0jCjyRS2m++kO44I//NqvXGpK
8Abq9fAkCre29104qvq8f/1rd/gVgSDPHFDrqRYbBCiZaU4NKZuVC3yzi/foQ9H2
nvF0vmzTlm7SDeziYw0AHiFWZCkvv+lD13q6Kh+Z5VM2bw5WNZ6MEMAsd248nUpP
cWCxTOztcMC9TWG1nFBAdF6G4v6NzQYYwLgBKQ5pIf+MZVGQLrzi94F5Ghxmlr8p
2wGERokYarFuhDWOKqfGAVMXVhknjp0QmsSuRmeYVrvslVEJRM05qBDg2npKI0Xa
M15PvZUBc3uljBTg5MckrMWTiQ8ZflcOCsUNPhYiNWnOGo4olOqMMewk1wImv8/b
kGvE5FyPe1UScKdqTM6fywzIWcQfv1FWssDewY1HOgDmkRrQgmoRWET4UzUN46v1
6d9zWbYE6XjcTM1DxvM0MTqdTDZwc9ioTkvcK6v8fvMQBJNweX4RS/w1BlQyuOQQ
CH3PVAX6KZJ4kE9XwL0FBDfoZY7Y8NzQaR2qwCA0JuffagkUmBfQ19qX5r0BLH5U
Qmertd1ub1BwlVcIS+Kmczr1ud6IeHEcLi4Bg7ObeGKzXNqkeUAZX0kJ1w0uQisU
9KNO8doV6W29EbYf1x+NsVo12NEPNmSUaHK8Qublu2iafWQlicqpKAAWIWD8myrQ
tSlUhB0oUEb6zQMKAAJrLtC6ce/q2xWARlhb8zWuhhufVfJpgyVHAL4kMkbAJgM6
Opt5ELSun0kZZRJM5z0s/UTyDo6HLGhn9woyP/4fuwWJ2VnyoHKh+huFxTFRbXWx
+A4cJybUdji84rPYqUH+pFx/zNjnz6FXF0nifoBi4PlSi60torw66GR7MYP8dnHb
t+8IiTarljubT4ECMqRF+0ZV2bOUvXe3UDYeHkN5JA8XsuypP9IT4ql+nnoCGmb7
JEeLHafkevA7q3diUrdNR2g9kVdshyPWHQOaJglS5fYlKbj8cfJqo4sYUwmYfc2V
IUjdQNFdFGA7V7yGQ10qN/Ecvsj4PqqAlsmZI5zpbHc8HdqN5mwv/vU51he4Doue
eU0de0dNvdtWUb6uvCYaIYGRSngI5j0Ho3mffxm7M8kJH97pJHFI78VGD9W+A3KF
DJw6xiOZJIqw7967q0WlnrG6S4PWRXYrLWn/3liFuBrdoXaVCayp+L/+pIlAugnW
aPiHMXVq/o4Sb7iq9HvYw6Fbq1KX6e0IIJwzw3O4ogiiKGrEdjZikKTk1RW+WCY7
X1baf3BX8+zl4FVdSkqu63zaNnPlqcWNbys5WI4cDXj+CgiIcIGd2UeuvLBZ2IC1
wbkgYak6SSKiGll2vu8lN+WaQs7fs3+M37x+yQdldA8t2hSgPlnGcFjxaOf6bgdf
8fN2KSwLJ9ETZ0mx53NckDV3GfJW2brflZ9U0NQbs5xQvEBzHytX941MoRiOfuD1
QjXB6HtD6nsu2Ad0MKgjpi5QHH6yAqE3/i9flSN5bl51bVo6xrbF4mLGg7VGL0RH
Xm9Or7iWk37d0o4lpOxtr6dj2H6J2BMbA9AR+8ah2GfYq1CCwE1/I6OKENe1bubH
6dZGS7U/YKlYFVbt0bsMzQej3ApeKkmmxOSIkp3+iXbu5B1wbEVYoVF4h3v1tuaN
hf5EXBE+1muOyyvaAqK/aZSfhE7js1hDowHi4Ppd8bAe8Lb4ByaKTDA9yP4ysTmf
yZ9wkly9ggL5ZZYRrL2HH8AOS0aDpfJznb0jrJ0zN0+y9zys7pWCyMTUbJii5DiL
YKw1BMLfAVBvwnw/bZ229hB6HkQMi23SiKm82fR+jOy7VZxBMkYTe3M633+sE1rV
j5i8tY8rvd31ZsQURn+F4pJZtE2RO8DRZk16WWajYMiTY5GJJZUtTig63IVmg/Id
9LJTBhEuDDQwe9W3VY0ylNaiK99wlJ2y94mW3EEE1LOUgh9TZWjZ/AgNxJHoG9bB
3bU8HfGEvkxlpLbPwDPPZxul02VjT3zrBTleGKJ18p9iwwpmABLHDh86UP0tPUap
xfPQdjrowfslEaRLRIQq++bAWtA45Ti/pLxMUtDYJF79FY/dkHMm+hTKdT8C3waa
fr66LtKLoCkdiRnS8uu41hFXCLqwibynCBDawHICBIeLHGJtacO2s/agSfl1IZs3
kHAW10mGSyYgDaHzC5NH4jeZ0jrM5KPzy0RQE6hEWEdZNYufnSp3OWC48y0ahid6
dtwEqXj1o9V7IBcma3XcMOBe3AR1KXdDTyG8pRFQxjRoGJ2oYe+GjbT25VPfVr2l
2Bpfot1C7TJOIUBfcJkQaEinYV2OTgI1ochLQwr9/5EHqKZxdOHI7OckIw8nc4bA
JHElH22J5VH6reTpQ4YJQHTjHxIifTzNQfH/wkzNKZY99My49rHx4UfGNmlRck3K
jJZX8VoKfnlDgXq5OlHeaQ6AZc79MOjpK0p/CSJB2pZ85oyplBFbgxS+ml/reOlh
DecOBdVMioZSfv2JaBSmGC9uFRUOltDbqlCEdRd83GzDmnV+H4lHDp0exAKdZhS4
gT2NMMAxudqEwEQN7HsGNwk/BpIG9EEoEJ7lKCD3xIp83ecH31kcVa1JqIYV37tc
SYiLZmfqHwrMyXBfzZRTGSEIp2xF043b0In2y4ZYKqbtW5rThXw89YYoOuAii9rv
1uGDK76ktXfv1FOSwMAyeZctNHUjH1vLXZ+ICBbyG7YC+5KmNsB+RmEO8sdY0mxK
3V9PdSf5cBc5IQ3ElRBMNYHqOqkGIizO3unnq7VKfnfhxu8QakuqVSAuCBNmF8HK
K8rwHORrgZJBWyoAhBFved3Zm91Rrks0PMjGFTT/sZY0ubaVvShLzBKe/ofXRV8D
sqpqjTfNiR5MFH7/NBVAIHgw0vSEJh0YPjBQeeEtrV2sA4+n9C9KhdkTxEy4LUgi
Vm437w0fWxPW5k/9L/UDnw9xuu0C6j6HMUjZDje0Qb8eku0ukcrrxDTZbrD2qxbn
tfHlOyaZnSj/s+2YDWHzWQd9r+/SVgQl735JtovFWmcSjt7OS6c0YDvWPFywdocV
7pI/g+tEvnbcWmlvUJqqa01YT0vy66+dl9jTtKIZtpyJ4A77I0QnlZ/+gnG1Qo7t
GCVsOWbROzdFnQHBBraQXpVda6ReMIG2Rn9GslFIkk5QffBAVsyDOqy+FrWV5Kbr
N+WCwscHJYSxlNGLN3CvIFSjLPSBlDzU0Tu6qyOpFCh9pGZGtGN8OWo4R+aJouq0
HDlYwMml/6Qsy7F6bVaESoK1luAsq0iR3SG/zizSXjgGSxjPhbLsXE7I+HWkZwOE
ZnDerO2dnDwSlco9FFS6C52kFzg9XhWIJ4QZxrE1Zl3O0DXK8JHFiDvDUBn2yj8O
4jNOJFSe0FI6fykdvr9PhCz3y5rR4rPDZTSm5wMKAvMIMNX0wiG3FiVRd6Pc3GPU
DQkEsQ9r8zzt/qnENX1TKKUvOugvNBCQFSrDD2gYXwxlnSWGIGPnacnszUCga2ix
R7B6+ZMmPIDS4CNCPsNZiyCaLlxB3XQFeE7nXbtQTEoY+RrV9BtKZKw6s23kYYdb
Bj7S6cTWbGnsFhAcC5PvqmaaggKDFe+6haQSA2sRX3Yu1L5b4vsQKfmH9byiJ7Az
ucBMJtjiOe+HipKGQ2W1/9gkHuImx8Zv0TwDSlSCGGA8uzaVFUiKiYpJJ3GLY+0R
8Xef3iGvK3ZrQFUVFRzZzPav0N5oTaf4TmKOe+NcIH4P7ny1r39OUpdG2FuaPiWu
LMlKpXhcpnp+b5W951K4JLK6Mt6m4SDPUin2HFC98y/D7g2rrZDUqDOUysUp6Khq
x+h6DO6m7ksQgGb/d6l9SPVFAuvl+5QU4YLjJOpJsXUCNbPmmD9WBZURawvcVeLZ
QpivmKZcjMLh3ZukihOUv10kuBxzV8QM49kV/HAa0EGN1Hwe+HU0QYiM5PzSCUrL
9HJ2AoDvR8YVhySEYqiErj5+UT2Mv0qZMiUtiO5s8mKP9xyksQQZ/NpqqXcP1GfK
Yoi13m9VGDCl0CvX7MyW6zoWqO0/aoXNYK8u/iTP0ZVq8oKKlkags4ApLROxkbe1
bAc5FvQ9eyTDJQyA0+oeMODNlJth4Kq/kLZVgUtKTt2yacNTTRghizkeyE3w9kDF
OMIdUarfGmfZq6wibyPNc5IDh9UgaJEWPjJk/Mje8Nu18PaVUOSioGCDH9DBPxP4
VjuUO79Vet1xYQMG7/anAP5ls9ezIayFrKvdKHZV5qg+9Yxc2mXpypAUTD957m+N
WuuVyS4xog/X3gfpl7emr+gitCoqSS2nMiV64ouBnVW5AApVZrHWBlD4vfCS3yNU
DD+l5YTyE4JBlMLlLLdlhPUArn3zj+4eRzhGqbh6MbSD700GJTolGnGp9FyeAhfA
RzNDuMVQEC7ejOsnF44nhlQ6B6mx3QfFsT9i7/0f4DsnypVxSPF9O2OmYzn9h2p2
9fl5lMyPVTNOEB83Buqqv0/L3KvFv0vO6VkFlC4QWJlDpY77OAFWvUCfjGgIu4wt
f3I3bv98qPLtLkuE2Vw+oB77psWfTyHc+KPmWEyk18Hdrks6z+taYzz31lIbFDXf
FRkS1v3BjzE4trG47PRI9V/ruKUpuIR/gsxT7sdD0KTnIqsDthGlihdWDdc7XkIN
ujFpx+CSiTltIaytwOEH5hhvKqc/JXg/dv4RWhS53CBlGjiOz+HeqpENwI21gOgA
GGyeAxsheLGmoBzWwwTgCzRU4eFOly5YS1gov5jR3ZB/KgXm662TN+CMaQFvlb6H
b5hat3ukvfZzSDN9rOXutof+jkPh1GakwjGVHT4/InU=
`protect END_PROTECTED
