`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPLPLMJ3weBBnOjWuGgUGDaCCJ5XUhRw9ii7vpnBt3WRZtzRM34AEUZtD5Yg5Kf6
BEVkZq8INvY1QX4v0/RIgL58pEVM+9uHSFAa9X92x4Yxg3gFi1oLtQsN67Pj+D9k
02cgYHun2+IkWJkeWRZHgCZGaQxvhQNlEvChk+0zSe1ny/yUIPsM0j4d2zeK/feJ
ouCuDbmuwNxq0uelSGu76L/m2U5IDjbNit4Q+hTcwCNqcZyCmeR0d6EET3moMSds
wIVvXHuP7O4pnSrhmQq86M4X3SZG/fyzR9eRzerw0xJ10qlrM1Yk8aPw9VtJmjtg
pR7x62GryAJ9o0/65xST9oHRYx8K8td7hUSbhLbv/veknOWMeWch00ExumIxuU6U
SR9VuKdCLMcaTAPRJ8q7GwXDr5mZrPZBl/Zae5mjUCjO7AzTr7QPfBOTyErsBqHw
NFQkQzs0dJPgXncjLAObMB5VbOW7t1h480cTCI09WsKMkCuIW7LKG221naHbMzVI
mNGJ0bAktmz+JOGnwRz8xSDgyPEja08J9NDPeMOHSs0oIZ7oYlZ6a7SPRqjHnncr
V6GiKwMG1qT/ui63Kjmh0nmTyZhczW3pPIseAYfih8h5FKAc5Lzzeb6hfqAPz7tY
LgvmawicY1ovM35C08Ioe7XrMVpnkKXI0oEE2vc0DcyeFzvHLO9diamzqi5gA+up
PLeCSNLnctCJOKTLMBtQmq4Nfix/OoESgle+lJcTjut7bjPpRyDVTSjlwnqR4Wtj
vRq0r/WJiRzszO5X5/PdgA8oO3IPgq85E8chr6ftsZaQvt+h55uOfV+lFzoxevCg
9DWybvNQhuGfACJoPP/8X+taqJ1v5D28RgOphOBFB+Hbtl17vavnrViXTU4suqXC
`protect END_PROTECTED
