`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZ1KxgffzqX9ZEHwPTDv7mAk+QbiMKbG2tQ1hTHALHCdB7Mcg3NcVXGg5Pg0LiYi
PBHVyMKMfipgydh/Uy1gbhpBmjlIx4zyVej38Mh+8d4EGfOF3rdoZ5qIk4iMe0Qx
Slgcj78vMPeODIChX8if/iKLuf5so4kL3/BbskU/vhxWujIwffv9zD8VgKj+OI8p
ClKIO3FU4be6dMjezMqJfGEnlSzT7DFVDJfJrH1NGZotrOZVDIZPhWu5S8oxBs0N
X9UjceGEFxUOOjpew/XGQ8qO+QyRP0ye1oGPZs7PZqd1FuYfjgDeoywWGJam1gOo
kODdoTgTOxbvt79vbKjcFurXJ4h3EZG0+p5G75yUy8oMuKWAlOcIXklvsOIbC9N0
V+5o+W7NuPjpYanjFl5vil156xE/Va/UeAohGo+tXqDPRt1zZOQmZ0xJuIqPVLWn
e7sQ1L7rc9ox5Q0DphSggrdww/oC6d3xgKfLK+JbFmirDFXc5XFQLpa9FkgRYJOW
i2F2d/aaKyH1BcNEPd7HQqulxM+pHv2ufN09D5jLvHnrWsLim18laLj5F1Euf0Rn
m1cy/472x0Qbs4uW0xOzIzv/1tGeRrfYY6tqxEkI9IOAqjO5C7ttweM/DnO8FnGs
ZB3cbKkQbLlOiR0dQdFGZYcJE4rHddP3yDbut4gzsMZYpWJ2Js1keoHkx0EBgN43
rL7Y/ykwGpH2sFourwdeXeB4ATgQQXD/CRH2J2Wnu/0=
`protect END_PROTECTED
