`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywObzGuiU0LhlBATQp7PKs9h9NYZE6cZBd87KF18MmpLtfnjd7+Fh1T9L0rbffaY
S/spy+jOA8wY8i9M1qOFy6JXKHauGkV3eogl2U0dwaV9ToCw+5Q7EN9qtTID8uGM
hSMLSOq+hpZJcLAmKSEEkgAlB2y4JHY09a5c/3U+Hv5Nzgsm3acxTm42hClDVUAu
2h596KujGFh1uP6JrXfqbDLbBejSWwfgkJEUXNaHg0wOqnXH5XHtYYuPxEHIQN6m
EOAWkoqyhggMFtLELtFCJM+0Ugvb8sgDItKWS/RFRX1iaB5wM6maoOot7pAkV3dl
7ZfFDFjZBNCNerfWYQ5DvzdHjmJApZxSveOUfDUAobnKZcGasibDco66ZJAIngr4
6VQyCAih23M0SwHtp68czy0Fu7E2CmllWcjJ4jy7p02sUcWKx6ItSIwhT37fvmnN
edlGY/q7zGdnLXKc40wwjTNdeckUtQoYKtakogOPTIK+0VL/xRc7AJRSKdL+DmBJ
NbgHj4rPHgeHyku4syJubxFpmgcsIhVOIJSQYssOmm1+x9+1+sZmGA7MKe8k5AcF
o36XgAELqo3rI4IXjeT/ZyxdmHWf6LFRvA+2KVHbyUXowXqFYl/DZJmt7iDlZwzq
r0VSDfnj+YmvL+m2w/KpDIFAmbLq8KkmdWReMEuQSFzRDHL9jNh2ulQytcJYxSNh
mop4LW3WwTxmkwupREsDwVm4HtbqIsZR16HgnGg0azJ8HO/i0kLs/UVcPofNvJrE
u2CBigLBTOBFRbfzdjKLpbBtsXlgWQPQOB/kUpcVheP8x/DSHHhLMDk6uWO6zrhA
7M06fVLqFGOoj8YzykkgUgrXXYyhYoCOpf3wDbLzwz50OLLwtSS3V51m02QnUY5S
+mcmQp+aLBLsWwPZvnBJu8vaSAqGq/F0r/4CeMNW0/kfKiWuoR/bIzpVg/vTIBg4
RFF+w3JXBVAgvK/fByfMprcAJmxoShBpwH99kYU5qsmB9Pc0P3K6jeoH/S1IhemQ
Gm3kj6xHk5+ckcCFh8EegcdDa5fj+GMg4OROwARqbCof3vAoZvArBoXsmDjBLw45
2bTvtqBSOigVNMVXfFWLX4yDQcL3mT1zAXWgfk/BnOARbwZFcjnM6J9LgpW//R6E
kv5lZ+IwL5C1NkzEdimiCyctuOq4qoNfY8BL2qoeEVVZvgjJOcTwEqFabX+Y+jbh
jbE94BbtyAKe6epAEnBBu2YI3B4SC27tkCedTCHEvCZ5Tnn9xkv81liA0ry9O7bm
UK+gNugptEjSIcRNU7AS+M5s2VWigOYJNyLKulv0nvnnsaUmRL4wFVybqv2JPffa
ml6DuRqNVhW6PqkAc85vopfHO3uLxnyaOdBcQnA9yDJh2gt/GAf/FAcpZmLH2kyg
jYoLIQ7zx/3ExFbnlN1nLXUcHVLtuo+8Xw8ze+8nG7ZID8P/baUwOxZkZ0Mcu4U7
Fpx+qOEsYGqNItjPHCC17L6siFnmepbiyMhryjzGIYameNBJPMeqm0DV6rtNlAzo
5G6nCC58fiGxW4kxf79YRFzdd1wd1qNbJDSREF3hEI+w+yq7KfwMae7tuGAIgNc2
QlAdW7bfTSHolnQwPTAfxKAxaApj4VYt4OJT90rDlrvgBqkyu9G2726darPglYcX
27KDFLxtB1RE1v53VTJcA++EoCG322/BHmsYFWIhUrbehBUnaUwX7KJJRRdByD40
P3TI4VO0oTZcH4cfjfi5GgRJ/dfzyE2kFGG/CwwXF2f1weqsnm5iqnKFbHA8MUj2
oTCIp9gCqb9fgpB1uKpHaAxy/7QqGOd7jIY3oDddG2Lh+h8RNB0u0SHu5cylbjws
b4+2BDVV+65MvQapSCbhPZxNyeI3iKkkk8mhdNEzrpLPeaW3B6VhJtcT5hnl/7AD
9OHISR0QAPhQ7WRzOfi3Rjs5AnkZlsO/cgTjuySNnn9hdAMeLxzC7pcw47URCL4O
loGJMQ7OSqUOKy3aeq4Uny68wiBhwCBzayep2ehDG4D7ehImJ7AHXB42AQHb2Xks
A8daYLyWvXNpvLIZAcUsvpMpsP9oEGa2tZsv/ZPKnYfJrbRTWSoOOOubZquLLN/n
j1b94K5IZ+8y8s0Yf5es7jLOH1vbCpapDSfGn5/j7Pa4sUevIXznehFXP6ZwFz07
ZjzBm444siwSB1sR05/DoFgNgX+5p/2LsdnIaKuewD/gafBTLCO3cQE0JL9Dnzw/
RJhsN3WnXOfpWb4XI3Pf1APliJaxKXUrbwXJ/+fUSGEmp7waITbJWpoRYxhyQE6h
e0CcGz+fiwoL5ky8vp1TsP+hpG75NMMD3TGeTUo0OKrZ1voY73R1cES58EIp5y8c
Ddb1yE2FdvOy1B4E+tXQkavgaaDoWCMSgTFKQ0NTMyJFXb6tDnxM5E/mzCJrkTP1
AeXbJQjLt94+caVbsz5CCfFDLBU27nUb1Q0y83yFKS3FDgGX0cZaM4ATNyiTHhJ8
GkcQFcmpX6qzYrBUpv0+ZvDqGMgK3k+YQTQWZ4yrzJMELtTwe2CjjFZ6eG/jqr4t
7cmKUVryJZPSXAuV6/4wUv7Pit+m65EZ11cfEh9rdKq4PMfEqaVIKwuBC4yfLWKr
VqUxidpF2t5Ro4SQijnJkVRzmDOKoVHdT5KaKGcAvsny02E99gzgUDlgkiyTDfWz
PiNQv8cFMUQcCoVzl9JUT/CRqY24NICArpRVvsb8t4HfSUh3Q1EyBeu23aSEUI/P
cXDtd/aQk+Mgf079Cm6K/Oce6uKEmR+ZuoN6wvCkNV+BjdwPD4vijJnJ6he5LrzK
04VGzs1AprfnEM5dJ244bhP+m4JmECbS3ZOLaSEf6SlnF7r/f1l8LhthVOvP8Xgs
He5RhGyQIi+nuTpHWvipJmiC4eECbwip2jE8fZsfOlb5d0rGNDi0ph3m+XjPtgBo
g6wja5j+wUCmh//zRa3cCO36nSZaAIUmUHo6stgLhYWuDGHOEC0tNUFR1QsNZqMk
lILD3y6TQ+URAWsEHcjATOKWcKfcuY5BYH23LKM9467HAbmpaNLrIDDR1EZSToWe
+86vbwZ2jUOqhE2p3GGgTnxXu1/uW2j20Hu4SeArQBM8NuLhb8U6foePo461nw1L
EuJ8zWsa62H2o41WOY6HBzWiQbVh5r6TXv78FoBV7utZvtDV4crJK17xso8e9JCs
di3hTQIKMkigOOOM1tB5s2m/VwVlsCtpJ7NEOjl/yxIibWgFtFnEGYljHMzD50Z7
JFd+1HVUbum2o+q/SBBPUhbL8hL4DFR7oI8tTJ3HEttOqYFpwEB2osCAhYPwC7dt
bx5nA07fVxIEk8S/9lUvTpvawiKVtDpKq1EkI8CKJ+vzPARLo67lnIAsCzMjCYYw
oQyCqkJ/1BiwOHsZDQ4MBN/DUd+F9OTFUulzpJRW2vF4qUWe+3xLY5UOj9awQbsp
FeMojyJjQdeMj7jxBK095+cxBAGEsXH4JlxBG29kivhkdAzZPJo1XnUapQE+Lqn2
OfVjndphjcp07+/wGZuxb378JvgulaaNwy13iKGUdAaxgxVUxBxiD26psu6Qlp+5
qrlOhhFIAs38rC84jmOnMNurdGzqPgYisSRhg0KPReCLI6SXcW7XyCSotLA8An3c
OYIE0QhY4XxHFto1PZ/u9i7RzM8sJXsbFSMrMvri4Vqk+OARc67sYVicjIQHdxRd
KytmbBvhF7D8lf49hSzv9euzyNiMz8FLttv4mtWuwwByi3CmhIJJeH2WxVKfbghI
Gq/ek+vhC+OP2cThd6ypV3G4jxelun4jaU0QzUrk9Mo/6zd3LqE1z+lVLgI+YQlw
N8/14YT6R66I+KEsMnb6izbvileF8AZ6TqY2rR3Q2L2tQ9ZZd3pLnRkJ7vttate2
3G+eolJPGDAaTD7BSWFgtazNJzdTrpVCbjGCGpPYafQ9Ww3gXci2mHRvKpBy8kMa
vGx2AhCQIdWe0mzkJEmffUHOaWMG6FSrFgiM0yi0tE2QWeaac/TAGjLF7yYV2rO6
TCf/JwR28Du4TPiKHI4nJe+5T32LMjSW9/IBKhvLgpD8LQtupBtIZ6oOT6wMEoCN
JOgFGGBqwX8suIm9mdQPpkzfxD+5XiyjWnFpHZPgvz05H0Zi48yrCB2lHpwooImv
enMRl2AqbIzEt6nPUxGiFkyA7oYfq5LYaTSSYxG3QuZUg3mRAOe7Bo1CqhmOpiB8
7jKe9ILQvglEmk/V/dPKMSoPx6qaFyoxNSJSxw2i5usbORGMNI110ejTWauX3APS
EYQsVO17Vuakn+fW1hdBnmonNudWK4JSLXyBNfq5LDgTQaJQkIo+lpD1XzjiUaUh
N7kkB2PI6eGZQFAE3Trmv+3IZa2HSAhHvcjQMIToglkJc2H/gVg3xb7PGyq+ejX1
3zr8wOFlArQwByra6tDq9SJ0BT36XnZgPlLSH1LHTV3hL/4YtNO0ih4qqMMZ+6WQ
yN/bzAClR0KcPfdFKRX/te23027jI7+XMMYNvIbOJOom9of4Z7K/qUoqTUuT9C7f
4b0Po54xtEYtSjmMIDtiwfrd/vlbItaGA9HWXPB2dxRkHDOEP1YNmgCQbD4qEWlV
DeMf0OOBWyj4X69AXUWXfJtomcX6QlDulDVWp6GC+2iL/a5NT9Q0kGtWzip3+S65
v0m/CgMRGjiuBRRgQtpx8kKP73dPv7wOxGOe/dQL3hVIx3DCrlSu/LoI5Ap7x1zD
qIsr3NEidXmngJUMHNZGUKx0tq7xeQ5ae4rO0O2zCqSTGCJ0vJXBPxM4NeSqHl7y
vBvog57SXB4ipOESu+P+RTl/T8bZWwrOIX1R/aibVdSI6ZlKPYSPPdoHMVhCjdjZ
EWg9pBMsfroo3Olcr/hY4NJduDc+QQ0oZVzyMyAFhAyrzcvrbGjgNITLuIRB/diJ
osAqMGb0wv07V3sXbZxe1avwMy6tXMA5W7XJm/pNDUBUXUDiKWmRPBM0/gDimPdo
WWYYguqicZHtJl4XZS5k0MZe9PSPa1/hREZRK8BGiYoMu93SioxhUKfVAN99tFdM
tp29tKmd8Rk1st5MuvvKy+2MYhW9B4a8ViQiM2KkMmapSgkkvmvbUe33VCNDtUX2
WUHsZu+45A8uR8kqdzv1pgGbeR+t6cqCzzExwjMWlqP3uqm3KJ61wd+lkzAIQR8l
28sugtO9UIKnWRfYIxKdRQ+o8jMhWT/Q7s5n3Pvmm9EmRo7n080tXXHSxdaN8k6Y
GnaqzgeU2vbIjuayESTK4PxFxv2E+/gsFZupvvGsa1FxIG2ohOJ1ylyTxP/e+IgM
1IE5gedijpagMFvLG9MGoC8G2S67wyY/HdNszIlRqUHkkXnzCU2NLFRseAFHvvyD
NRCddmdHEleEwq6BipB2VoBPnYGXlT1VAJEnr854arN+NHC47Oic+6s51OrGaWb8
Nz/OczHUlyQNa9J9lZFoT6Ox9Qn8qEk0K/Tn61z/M98o95ltwE7E6mb2S1D+WHSo
Vd8vnSuI5eVPL3UxwzsesW8B58nZE2FwZxyUaSu4qGdIhN9moa4CH+7fSELZmzUl
n4s3a48BoPdfRTeG89/Br73ZwQLbsrxv2MxvNZLrCrIKGDbaqpKPKqHOHbG0mb1J
T7pKNmK5BV9b9c3KjIaqO/QLWZkmubNCdhrTQec2pMVR5VzPOnMKAZqPN4nR+ds5
iXfamexkPGApxUwsYwWht8w7ErMFviabG6Fh1niReszrJ6rbGlwKlTLmSHHiUuns
nF4HfYQkqlE7TKI+GArR07VSSfyvT3m0C3MoxSB8ix8RP3tblaI46rEDESPJNvr5
O5gXEdNh1Tiz4HWv0wJo7q777MCRGyZccz4uNLKjnvsMnciAj5PgteCgZRXlyV91
mstIdTRO9a5ItNg3kuhdnGv7hsmWhJtODouQq8DwBCLnu1mjtdhNuobXEAlxmZ/E
zNJX02z3zdNSdzQ0ieNUFEjuO7SZPbYyCukCZyzyV7Z8hwvvMvlHWoAe2C7JnfYa
IpcZKQngFpNp+DAhssnk0RAOwVG0+dIoSKgULAeGE5w=
`protect END_PROTECTED
