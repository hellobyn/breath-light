`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73Z+xZrSWrGZgMf5ADzleCUkyG5IDqQXQtOLtOlZAb0RMig4mIAOiGgi+w2zb7ba
DVUVtOfCH+2Ri+Nbbqxa1fh8BVCsQgz3fTxtt+6UbnsLXZUkrmKBedlReDYM8Bzc
Sad8oF7R60ZBEgAkCiqvN71C/M7V4sdG+DfWrFeCT4vomrF8F1+h+LDXazQW21Vv
7EWT63zNOhENgBrzcXFkbzT3u8NgEJFCw+5oMRd9W5BDMSVf+uksszKyNeE4zlpZ
LRJWVRNfqHT7+6e8uMEiKALNhnOOT53KtdKiNOb0EbkoYSXGkpU4hcynB4s1bruf
yVVmUDUhZsipc50mMpnrH6mPGrvScKSZyfVCC1MJZKx15tIxH+ecdC/v71JU+6rS
Dkwd6PZwzEawJ1q3k1TuvlzeVKWmvEGTU4MNbmsJABNrPMsh6dyJ6SuE50YjLQlI
yHIKCTuX5+XJ/jMWTtxfOudXJSU70bNTQR2M79U47wXfbGISVRG6vjVf4v8mUjwU
A4mJTyXrAB1l9RhbPCcv97ahQxCV/LnNAUbbntAj/er/qlUqz1vNKvALbaiCZLxy
k3ZJcQ4XvJC+YFYj5abpSttRA2AIm92P4gVZis3KxapNC+VHx8rY1K8nH0kbodZN
TKjOFND1nP++qtH1875p1x85K6F1SHgvvwpHkMbdEV0Gq76OcLkrg5LpY4Tp9dfs
kUS0uQkIssmySCDpCE55LiVI4dbs7jwhcJWEynlUXXtp8d4s0Zts7fOQgpS4HPuk
70hwWTPogMkgsgZhUOCUJ9eaq0YJAAJhSFkArAq6dBC8DDIq+XzRtHt0oy72sIIP
Ks7SD0ob17XwnG5uBGvnoNcnUG3AvhM93zUALTzJst0DDCm7LNEHqQerD/hLX2wW
ijk4/V0ibGialSzS9uMmVihiEiKXHKrMBK+O8CHwJr38gCdaxm2+sCXov7RRb15T
+8eCE6uSETd/UjtTBN/6/oJu7KDueW+DtMrmdF1C3tN4bMEmP8eLMQJzL4eMkptw
/TuD6Pb75z8d/H9CLb76rLFFFu1clvkVvP9mI1c8pCnhFjk+0jMSZs5VF+VOXn4g
fBoOGlgR0Yy5JVDq3hyaB0i851Xc/2rZ6aBigAx9bjNJUoFeQ8Yce1WBxPzd8UsX
pmmvxri3tfv26MDst3ioS+n8VlUZGlq+mroUXh2vVjolVkdvKZIanrmNntCU5rer
CHgytIQ4txZI8iAK2rl13cfMps8c0qHhFe/AxK499CAFy2zotzdTbES3UlhZJiwb
8F4WNEDeMpNbwj524Gj8YDGp5tjawh3Dbr4TWv3COUxgxQBjzkxFvPOPXJAB9hSb
ApMjzx7+NjkwBz6rJmNx+G8OmcuQ9LJmf7R0+fruDaeWCjvey58BhPSEP2mB99j0
wNQw/OftjZMSwEMiwBWk1rNALyZzkGvMUf+URLMfuWkqdtd5k62Vd2GHh/ar9gMI
OoyluysmzSbUohdblDCnge5/b+OWqsfK9aaQff8ljJufAT4N/TbO1KB0VaoEVXtV
PsWUH+dgge8matt3VEdVHZ4HjLKIEdDzvQoUWUAUq/BbG0o6eefMBjtfIp3bR+ui
boQb4VK2n7mc+95uZLEYgtFc+PRdqJHXB/fcfmaM4DVoMUCNGxe6R8snLcxBfwja
oyr2OVYrvnLusi1A5XUT4uM7nv6ZFF8hy3NrU3luyT953WlBsNHPUu3ZtTlSC24b
BlzIC9YFYfSiRz0leMSpx8pshIFrXtyxq4tbyyKYks8AykK0TSGBh80TZbi8sJIa
rY4M1tCwrlwt8H2aWqa/kg==
`protect END_PROTECTED
