`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLwqb5NWE/EZE2NHgYNCg6Y7wakpbcow2Wr2U2GqxfiO4+zVS0Nw/DSZfHHTSZcJ
rNqM3A307C1ZS7HX7FBK5wMRs8Cc2l+RxHR2uAOtJlTtpiY6MSxieDauw8dFZ5EI
nwrQyWRtkMczYrVZ2cleQv3/Int18MJvzGefa5Rgl6bzOFQ5+4ccYmFa3L3fmXlo
IktzVkMo+hfhPfklgqbAENBE5/917GuSkhiDykXjy1HDMLwSmPgsabmdaeD3NsLV
qZnukJ8dgd85u+SpHnjMF5hpzPcBr7y3tkQzlQ8dE9puuPpY8KIw3v6jGmCWL8Eo
u1EMueaD0UVDxKzTK0ICb1IOWlI8L6v/RHaCqtoe+Cj/nGqSAnG68hTmYozfn6PQ
TNzoJohU+7YRHx37hf+bWlF0hUFGciZzRkgJ2y1wJYWJ7Cspwmx/d5aPg7a28ZFp
I1brbCgKL/ZNef6LbK1vPo8rdWOum5mYF9FJjNMWe0e6fJJGaijTipk4x4RdMom6
OgoDfwedAZ+wiegZBoo+OYxA7EqxbDfOD5l0Q+cNQ9MM4SQowB8ZSdwM+38I/Fv4
expnkOpmqzjtqd6ApeUi6daBrASR4UYq+BcquVCfmR6wZJuh4CDLpiMBlgjlLo6x
ZPAXk5v51MdD01uf1F3uKfiOyMiBT5keGFx05UxkwUTKjzkMiprmlrf3l0Qv6iS2
a6UHqvymLrXAGDYnf/U6aRrug81Rduq4U8WHVWXB9ho2IjZOBvNF/NFdFn53WKrE
5xLyPCDtNaJejmnmQoBDx8MR2LlDBwxf/xdo3GRdkjanv4NbyPgYcijb4IXqd1Ke
gtrwUOr7pH2/sSgZrC3QGg==
`protect END_PROTECTED
