`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgjedwcFICRuqEKLqbeLc+wei1zuHgqJN1pHMN7Dc5NH5CMDii+cArggBgPyoQaB
h1l9SGWnLZlA1asDRgwsoJ64po+cK3VarM9XbXaUMJrOvEZUNW7cNcjkRiSpmIVw
bxRUZgutE/ucBlGpsBcAxT20K2mLNrFtIVYoMb/iRvdPuUlN3BsQ28NI5ae16r5O
+ZaToNXKA8xDu7btrNtlP/uIiCR9YvDzxBwvsvr4BJ9sjR9OuQw8Cod14arH02EZ
L8aiDRk3qlLinvt6XL5jJL0ttlCd0tSwQxoNRQLeHzwrOBBe9sLwfrEZDpkSvt+j
1YccbVWLqypq4w5BpTCMGjveOu1P5fOkIC0HUrhqA97LbXxYPnw4QKrZ7F52ECxz
GDhdXbdz1uRc2L0x2iy8W/OZ6POYbkcbPGSv7WmJ0vtvOkHACQeLXlmAub/rE1/3
s/Lou4ZAII85a6lOd3OPv5MWFWhLh8b8ZOcFsQ8FaS0g/9zWH+HNJ70AcW8Kalbc
k6FzIdfL410tvLSVVygsbXZK8RvhHmIjKG6bYn8R6OHVH6hpAFesxb+9ejKuHCSr
PVSTbS5NNI57NCoLmGdP4I/rMReplgQrDLxMqxraRMH4X69RqtA0l2Hyl/4OCOia
sKNEsrIRLVLXzcat9iERRcAmoiBEeKrs0UdJUY+QTL5tv/lmOPegbjRjIMLnTJAP
KyUPcmh3ZNyNQ7ksZ5o7fHuOsR8z5zX6fVYITDjaHxJlK+JS8i91xCgAD3gQsanH
nbnhdQjfgWf8N3mr/e0fLWqeQFL+8LuQVpIccpAVQrW+YGE6atjgc0cwmO1NO1Qe
nrGQkW1XTT9LbBnRLuY8EYCBfNwTF1B21JunRXOpaKv2xWnxap3HrNtnIziRholk
7f0dZ7V6O7obveUMLCYzjHy8GqEDhxm4qGwHgE8lZqNIz6WcHx57BLjjvOds/vFh
SmFrly5Ae0baSp8c8CJ08sqRa/K+3o3jwpSFoJJsfNMv6/4gaZl+JPVQ7D9/Gj0s
/IZFydRxgpEkPrDCNh2lgGLkurXleDg9R8V5/4yz6aNXUMafb4dy5PrWfAFxOzIH
nJet1mprtuwyTrwx9C4dyAXYjQdiC9CjB1FEIRMx+J2oDTZqt4EiWRx6/72hxWqZ
rcLbSVeeifeH7yMM6U5hFcjkKgWLsyfO/5DPMlsT68ivNsusiGpRF1d6e0KqJ53l
DNGlbUq4S6/1hIpGKemIvj1sAdlrOGp8q2wrJtdIjYpN4MhW1zuA2R8Lj3FgZfm+
0ciaVOVOpc13lXOqAIfJ8jDIs0PThJkq6ZgtTOODf35KsNqwuWGCt2p6PNWnDkXS
1zt9/SQJntmyDUHm2ocUuNQkOXuB+6dn0/kPxFJ1kCvlpPJRgw0AEw9k77U8s2F6
mooSFpQ1zS/zdreotdmYAwoxUoIYC5OGd7trSpu58Yx+SF9NH+WQyT6Ri05Yi+kE
QOEiGyl1YE3XyusiY22DAEOemn0evnjLVGoQ1aWaQBjvCd3Gw7/58ITyihtdW9S0
ODWU9lUB7HJ+hlYSoiPUbW4vvKc2Iq1q1dkii/7gnb5rj5t3vryl5Vb73ljqa3zZ
NA9oh59Emyq5kLc5pZhoyBfSAzkteG4ESdHCk9uST0tjVUtFv3iTWPnNpJyocHj+
yGGXOitSOevwKokHjeJVqNIN2s4bndmuqQrpdsMknTBwgwc3bbccwBmW9dFV1YYb
2jOD//jQOeHeST7q0IZ4p8O8WEovEpodCUkmBoXaQYUpCJ/Mx6v9jYY5seNpCFYA
ajELVJ9fB9fwg9WjLL7i+AsQxHwtpB0JtBlQUYVBFPsdeinU2eO8KCHFQ4Db6Cq8
QXIj6wQph4hCar/mkBEuMkIo4zkz+gzVTi4VdsGUQoOd2z8u86gNB3qD/Wr838He
BsmnDibFkMhtfB8tC7NExUkfODkxlhdaXY2JKAspK0oVoRbdaHycEKZbp5CyJQrz
+P0LDf6uVvXEl9UwmlEvn1nscQrKSHY1J40E757yNZJ70OOe5Ztu85sxX+5tFySI
SP9khy8sh/90tINzY9xtoSHm6K/2mtfd3c8wQOlgkTFOlXT253bGEQLmO7bZ57Il
Q+qfsTFvtvQT8ORX+E13NFzj8izBoTIN7nEZNS5Y2B10OdYxkgA4SqD8k3Jjolxs
iRgnxgy1NBIZX6DpJuvZ0MxmbeZum6EA3yTNpo33/topB6XBrsJTDq41QCxUG4qE
QOAO4keiZ+qJtqZaIQ/5r9h86hc/NUej5P+dzgrT/EacuiWxaDR4qkAoJ0v75jHQ
ddlSC0Us1b7oUggn63wIWuXYpRUYCc2IQ6/Lve8RhDiBzlsmw1soI0+e1i0Wpgl+
6g/6k0yUzTHxuLJyh1+PdEiFfWML9cA9UXhKtUswpf6P142SkVckhG9ny5Fok0NE
FeuRVCaDZIT5IYdBzmTdIah+ZnrYi6+kNBhkKHL+srmVjffY3mJq90a2LnBFCEWI
Crc82JeeYVj55d3mL1kTAEq5V2tjlCb1FS7ZTcKNMjuFvbrkMspK/vgybhq/O0Bl
qTkB0EC4NHz0xusLgECp4rgD3nR4tmpFL+duQSfFgpLD2kwg71ybVLCzjbY6oqpX
WPk94PLd5Z4JIjbGgQkpMErRvtHizWHuEy1eHojzQcqtZHM0JtPpUkyJkrZyDO7G
vnhIhm2BdaUWQzpAY6C+YZ/GLUlQ0kciIfJz4iuKFovJ4VjYvRM71ie/9PuO9z1c
+RQ8SOV31Quj/Bz/X0fIyhFZyunOvVEXGhN7CAGZpAG90wiQmFbCObB52OUGMVK1
XVpOKlC+iochoGSVIu+iMtTmkVowYfs3qF36ivLaNKL4lSYyvWdZmj2yJvNfB5BQ
qBBh4Xsbs9cBCayQXUHKHSpALh//1SjyqjLRD9ba4IJ+0C8TnonXai1lkfoNt79v
+nDOGiz8Xx1/uYJJaI7D7355bbQsO3VGqQuyHHu6vCvuzW55ViQc2FonN8T5WWYc
X/O3ZELGyJDEr3EZRWZRNfrRq78+sqPPIPGQlGaCU6ASulVnt6lp7OKlXdRwf5yx
ekrajbcNBqk1x6WBNA6hYoN0EtA42WM9rTKl57sMdMd8JaChsgaU9Gn4Z2oWy4Pa
DRFf95bGpmohY9ckpB/YioFfPE7RF6mjOGhBBWnUDIi74u3uAFncPPJJ/4CsNM00
HxTRv/4BFnUj2elNXVWvMvKjgMeq5JCvpZPvmrClb1LjwJeCWPrIrHsm9NcUv6DH
XQY9kVAuMsPaKRPDQGh+FFYFfzHa2/ZFS8buf+ABXsW6uJIzoheGEIE7ZFRfu/6b
9hEjz3Bf+oQQ35+yYRuCIF5Lax8W4ngSwmuDyjfayRnnx97nM/XoYqL0iLua5ZzU
OdIFo7p3R2ZWC/p3KqsqlQalk5SE1wy/Box/tnO3QHMLluchhycSfCSvNY7EBhK8
x+IDwql0jHCLZWVWq8401lBeyPCXH6kNI07l5RGB2dZL1JAksZhKAxcBgBycvCuf
/wPdq6pORdvMLCzrrFqHnTy1JAT37a46XandEaPMdgurOd/FOrPtgzcToYY0npvW
ZbsRtMMlNC0t7ipackeoyLQwkh4oIqqGk1edw3B8Jb3pEtkjbRLTdYhdDYwAJIq3
9gx6VzVwylTFAxCYm1iJo664LD2t16t2/7g1+Zc2iv7BfSTohvyOcMDg0Xh/Ao0k
ik8gIgWAz1NR1Oqepv5FGwmB1QgBZvgeH/blN58bMmgVG0hODJflhhhSMCLfK7vN
RDnwPoShpyQHjaxUl+i8b08CGNrVi6ZUx/7nt/kc7EA4pjWaTBe6psBZTT0lrT4f
CI3lrIPHXh4L4Fzn+xPVJjNz9cvYSlB8p401KMqSD3v0uHSTPoWd0k7jmW8XM05c
6z7xpJzik3/Z/GqTbMtuaZSBLSOQ//4cdMqZt3Ey/FRRZJDjVcEMvk3RBGV27oRq
fuXki1jiqK7X5SShzRFvhW1UxnQxiYEdtjJGBY3x5D4aQWVl4gPjEk8TCWU0n8xU
ZTKqguctoQ6cPOzvJg58HZpyZUZa1QZ5USedfAu2r2IKxWcv0UlQWC1xR4knILvk
XjKJV19OFbfvaJhdPUNlELnJ8g21bU8rVZLjxCanLQO6qSyNScgKhhUPoRB2LyFz
np/87hLINi/qeeryV/ZtdZLRot3SSX7I7VX726JuE1tgqlppr5aCFhmMCsA7OaTg
bZq+ta5ilJr/4OtA/NtJ6PaXUMIMdF46ZRq+6LSAoWCOB0CFr0YcXEx4dbtn1r/r
Wg0Vu9YM8LERPx/s6zeNy9ZLh4bwzwj2BwsZ8jSuXNviqzbaJ+XJTbLF/bepzbi+
wvtG5OKznEdH93jaEZ1YvRT4CD/TKiuLRWrqyXCfKGvvXDIRl9ic7boWw0kYtzV1
gADBda2VDv67jY65UW2nSJqmhrRLbJrqw9yBfhfQbK3E58qhUhuWRhWjN0He0kkC
qkc+/WI5vlQbAYoDKSffyv3eQUFcGPpBv5dxdrSYdXNZc7Ja+UA6bYFmBaQ3r90U
IzYvS6yVr7rN5kypGtitL165cF7pl5r37tzgsa65/KtOAJQja6CENmliOYms5hJZ
8H+Yx/ANw00eAVEdNvdDFJXJoHqNbiKvDnnHsXvkhBr/raTfGObwD8RN7Fb1WCSH
sEtLWyn48iAc0hmAqvrRKg0y/KUneUleqGrNxp1fVVo=
`protect END_PROTECTED
