`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNOhfd4Hls7jYe3+uq3U5iEj+K/BlEnJ6PncOVj0RBhVbaL5P63W+0Hy8tacXSD8
VuZDRPcg+81TxAwzSBDg3JEb2y/iccgVWo+kztH8LswNtVLq0hHzxfO8L/LIX3FX
bYSpWwki1M6InzCGzC8Z8jAeu0N9BSpMk/oi6YM0MMhHw5EbrTom5JBln31X9EVP
xHhfA9xbxM/mUVgCmsVQ5yALS4afgTOsGJo0L26MToAyr2RMNWQW0yTWvEQnsXm1
+d8n9X59YUm950WzDcAjwXvCALcaYsolkqoMoV791HyftKWU4vDT84HeBJe1mD7k
QHoduExDo5d/kNvOSw08VZO8/9Z0AHusbl07f8SMjjIugLeSYRIGtrEz8ceC0/Ch
nPqFGpn8vStyyLsZHOo8XuIb5LQ0F/ZGPrgZ6G9zU0V0Dz5j8kMfUhOroCnTSw3Y
Wg4y2UcnHgsuDFU0JMbBE38MsaEdamY0pY/ARQthCaEtkHywJ4YKMKG4bUJ+3BVb
ZTZDE4q9JXwwQk4WPxPVWPB/1kbbe0agzSExpkBQSFk=
`protect END_PROTECTED
