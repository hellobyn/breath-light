`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4cgUYVgzZJVSnNdd7XBRHKGoR8rloQDYK5IY2QoeoaD9KbniDP6wvSxVzaMHZ9C
q0TVFH4IT+GEEdxILjOArpIH3ykucs7/4kDvozqiZCRnKlCL5Y5O6aWc5CA2WnVC
YGAYwu2IqR5vHulEcYklDscf2DRC+vnGYsQ4S1N3AT5isW6IreZ8bYXcP0OmddJH
c0wERMlQW8l67c5GRHDeUGMQ2vuR7i50+AK7HJk7kqffLse5M+MmF3t35PghnfEc
GM2n2wc55TqR1GxZ+1QLBeglb7UKHkI6xkq5VAd52hWlzvgH4jHPaGYtILJevJyJ
hmflEIBlf1doS9OkAOvvBuJvo0QBBfTTs+34HT08mNZSuvFNcDySVGwkUu+8wPIy
LZQ8LmoGePL75XPHRsrtLV2HTYfB2fz+U5adBkKcJKaE6iaz8OA/Q26rY/MI+hgv
Boe0xWtYiuWwqBmC2AJQOcHwQ3QXG8tDjAGiZ9c0gr8k9IC90mDzILhFjVvWkbWv
8eet4afe/eBiG3jD7/ql/9dXFrtJ1Ms8GMk4d4AnCBS2Uf8H3usJt/J7+mpVqDt2
kouqntLdfSkGx6WE6BZEZKbkZ5aUYfGulEBH6FQXVvoEhiUGt0wzPG47RwEWGhOH
FiM4uTSKJwV7LK5TDBqX9j9kAttlzFskPzHwXFXn2mF0YEX3ZH/sJqt/m00EFCFU
FCg1uXlRupUU0kv2Hs4h3axZynuDkVtt9GHBX2nVndDCygl1Jr5xCOoikgwqLbsn
pkGY4bEdLOXDz4oPJ+BAutyVJP45wBFdd6SSawgxKZNCStYRU9wT5IZR4GTIejDP
irylqQSM222cxvsJlt4gzrJOJ0FMLWPzaigFJh0aUlBbcIghkExXYdOXlblgJ11u
rUAx1m81/wf14pm/ONMiHwVkixDzQ38H1ymVBFi0A++oNx5AnXHOB5Y4KBrSCeS8
Zfhkj+JLcOtL4YCbS8Prrf9CtuvqZk5bRT0fyQHfQAh4ElRwvqVWMNCNj9/QYm+t
IsnuVRjW6ClmZjcBu9MCnSHW+wdXjWHbzTFpoC6MYjmOgJtMArPRmvlg2aFWYfEa
ht46fm4aRO3gIzhyFvnHAjtgD48YW94xRyIYj+ksiY9aPYNIrDf/e8GPG0q8sl06
S8gHpeTNM5yEjjTIRknMVTnB4zXpp5kHuGc5JNNy4dkI4czdLPdl0fL+mB4sJTOA
N0EtdLc21smmMUAoLYWqjKJGvCP2VxUtDWeglSSFWiDQ7ahIqgR4DJQJr34RpFaV
ey8gxVGWVnp8UghbyQJ7uO0XdgzG2NLvOKrhqy7T6Bt2QYBbXftEbQ9CBpnlUfjT
KPRuR8mm26H4k0k4Z9XbWOOSYISPrD0HfLGSJUSe0ds=
`protect END_PROTECTED
