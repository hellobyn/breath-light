`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bL0V85ojc7Rao/J3iR2TsQhJpq32PHtH3OYXwZtxm6CeqwYkNhEB6sSnfUm2Amd5
TADSACC3mgqO3Dv1Ldi9gJPu8zMztoJ4XIlUmqP7RM9fePbalidx5wMYa66ZNiK7
wc4TRQDsUQJPNZgyLDCWbRU4GlopuCJHtaYg/CR8GNvlSmV4wCG7XwWvZEkE+NtN
ykbSMDulnDkxU5msibt0alvcI/bC1erjPbkmx5uJIz+O9mAydH6AmUHWdfd/Oq+Q
XP558/1E7jNUu/iobmxYXF1fD+P5QUL5Mc55D6RQbu27XvQXO5nITompAYZbeBVG
osRemCz8l3kCJoYb3hU6JeDkO3sITKpRUQ7wnGKECdkjT4ozzSu669+E8wBHZEte
0qix7tyi6sdQM0ehxV0nMTR839agX55jdHTZN87lULRIw2UKNKa4drZ34qgfRTmP
dirb1bNiOP1Sq2N8lOIjhU1cL6uzLAbF8X4Hpm9ZxanixCSI56Ncklejz13tGdBH
wtEjdG9opsEDWGL+6Q+GP2kz1TX0VzdnPA766HnMKTFmeP7Z7y1h/LZQxJUgV4rQ
bwJ78tKe2yYJ6imGyZX0qmCldSA9z8iX7zB3l4vOcFRb6kTAClOrzZwETx6DfuHe
6QR3ridNTTD6raITknhaIq1Z1PVR0wneOCCj4fT41Odn80FWKYZVhiWDiNzvZ42w
U5r8s51RayFrpTnb5JKawNQvHcpBlS/EM4TD5m6hfv9ikges8BhcBQg5D/ZWfiLo
rYZUqFfcrEEWahxed7RtkN7Y/xO3YYzMFgBTIsboMb8Ra1R7Kx1rsAV0Y+tWLu4v
TV08fLRq0jpBVN497PKrb4Bo0wbBil7JLZ1cd94vjAKcHNQKjHnxHFkFslw2oOCO
TAenvTvo7/GDjnzfGrYeu08Wa1Rz4SW7Z15Xjh2EGqHadz2T3A5kiKm/PMgx4ZXF
qnG6J2xNLjVoPZpybPKh1fJ1JNkPKGWrcV9KYETl3fExJ5VguAyDy1Fy4txCwv4m
HWLBeMkXogJt/jV1lJaQcaPVR2hzaVUhNKqW/PYo2E37Qz3xBYjnrghB4uK0Gzmm
iEccnrzGaZaMl0/Mj8zrW1OPv+lj+QJQ8TEcU3KHsFZzliLbpQkmh6yoX9iCLKlR
RHpYed0zNeCOHo0tB6S7nzABaMcTJm0b7dong052AAIJqhm/LUCoqbvWNyeUKHcl
pG5fE1rIdifuzmdbWJFTnpQMlZZgUrgKc3DLMrFK4Eo579T3tEs7e070hgIK83z1
rYvtgZibiZOHecI+3HOhZdDauBxngp2akCTrTo5z0Ca0QaQ2RcCDmh26E2E/YbvC
/eFKUPG500xR72wUKTY8IwASEAv4dCnbmbVJS8BKgiUb/7bXiH3PPxJjOiApjgLZ
27T2WWQUJCZqiR9tILINeG/20bbC5oPylIB0RKdOoD7cL9d5hz5XmJDJ5khl/9Gw
sRGUM/DviEukX5gRxl+AMD0HZd7mq/5O784RBjsNIG2bT2GO2WfU9C5dPP4mt1d8
MQxSCzL4PbET5byWRxXiLIawNSE9nOTOiAV6kXds3H0Iuw+ScnQBct/O+Sr7SqFv
oFKcy96r2n39Fu7oOh5lciKVeZ6zW3zfeDzR5Akjy+GwJkEHhhsKICFVdk1upiaV
+BPF6CJZzq6Oh0I2Qa/ANMLMRKijQzg00JfBJqHtixHtZubUe3EXEKS7KZMzNwAu
o49y1+CYz9n0DDesLwQhOq59Bg5YWsMwgEprARK0MxBFo321ow9SguN2xr9mXpeH
GyddSWJpkeJqTldEDe3CI4xKjhMpDJN+7bPgbAV5QTLUsPv+MRp19PnIdoI8dWSK
lf3wLqWWAMkk2vf1g2VQEVHjp4ErEOO4QV8MaGuhwfobqpgVLNjj9LydfkQFOES6
9F3RjEUouipwYQhroqaLutoigFY+3m2jDMkp7yIKvDXiw+sKmHAcvNbng2CmA4VF
JjrYL1s9OFaUge35rkhtEnsbb4YEvjxtXSFXNNutdrwtQIFEOQu2p7Pa5At8DNQG
coUFZ2Y+Y0PtylG64EZGWuqkEqgepcYdIG1lwHQd9Dw+mZbMou3/GtZrU8loVDb0
UX3yllvqenveiMKZa6f0hkr0EehESTPKRGEateqF8Pz7x+/AsIFGIDT7CF2nK+VT
xhyWXkGGA1Ek/uv1/9750Q1Mf/aCQdGOE5jdc8BDToFZlf27Sopi7OScnjnTp8Q6
IUw5Xl+xuAQPclcelF3rnP/3Uf9MOSwWILyOz81zrEczZBeh2buNzoIoSm7Y90J7
xDQYiHWOu4eOtAGkgsPAQ9zY9LoZAJnsU9gF6T8y7i7iPRCE2G9FWIzeExWXLdiP
OgMIHbcMBTxxgwnSnVcAnPL92e9KNqPsXXI4InJNh5cshwPmlJA9XvD87r938G1A
W8IQlaOWsNZyE2qJv3jdIsY5KokIKtkx+2h4PY9xeWPWKhl05QCsGfQDbxmGKBLQ
+/96925/0IzNmJZqAzx/uEAdbkjUV6XYf1b8SSgBRm7qnxDg3TVBkbQav+3JxeY8
S3xidMwhOYnQS5xJHOI1LeH7GKNGDUU0LMEOmoq5vjcaWCmPXGkgldeAnQ9F4Blu
V0hbirEkjylnEA8tLERXLQ==
`protect END_PROTECTED
