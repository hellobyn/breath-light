`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eOvHn7DwJKWCaDUCWRXBSuBUf9DiIwob/JSWoXgmeFTLHrupbv/go+PNmtYovmty
b2vj26a9watv4F7k1oiNNSUZAPRKp51Scmsf3lvpA9SFFyvb9EtCC4y2O+xlvgbv
isdUMKeen41fNwxu1ic/3N2gKTQXnFxNPaW2NzVJ16DJ/9ZygwMzvZfTCaPWhIVf
Z+NYJh6uNQJ65Ir0MQoCLzNiLesTBx8L4H6pt3gsiF3YZXaMR528X/w7Mba3amfp
gFiou2tn1TorI2uFxJyTHeH5MmMnHqFFnPrQy+EFl6XCnIbCOIK1s6cQF9uJn9Us
0XfALvEE/+L7Bn9fE7zFxD0J/P59X+tsqkUT/xcZCUONuu0HpRMTKqyNlv6ja/Jv
1qkC+4Xzm6nsuHEUOfpmpJlkeTchRpCNsy89X3n0A1COhWic8MGnMzfma9RmcdUk
HdQ36yBYvJ6U/Gs0/606cQ==
`protect END_PROTECTED
