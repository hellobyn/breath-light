`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Abx0LKCCnEHHHO84m2dVam0cDbLxTrf5/hz++Nb2hdMkzR29oXVj6syLevN1J7Cd
gK2ARFoI12fvnxpOFZavrj9FcwkzUJOZWg22+E0Q07jYgqIphB3y2b36SJPZaO7O
4tK0TeNXhggnA7DtpfwLyhdyvn1cucOXma/dVjx5yM1d8khuGDmM8ZD83Rqpz765
dwP0sq6Lh7YfkJMsYu2z4kGyCAIVfhsYfoPuhlh0w8aBGqOpICdGPmPQqh1ga/y7
gEazmpVah5V8qZDyVVdK4Wh2u8S2bgbD5sX3L7jjljdCX4jDj595g8/PytI/CmhJ
2OIviz8LEU4L+c8iw0J7KSnmHhhHforfjSTJtX7yizuXkaGkptAGKZd8JbvJGGWd
G4JmVi9iK7B5ObUDIPUge6Rlw4BVtFZSkQ02grhD0y9QJhbA+AT4uka/jtJwMstb
I3dfLg6BWsfwPNhhXZMPZfPPfGnw5aBK+KfbK++XZNfIQ7j5Wd//clWOYb5tNTCA
Lz2MJwrEbpS26OMqrbk4rNW0B5tFL1DF7d9KYBepL7Io940AMKP4QnE0h023h1S0
ED01ko898EK9rpVsRLKEXMmfQVmZFpfIfn7GRvZegnyzWiD0ifHxMZ8b0uoYbcjh
OG35ZjTzWzkzqqeHEQPANAr60bQyIDXQ0Lw16KPjcPQGQEn+d5n2K1nQNNANIHHA
T7TyTFfUthm20oqaKhAKvHQ8DaswS9tXGRMx7aYVzLqceU4wC/Ulgr2+2WWMH4rs
wwJDe0B5t1/LsoibJY7hZFTFq86a0N6DUSjcbj1ddrwLrskYL85IzHuXAyH7gz7a
SPk6z6fVgA0Tf8LNidqN5IgTfLYdFrUWgfQSDFnW2AuI1g8MbKLTUuDPkKesyZX9
c6TutL2qyoupiU+10/VBmLkF+x9EnalYFa7zcG8S4NBE3dlq0gjYn7xrZ/FnGZ3q
RQTXAtpTDmU0uAlGLNyI23igFovNCl+M0BiLLclJidqX4tKYS5c/IOc24rqikCXc
VBBZ1525rVTxyHRGxTIXUTXRVYH5D9pcEhvx/qT1TGdtmekGy+XpjouerQWJ6ywt
zydeH6gqfRp6VzPtnVisWcc39vJrZGUT1Sadi0drI4Bsycbn31UNjPSlOhezQMxK
izyOQM4ksw5yPvQ0jx9btiU/RSr1rY/wQg+d9yc2Yj6VidwhEO9F6i0V92e9RLpM
BE89Y+8C1dSeFEUbL/EJdwpW9r9Fb9s/LTmMfW8obhs3Sfnt8aQ5lQ13u35tOVY+
sazTT6E11dQTqnUFQfcdwFsiX1b8cWNDHP42/E9CZOp/0Tr7eab5zcHEd9wO5jH6
c9/GJh58eodCL+4BenuDVwYSrSD/jL+QtpgaMDCwqYfaXfEgihr3OZBLiHN+ocMB
Wx1Dq4Aj3bOll9oShsxwWbg9+qR4FyPCzmXY8iginS9TSP3zqaWQVQGQH2cqslwp
UnjI6icksj7NHtQquLkd0mcdbFEewTDfiwbvcZH1fGjEPZckpSjuqVX9h4C5WTdc
S7/gDlgOuFa+bTEeWwKLSic4+L2OaMJLCajyuVYGpF48DDciAkup/rt14wq1/MPZ
cEzQQOT3oidOBE3tf2OAx4tIb5GchSw+MsUPD+RPX8slHqQAvvB4Gb7h/cLb26ue
VcnJqy2URTfpXpmFBYCOddFcfxYe2tFHD8hoDwWJXm9kl5+9d/xiDkHniG8qnk7L
lGJJ8d7J4VVIeo2GEx8Lh3H/EAQzmNbEzLVXONKqEaNV64crvdEkMpBWQiD89npV
E1MPXLB4RTK9ah8uc/cIzV7h9pXAxO6Te4bZ5zEWB4Glh0zzqRzeFMRXZW1nj/VF
fljmrrJILrnbui/oso9aWg==
`protect END_PROTECTED
