`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yKuC5gErv+BE5t5zBxjeph93tzdgKns3IRXMx8dYGgvWf6xKv1AY1e+95R9nVVig
0/BiabWvcceA+sif2sDPZa3Bq0ZN4nYqCENvx1FyTV9bU7U3hYl8ZKIwfCK8WILf
Oo//mw27PPFOhAns3lbH3/QMHA7cubnu0FtBAbdpVqNXzhuj3yFM0bRytG04wDB8
aYy29A/Ev+F6n3dcSOXRy//jMyVhSV5PO8wp9SnbLFyXTNbD2kr/BbWDFbx93zNY
Hd1Vwm68qw4yUvSFGZLU9MJ2wyHOMaf6qEq6zEgXpYKL+95I+YMIp/1naAlMUZND
d27d69ADsQUlmbR3pzZYuLYljR/dbei1s9t+20H+2n0ogq+XSa2gFhu6mvRjKbXb
OJZ/nLmmGfktU4RaWlSIcNKDfZT92C3UyxDx5mQ2lj2oPsb9qiTt0Smf5hGx2sli
Mky3egglCVyq1nUif6L3sGtebCA7RON0f0qWbLrE1doSgCVrdyTMb4IsJpKueqtk
abHlwGYkZnypXfs+OBGWD2qYivumr2WYXD1fAE6NILmgqHKj21jl00fJR5bVE2/S
JDUyEkbJx+w2OBPEwJvO1IU9OmHAtBa8a+ovvtIv8jcQBzW20N0cSZVK4mmWsKXN
ZbRbFMUGGypOi5k0hyRsjN+KrzpnkVtaH3cO92XKF5K4S+TtHEFST6cinGcys/By
MpAkovote29eFewBUKHCDkykdICHm0ddICXb0g43UX7CwOUw/CjdR4ZBlHAZOXSr
0KzmV8YkcAjNp+4qzai2sCeq6mxStmENGMe+e5F/V0Ps21EGHMxCD9lanD38Us0O
KeR/jGZDE1OyQ7OWkAtQfqxDnWv7Sd5u4SZbQ5y5q31uM7/ah6rDneR5vGNIhejk
CIZUFTr4oECUAgLPAFhv5vkI8uZmAn/VgZXxTbyrbN5zcJIAXt50hJsoNJAEdTNP
Rzj1/OEJXOHeTwRUE7mZvD3XIeQuzA/P1eGswoR78uNSnyuisRswIqXDf4u6/sCG
zcFy/nLh24yRDB/zilpYz+OThwNfQLxQ0Dl5y0L3QMYTYQy8veFczc1UEuT/ugmG
`protect END_PROTECTED
