`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUT9vPjUoD9llUTu3SIUmGcQttCd2MkYHg2c8MuznqzDvfxob9/+XZlxrnF/Rq/l
J5r70o1Re0HkrWLFPWYkORNRLnziyZKQh1OhHYG3OPqqEVeKgIyKtVdTgY8Ktwkz
ZLkudK8cIt6zfG8KFhvWWZPlyoKTr10qMtITK62B4f3S1IVMg6wYULxWmFmrTkOG
0BJJ+d3SSe+dTIPEDmDMN65S/mAsyzk3J7mJAH87BNcL6Ixbj40Jdy6TDWDyqfUk
9lM04rmrYwxX2AJPCaGLH5XQaZnMlBcKhdY2AKcMQVFdPVliywDnDWU8pKhaNumu
LOa9DUhojsn3432P0vtjgi7lqtC3PTeyWYArHjfCU7hj5jj7vwBFM4AQT1yyJ0X4
poM3CRD9u+1p7TzrMylXcOCdCEZ3On1j/OopO0zWVZMtZBdU3OlnicgBTqZtEKCB
rkzVnOuTozpWyvP74pBNVhilIrxC/KDleJtYyMk9cWJMBh42Bi8PmnKLPa5eMnjc
yB0prENBWa244j37zEGLz3akgtvgW6NXU4tJKL7ixJQwiP3JD/78rE28HtTnxtit
XVn5sUtxrB0A2a6ShiU7s3/AcJna1WKIcvllYPGQn9VUHfC5bvFG/rOXSs5XhXK9
9hJrVn5Mj2uUKSN8P05UWm9EukLICxXg7K0lsUHfGSq5AXN6p2q+ubnE8OJDLU7t
6HbtlvIxpFhp/+7PWZMqlpxbod532pHNdlIbwgXn8H4nr8tGxJEl4OY5MiHfoiKz
6vOvbJshvBM3JFIgIzYRdTTnH5jeeSkAb0j6uT/yL8DYxewCx+Vwd8DBoe5WQ4DN
jMx+Nh7axRB8ta3H1J74PBk3jPu4KEdKw6K4VWqHKRGtm7KFbhO8VWbr230flekW
mCABhg92gqRZo5rJQTVlos2qLFqUAgCm5IrS6WLlUso=
`protect END_PROTECTED
