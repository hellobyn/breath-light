`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xpqd4s5TiPIRi95Ks8iCO13w3eGULDRzBOzAbJUaUheemPvv6AHFOt0CFqVPz39z
hQkNSgCRcfUorCnEonX/5jD6VMBPvdjWTUWOppe+9Tq1YRivvYTCDLvc54oith5A
eRmgydh6HHcNo0MEc4LiJiZ28jYDVR8yiBtS5NeDIlDQTa2ryPAtOwRlMIihjDXt
77BKDajafpJbtzgtfPio96W1v0e9YuFvdjGtH47geWDvLmrqaQ+tJfBiTRvfZZm7
fNODOT95NBzYaKz3/Q5rW0pzxaKOIMM2VYOSKGHoVvJZnTXPjCFFmoJn14G2vaGd
8bIxkdAP7mBl1QbsX9KYw/iuBcOp2+/Mb/vevt4q/qOtxef645S3fu8m89MuLY0D
wKDhXNj6fq9oU+SNxGDMWlRIi841MD/wmRBDD52z95J8POC/yNFdd34vehP0TIl4
etkIr/ZOaeWvnvhYMS3FshiorOc0gEiBq2xXRdmpHNW4z2YaxeQDQgg/aj15ChH3
74gZJsUtaZul5lqu5QoiW953S8U6i858KRRbsgXCM8VFD4cPB2Ml8ZljJcy0ffEq
9QZXFQ+vtZPo1dD2Veffpp/I+bcmbdXRPLGa0Wlg6BJCkTLgufBZYurWHkvU5T6W
XNiZxTCzfRA/EP4stJmCZRERUEie77n+4u8hhgf7xVKGbL5zyZ3LOi7l7sG29qr7
MyAh4iRiQjAoY7pCEGTaUhUhOdYchzmOO1b4MIlKXU9odSCLrqjswIETEyQB/fOA
Mlb0eYgkQ1KK+EYJkdoX4yfNO+vocOfs2enBrtjrZ2q9kwHhighIGejf7t5DsU3Z
HbT/CVrobzEjj6Ni8ZvfEHZg7efMHd5/UfiDmSskgN7ss8rlmL1dnufwyJFjeeId
qO3RqB0gvk1YzpVc9MaXIqFu+imPpPXf4YLqIkQnvuNU02HANX8uLokojrMUQZUg
Kfxqackfw8XbSw/OWXxwZ3yauqbP4O3Zm62wdZW6S8EqzgKdNauyJjg8Nrt5ywoK
TzTabrbzgY2WzT9oWzLRds7KlmVbsh4WVRisjYQGw2ktk110UNJrFgjr6isrOIU/
vvG2sv3BNj+DCzV8DNary4Wxaxz47GWmgTVJXXIqwWz9D2ppLp2bPHJThBIIpvRQ
xAirQ45WhYRd4f7h3OEKp0pilfyO+UJljWA9uaI4VvaqwQD03lcyn3EUBvsAeTqc
`protect END_PROTECTED
