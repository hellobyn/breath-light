`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/wHc97e2d7j5vH2bOlCNfI0z+N8MU/GSXnxFdMpjWmZ8YleTLJiLFDNUy0Y6DvB/
ENVk/cZ/q1qDkBA2M2C0eHnyju8Fy2ax3rrEkWS5nq9NvV7RrG4wn64pKh6qElHe
zBiixGR5pflyRazR4TVW8rZ7jwfs73ACQJEAoLsACiajMfQfUYe9H2tZdnrs7D3u
ORfhrxINh3wu5JX3cqKxOuZDX/evOqadiFOszdKE3W9+7+feT+8UEWE/0XZplVjt
epSzZPXGPTrxVqpuKg4fGVbZ2kC1NRFpNsBJk3t1bivFS+utDm/+BdNTR6UlzoHV
eY6YtDos27D1IZ/NAaLHiHRfUaIwnoda76YgMQsDP+gWCfA0sbPNQFoCtC4KHWgU
9qom2n/9S3QWYbVKSXsvP1TrHiu9xZ05fGTxmuo1vurH+8PZy2Hu3NnAugW3WwLV
iSzQp1n6rHdJdjdk5DxsLLPfSrgStZsxbnfJdCzogs88mN3zuxzMf95KMsSL0vUa
kTdFEc21bXGVtfSzTXX9kLTaL7IPjPCJuc/BenfqMLYBZzfBGGaQ+JUm8+caoYNz
K5CRvjECEFsQyaHHA2li08eAQcpukwpQDrzcSzw7CHF5z3R0t1ssdI3kEwG4Y5F6
GbtHsXu6fuVJscKwybCo4rBKzxFSiVqmUq9TP6wTwFMiJpMtkdRFYjfuV1RvkYN/
WcqsIGkMsUvuf3pt3gwMSerG+C19rXbp8CBGAkVG9LoTry6tWKg3Eazkddalu958
qQj4+33Zh2D7ON1GmAACXAdZGD5y9wCF7eOKZC6sI3tulgOtpCbq8qIrPr31umdF
To82U3jWR0HzDZrnS5mzi0Id/z20S/moNMMIiJ5QKY3/yJu6NrorCm/LzkpuNQTe
viGQW9CIlMF4sDG1KIjj1OJSK2BiH59ppq5qd2mgCXeZ/T5EvgSn7qgqpmYTk2cR
dfFKZr8E909TFcZXuxIPxFKDrrvZmvisnhadvPtSOmaH9tZamdbYLJHwooDW6nXm
gqZyC7gH36IFLn7SdMsvQNrFVaxJ/uIRePyRis/ivzBu3lHBvU/MxO+7gaVjVS9O
4209hQOklvkQS0gYJWTmGAs9iehYEhshEefPqnaaajqYZuyl1k2svx1RJN8mhlNV
CRoMHssSL6YqnWdGLp/TbD0RpnKJUDwaX7Opj3voQbxM81M58Ilt5qjrChLc5zhg
HTe6vqH6afw217933LNXqevtHyPd3osP07mw0yyo1I/ipta73LmBPX32cRbEf+mu
4penDX3V5X9HMO1ey90fM73QvpQTTIFE4SSeU18gETQU5MXuCw3uBiT9ebZwIlsl
tkWHR02ye1qRu8MQNoZENEShjcexcBfF9B2bHYNt1MSoUZQJg0uy8dx6Mag6GPBG
eKcSKNAJiu/wD2pqE4Idwika5OHxP8vBsRE+NCQd5mCbYTJHqn40uqg+lZ2EJu/A
9tWLO/dHgpl8QYUTofbxXETYDqjzyeBmLT1JOgCSVrl6as28/muX+Q6V1bdHH1H0
584sLlkeS1ggRLgFGizhW6zY/Yc7e8WD+Tw6G89lRkmTC3XHQXiOqAQSN3LTiNxo
5naAO6EL+ypoMbgIs3kosMB7GT9v8Fw7qlpVAjPFcX93i2+WkNnMPQRMeFANWHk/
UIahdo8tLDz5VDriEfOl8V1P3LtzSdCo7KW8tgMpskWzvvXEF/iblX6JpzsMVps7
hEbsDIhICNyFJ8Wgi97MUSGEUFZEntiqvtS7fu+BASkM4m22wqtP7jtE9jsMkr1i
4d3voQy5nfvLIgSO8yTpKkytnmkxoJGX1R8Urc+vR4f2X6Kj2Hpd5HgIHsCaCGkH
9nyfDlpfVZxudj+6ex1DgtSnMnz+ynMM6wvZ67/6rCwITVToHWbcHoK+lZIwJfJA
wWirBCnoQHpEPr81PE5Y9upj4aTa0TSADyvNGspww3N7G85bF4pjgYWYzIQol04Y
bEmfG/BCBQhemR5F4WHrxny4o8OqjAnyTQyOX2/Nkt+i14uKKhYEVPeni5/7KWBS
ONA+wYS5LCNRBYLC7+DGJ5wkaHbkqY3gaTR3578MTnmQDEi6SUYEa8FkwgM4CwrQ
Aabti6JR9MGn2mMDDdL/I6W2Brb0SoXrwFeHo4UMu1jBnLNTE+bjxuXWy+FrzAlv
sM9QtAJlH+15tQ/PSBNCBBI8FpXA/f+Xv5NDtOovhCaRWNEZ7k/DNfx+LL2g3hxP
GvEWL6p/6EK9/ktbmdOMZqRdWl91RBf3NZQHUz3u22tfdHLI53f+QroBdE8LtwgP
+qq6pJkiD9zrqG6a7efPCkQzqlSyYudnu26QNM1NxX/2HByBhsFdmMiGn1/Ax1Pq
vyUiFJbrRQ2s2sE/l8emp4Y5kS9hST/RpPZV86GZ5GQGS9ip66W9fEzZK8ahKiCa
bv9WUSWNwmHeLFVDh+NgsZj4loOLd2sRhhiK8gfryFj9sBRfZ000vCo8agnW+j4D
RWC6J88fdPy3/Yx/dijRGJ3+a4i+uADOgQZCIlcty3VQmbemniG08AYSqMcq4ND0
rsEF3aLWmDFjdyIPtbMJzUCJ8ziV/eLv6Ku9i0mrSy9ieE4MFoqAXe/rIsYBhfFc
upcNqqQZoVcBt3tdNNURcE7jDtuKSQGbX+zQQrbxyTmM8hhJsP5GPhh1WZHfgWdU
V6HKsOcDZJNsUiKhRrzkIHGBr/yZV/gFwTYnrCIZqW/lWix7z0HWZGAH2LqquKhH
hNdkhYXTqLIusx965n1NyHeuzSw0vwawWKvczWMyeyn14cjtSKM4RpKRhRKhuAHm
NE8OZlOXc3wPYcONJuzO4BeAWx81LBBxKiuCPEPyFEF0NUM2849TrB9YYonHhQa2
ryHoqmXdhowcOkghfZYSjJ2U/3VyEfpD4c8QWn07XdGOdNICg1eumJO6yXRuk3Ge
XmcX+6qXUhI7ZAYd4f5hUz9ePoyPbfgiJWU4L6224gnAQIdOaYJY/dCZnWf40HTb
Sf7qnGC3ZIe+iK3sHGGT6T0rtyPp5Fi+MfFZMWqCnERK8RP4qYSkv3ouq9Smlrrf
XO4fNjJupuH6qSussqdvB4yDcrnsCFpYZL0UTRB+w56RuX65hAsEKcQdvBjSuUEy
G9le8mBhW26o5H7PBH93d2+ezP8SN6ZqN2hXFq8ft3jVLzVPEkM04xdLRM5MC16q
A4R/HZVzyGaNpvyN3+qVafJeKzsJiviM0ed9MrxAB3q0gxJVjF/Jre8+xbaEwXLL
UxPnNUFk5+cOlU1YFCiWy+/x4t9DHXZtEXkBPWJ+aeMU/YA7YVprBDJ/Sl2zx+YX
BvCXTb7vtqHEixlk6OOHlXRINQMy9ZTPTwoBfHL967S53anf4Llt+FwQcEuLCvfq
/dyKdJH4nF4xLkbLfnVbkC6bq+s6OgT8HjIZoysF81p+579/W93AdUEmZ365b9cI
+ByJkqPnjXWwR2g4kD/hEdU3Gh8M9ucJxTf7lm0Q5ksI5hnWtVZfMaRPmD2ZoW1f
FlLfkzb9Uarw05qyJ4gd347sox27DaGvjqBahbNeufXnEU5su+0TDnvUg9bXV0k5
owxYKoQI+6o0Qkc0a9Ojp/1Jk/TqM/ZGSj5cHA/Xf01rUK3eMSvfadK9k0uLyeXS
wztmBnzIUZup9fXn1efDhbD2XjPfyy0AQynQocpaGoPXb8BNpsajx2N642lz7Ny6
WTUbE0TLldytIy8Z9X2x0n1PEhavjZaUpiReXJrzpIn9zPaHlVoX3tmEKTUibOKj
nv5ToIj2pefAfrNJG0NmEsBQmCw113241W8sBMyk1QCpoXpKRqaW4w1p+j8b1p35
KW56gIDhiu5Mh15NqbGDv6yxvOjoiJx3MPUT5iHo56XNXN+ZhAndIGsvNFBcmta7
A9B1C95pV/VsWj6NV+8mioAuueNWU1wikrvCCeLAOqeKhgxzYmC2zsROOEgN56GB
/kUdk/5wZKdGb28K1taGI7DogjtXFUPSWmIOTxz/V1QyVKp5ESUsgbcRohIWUHlA
Apkui6K6pEjUpNHKmT00adRbmcok9yDprAw1bEff0PPkeYMgzi3COROvIaFoGyGr
8ASxedEYXdsDWEsm3+e3vZ+YLqw40b6cw6vSPGYZ0swSp1jiQCOmpC6mSRXK0bua
akMIJc72F9XBMWN6ZxxlGMqhSiEy5b9zDxZH9f+1ET442D1Mh3/p9dlZc2Z/jFCX
Fya1OQjmmbWTmDRb1jnu6IUmayFxa1wBftXAkbcbkh38Vs+/tQNAheE8YlSJ2GT/
pwZ50fzhTk28DgTxjSFcj2hcukJcRuVn46oqHLMCcP58P1/y1/LROnjHQOch0Z7Q
jeEPv647n0p7TCIJiMq4+4yiB6KIYbx4RY1qS20QmWf1t8dukrLmsMsL2pYQ+Pez
6jHawn/d6ENF+eoDVc51bF3oIWbtAfc48txrmvVlSZsZIuOfECpwumVHuZYC9Ykn
/nk1ZF5hHt10gPiHdKojAd1dIKqYh6XWcGLbRe+r8w9nFXTeduLcp3QyHoK30wdY
B+TN+eR48k+942tCm0ioF0tGIG/swj7iF8XRn31M3XQHnm78LXqJK1sqjDcyOGJo
ulZ8+76rmvJrB9sgJPM077z8sLJ2gTF+CJn2HwTcv+ym2F/nOPsPhJcEJNfCJ4de
7dWAHUeybZMEMN2qMyd8MIz83yCSRyH7/od1NFnZjhL63+s+UYIDyqeMnko4sgwp
cNrpCWxnCwbcrAGh4923eifySku/CNQxdaQIq/gV/jIdH8KSoKJO4J+oP0azyrM4
ii0r5+3V6zb/ryX5K3R+zCXBK/CcTG+HRkYmv8VQES/XhOiBlaAfPAVGoYY3zVKd
IYWjn9BJ+B1pD/2zm6jv1G1g9s7fBiK4p1mxvjxmkHE/VQB3ENSgo49xIuLD0bY/
OWYQbjVBItt7GIngc6CiKa0B5MPbWG0qtzTPxvQIbZOgEa0NPNyaqEfSS9/utQ8+
8m71/Wj+FZsYjqpFZJ8acaQf3DQWMoJBihGauSQXnJDQrm+eZsM5cPaUS0HQ0O8+
QlDlhjSEEhJ/O9jIdewjmflty2+NinW0MARziS7Ep7nMRflTF5VfZ1SDtWFP79s5
uwzmMRafWNo5xvLrcKL9NheC4Ap3b/zevOVkjecLGA0IjhImCQtf7kriO0bF6tmD
PYyeRKIoWW/M/xbZxRm2VSs3Qzkdx3JGa3xBP7iLnSCeyxvDO/nJBtZzSOl02Ze+
sHDL6nXMg80ufnQlrrul0nVwujjR9KFchvfHfVBct2MULmWyZjDi/eWzP1TkkatP
Y0QSgMlf7EHy5NSWq3G7+aTvii04CT6y5Yshf+WvPzokSBfyzDC8qV3Ottj1Q6fX
75yVnr+elW7eNug4vVeS2k1Yvvdo9wAP4edeLxY8ixJ+o5L4UxB8NtDYD70r4Xx1
8KHHn/NKCupbo62BTjW3VbmP4RUm30vFS8nnw3D/I5NiicfG1TVQuG25y1yzWsOB
u3LJp/dVvooc/UgkQtLaYW9coG/3d3aYdSl7bm9YwZVfyomwyp2KliumhkTsKlys
u0XrxbrDZT09E/nfuqI7le3ZZcjbEN/jEad647Ehqrg94E6EIaP98ukMZIRKSmfH
6XmRbGikbBjuKYYo6s2xQNSnKqVTGz9Ctb+lXiUe3M31tnRvJtHafKhvbBguYc/e
+L46DTnIy8JwpBBKTzdYnpL8aEJRPSD/+sdRrBmmdeT7H5mbVAqN6p5nDQeAPJmw
kxI0F2RT1zSMERoQ8PwNwIM1OLxybExXb22ejaR4h8vL8IScL37z1n93XCmp2qNI
pbvHm3NK2TB3Nl+wJqHsBQD1WaWcK/VNOvLJsQRdo/4xbPYM6XfbkB4RQklRwrSk
2vJc2yyxnbgg9gUF5qHqJdny9xFpI+U9Eqg/zX7xxcez0BhMCL20SD6x3arvSxSa
Q3leMd8i8G1YGK3jSfNYy3boAd9d5ZMQYJhqxcW82WLJBLhIHJbhuTs8iAZe85pk
WR4Ou8kIaJcJe4+b+bJis4gNItrZ6M+7/srAyiv0xvzQtkpLfDzoQrbcBcntHC5Q
XKZZ81utF7BGszOtWDExbpTct95Ih30PxYKvfWzoorfw0gyiKy4d+KjiHld00uBs
hdti1l+ClUicwYTOpG7RYxzJfAkgphj+qYoAxOinwOP7i5pJJraXrpsFDAVBvLch
uYu+pBBwSbsn/1oV5RZ95SE0gseYck+HntdaLgMl38jlTnoekpbuWVcKyE9DhrMm
kROItCaeyV01Eq9ONu9f5Sv/Y+IBAND8ssdkQn3d1SfAeFlbjXXI8b5D6jpyhL4P
Efz3fTni0TrNfDGQk5YFArrdnOW+g75uIJ+4RjWG8h5BrT/sFtCZXTRsHBFVBket
oJFyz3juf0YFJBch4y1ckR0JeIY+Lwgi4N88o1WXbPGQ67N7r70ujKpqfKtyqTkA
1PbzWzoAsMFinVnq49/xx3BQJ22a357YpZ/lQAJY4EYI5M1PhI+c2yMraS0ObypE
fmsorMrnN1WKKeSoFCQRUudWDd8dPlKy5JvUhiz8bQocMZXDkN8dyDBtMEaWUVYG
k76KUbE1gEVsB81/WSCe+UdwQNiaQWPr5dQ25APm9FBLZYx1akiAVx3eVNYfhiRY
SydanER4ADDCb9KOPfhAcsLlPRC94tTFQnTpTOslEzZwSPeg3gX6D0UF9Akbo4tF
1IRiwcU4VFsDCBIqpQAK/61jkE9eQIUP7e8jejBZyfTv6QxqMPO39tA+r6iiWdLX
A3nfWljkvid2j6RIY0jzFJSaR50iBKAjPrbMvDE7GvGGF3yX+zWX8rl/m3zl2I5c
9Jg6RV8zg6igTi4xmbwjMnKyNKufW70cEBmAlBYC+LGCmFDdtonsvQr4envd/CKj
iU/hv0NW+JhiuJ4WUeiqCrhTWFrK018QQOhPTdWhSFY0VUBL5A/ExbKh818FUtwi
ss9YUrrEQ6FT0mS/IV5dd5+L8UoeQhML9WdoXrQNP6Un3Oyw7B+Ki0cp8DpT4a6+
brYFN6OmXo4PXzgLB3bJ8k7Aq8S8HnN5oG9rbgEGpKV7OjRvhYXPPSCCsm8CuQi3
WapReeCvPz3408qDSnWVI+TQLQEMjmxkCuYaA0q7EdF/i5P9O63Su7JRSI/nDkzq
hOyHsaXOlUxDkQHHsDdwZjb+oU85ny0M6h7/gqCPR9Y8vVU59K+5pTbY1pAVGeX9
fhGzkvoJbFVgTl5nyBm5yvQ3wT0yPLffWICgPwDLjWIZlUyfu0KIs5jafKe2bnPz
ciT4bKunXSxL68sWUcR6vN8eEuntsxmb6WF0RP3WX6HF70+ORaacu09myf5xYfe7
tjladSUK1dqJT24QSvCBGyjM6/3E2DEQzo67RagXRKZJ5aTIoWZH7TJQN01YtrZt
pgDeVfeyvf3YJJRl9c8MyW4cy8BfvwOrih+PhIhLQd/TK0Qhc3sqKBGNBugQoAFZ
jBMzvc0TnOE0X9IFdAmExF2O5wzi+ZWeSOO23Ym5blxkhLmHigoNH0fiBTwR6t9H
W7255GhTxYIQoXKJfZtW8hmyNXE1TwI/fJPkLgZPkYeke4BumvQ2cCkF8dLx6cuf
OUsAivuUyv5LAsv38abEaZv8z/3r06P4ooxbwW4kQGG+b0uQ/yxB2TMno/plGNb/
UaM4L9I3JC8tYgEtPzoCilm3A/T/MWSbq+LhRcl398GGAR080QVslaLh+Z09bkmT
d0BKoYOm76gw2h45Vu1nh4hXav3Dpa661Qs0K0BVjuT4mFCho2oyLSbhpGZQlpkI
/x3fssw0Nfz8JvUHNc3APUdC0N4+skGO7Cw1L7LC5gf4/Q+hDHI/pJR5Hyr8IE+N
AqYBagJGLGsrSRvjEyCvjfpa7OOrq7oiSSPdEJwmEHECiMxcLrYjmYMrgupPnJi9
j3VkFoy6jptQyYh37kZ5YbS+rpmuZTem2j+cO6qwxmO9WesgSWC2um5H2n9fOFDQ
y0Kviz15jSl7l2WDZK+0/SLvK2bB/gUPcvpFggxtHzlVHB/TMjarGbQhQubMEvvl
vpgAL1klXPG2zPxVgYRver3/VZjkIswKgsv38E7SffaDmDT1Gkq6uiQQRc/rTVPG
GAkcJ9jL6CREa6xQn1xnkoH8l2MHsBgbIkUENpzQNpiTAPJjrbKjKch+u70kxA1t
J2tDeIBy7DoetCRQWFACpzAtcl/wqcB6wQG9nvpupglP5wRcK03s1OaKx32xTrm3
LK50F3M8LGT/KYoJXLEzPuBGAFacddWnB9b7i0kTwje3jTCg4HGAY2wYk1TEIz+N
wx7b4/mFZQOsOlIX5medVwgYpcXfzM8iOJ5M/KA867UmbqrMQd+HK/VypEd7GOB7
O/4JME7LYZLPZaLr77Mx/gfwez2NJXrCwuMCwxmUxiSIpNGmoGUjvcT8PRhflWIu
TOH/VNN9vdGwJwOhyfL4tI/UAclqnaHswg5C4IhG5MT0EyGTJr8GhGdndeEdWPjo
Y9dHtzmjrmRFkgt92hCFQPavCJd9lEci+v3YWKzfQ4IeKTwRncQFms8/IsRiHWe8
yrmJaJgyO07R2599mMWmoa5kawaFWmOeVqpmtLm7CiAQwGsteiadggGdmX+MZPKu
Y2fOVmYJi5rW6KHUpo/MeSTWFC+u/2uPqKxE5+IzSwoPmqg+BzNHj0n3XyQIwWpe
iV1c1Px0Np+DZOPTn2xVwuELAqhpXte1Eme8t4sDpgjbx/n2S6iKIVqgBVCpyLDm
UzZ7tOcSdwEDUSG+a1M+Q3vDvepRnH3J8lSP8aDRMv5Bs7YzAcSZAXd8zh7aGeLJ
Li4Nrn1dluTmAMCmcbbqbXrocx0ULI6Y+djCaqFNDVL6wfk8Or6VPp7q/Q/FmC8R
6eNs13zYNke7P16Qo/6KxlGSym2x4fPgjADdUnplv9nbhbxaEk6BPuBVBDwr709z
ccbw2DqBXSzjIdIzAT1Uc3bngKpbr8Jmvi63YiVM8dXumgExg2Op2cQafKDXJqYJ
CWjTqa5q+uMq1yee7oSZamKg71OaI7Hm5bqInO1FlCNNDQKb9XSFojnnMW3y9uQB
Wdq0yf9Gj1vPgX9MaOkeYHQgX0imq/Iev3O5HxHTPzmRkjGJuAFiCT8zN7M6Oh9B
f+C2MDu44Q3KKc9F9pVSnnJ4EVavj5tgqAbw3ehXNMOA+JHtMcR9HDNp/d6My5jG
QDLNNvjbHpglAAIbH1xTYvBhcstwh0k2Bu0qmeTBmLrR74K1LIcw27bHyMeaDNEY
yftS3R7BpdB/vAkclEzDIR1IftgnfquHqL5iDaboybhO/qln7XA7tChBJTdmL1WE
w+f0F0e4YaXRkn5edTziFfktLU3s9AY3JptWCrvrJ++LZTD1iN0Uw6sTUiV+MuDZ
vFhyAt476VRTR+2NedouLCF31CbcJ8V6lxRhfyQFuhGuXH9FxBjxLs0E81vxQcSy
6BHMIf4xtUERdO/mxTuquTFQouU+QI58aNm9bhtGY6AowNQ5ub0/l1wl6/A2AXxv
ORJKHhKWbcKaM230+w13F8I3U6rHzMCYXN7KDuKNV7wSg0n8YVha8pHMArCIjykr
DrOnu2G1/hphEYt+5Yb3xxqCnklrGZKPtr5Ru5oniWW6ty3lmFU0GoW/1KfOazF5
F+D/rD4xwGrVhB8hpVC3ALRpY7AVBsDhfnTwawauUlgu729702lZiVls8H8bG3lX
oWlinjVtTKW5878yMrCMe+SwPDm4hTuOu4uqXK9m+yYKzWDCnwMkN8bDOcbw2u6p
CFueCome69nrLZlPVd5jm1MziJcWDfMFbqdyL7+dO7dBShBkuD9DGQdC8/y0uwg4
AcoFyH4pl4hZkAJMgAEzgHAkCFMHPINzclk5AyFSm3senD7nSY+stNKUpnCfxwre
VSsD3W9lm/z+sza9wrQ6ySURa5l8NK2golGHnXZHOcTRg+lUTjRKPGjYKwJx4GmL
SrODH/qiWbpsxO7LqXgTiNGnbslUcWRnt4ezV3vYlSteMgvI5mDyyUwrPyGQTrVi
zdxOTIWV0JEHs9YNXfZBarVue6RAGlPrI7DRFxQW3U8dmCccnghMjl+1Ce/NFA2m
4MxxETWGNZtGKHsOg/FhWS/FZeEaxnQlk/HjldFUDAV8QRBKZLj+DMbvrMdih9Cg
nGV3jHEB+IA/rw+cqjtdtJOVzipvn4d8asGtwS9QvGaYbPWXXJuc9Lb1nd96k38u
WpVz6WAbImS83nEVQmVkEHZyV/ZQGSmZ4B02sjpwf9z+FIQJytG2lwDXlSGCto+o
vCA1QQckb9Mkc7vt2h749VshvRRUTml0oyn4PhAmTZpaCe9uQg5iSv537U5t/VWC
B6evCQnY7HJKlg+GBozpCOxqnRR2i869F8Kp+wyw6ytLMjW9J+4BCNaXlDu0uBYa
8GETGTyS1BgE4t7c6Y4KvqWXf568WM0/8xVlhy8OEhrcaFAB3eJs2PhaJedcYLDm
mQaJL73o4Z8Ki2vZO/3NaMz7JtJBNSLqMSFjSkLHEgNJ45HsZPxGC9vkb8Jm/xvs
sAo/3P43toA1UdLTb4joZDAFpLQsGiZiC8SqYceWBv7ItEtfXbNtTzWshkcIyJJP
pV7mhsdJcEwkwo0RKwnYiQ2ORs3WSKcBt5QIR56UR0BIZpIRnAQsHoEDMsl7wD+k
0RZ13kbRR4Q14Q/5L1FLuubAJ//2VUVur8IC6KX6TFrUxWvZ7Bq8WPY270DuEn5z
mj7rk/dI5ZhU3JffBaxV0C6lTJh/b4HT3Xn8eBfBGfoYerP+y37mSNRmivv1RJ2W
zQgfqliYuOv9T6PySFW9KSbD1VJAHcoJYs1ugG4ZpFdA1yQBneGPxW33McgWEYZn
kMFKGT5FGMtkuvjV+/OlOX8z7i7zApVC+0YZNV3Z8tFRBxyVZwsNJfRLMjTI5Cnx
amK0idnerP6tOuVPaf3sIGjb6PVc02S1o+DaE6lPZAlnSC5rhVcZoCQV40GHGWfk
tedut16Ul0SwksbPyXbVtdsM1riAaLAlfsWGZERbiHCs74XZCdxyLfhytJ2F+G4p
KZDjmn8jcmwASTWDMxC3AsrN55JzgEu+VKqEcPjKZw8PVjdnIGX3bJTucTTvRLXc
0SNBrS4zolNpHT1Yy6aN0x0lVL9/McDisCgKMjzf69OBtFvR9rNihBO9QZ24XtyV
zpBlQwy/TAxn6W5aCvmJY7ppnVH+vWJCkUcejTMnkUpknr4Q21SaQ4cnfK+8TObU
rme3rWSL3hwru2s0COwJBwiVW8FwS1/NFCb0NKwtnUjTbNJr9lGJTWbkrLADkn8k
OcdQujlUYpesZDuoQA4Mfue1a5/PTZ984xkWLSBDv7SrxveydAMHCDrbsp8CcpMP
vHYVq+Zj0WNzyY56txMKv7omBVSmAo4jPM9FJ2vPMqZZ6rpp1Ct2pB5JLkvTok2x
V0jQiajVgDmr5WZxY00FyJR+HjSWRLKVdtiHJdvQ5KN2JOeLZrzQurWcbeoDGUqR
gClwQp/6bkVq0n8qbBIs5UPhIvDk6dKXWVWGQyTuGezXwH3izZEzW0sPH8H+qXpc
jPRwWPXpytZZMTGcMtve9LtKSr8lJU0yiE1+o8pTsu+OPOQxRI6jNnLvqmrH9Mga
Hlqiy16Pf+kYbhUC75Wvlz0PJP4vyC13OWmp1roFAqgXZO3kVs7tRp6z0IAqFjIa
gfnosBcxpwORp5UkNhBSXZFf3wwwI+sy83VLl919tVdTCpLMMlZUSTieCCpxyb3b
Xd0VgkSVuZt1bJ/4gx3TL25w9KP6gPx4+eTGcT+FJ0ItMU039QXDOMyg1R8MkYSO
HyZ6TLJhSR6zWlJi29bowQTTKVd++U74NQIt8trjA6PAtfHHV65lQuWOM/qFjdJk
4NQVXvXgFwF0GdEGj7PA9zQnSCWVKUu2Lty7OzSJIqqYNVMskFarzvhkveW8x7Ai
jA71yAyPLs3k+ardqMJlukLdpbEfpPK398MxJ6BOid9wzsY3Sk4CiZZ9OCW7R0HH
ZRYN2ZS/HqyTGPc+mdpzxEn3RtuzSkItebKWKaMIuipwnoNBrmfce0OUCmSe401K
zungXLVN/0AZ5U7xD+SJfxnLaFXBLkIkfKm6Uec5a2Aj7D7m+tbpDgMtmBE4YkFX
fMCRH1/cTaJIiT4aB8bfsy7fQscOegBxVq19/kEjpzOmBACdrSFDz4JbXbZacfyd
J9AGs4rgRRJH7MMAQI1UVkxDXg3ecLPMS/rnY0bIPXO9gVKhGTN5C/x5XtmY8vqg
y42SFSkmuVGxNLmiLNXEdWSS7vRlfsIHNvwjd0VO3DMzBjPSKildSXNqbxrdpltB
9UO9GYdZ2S82kZZEsm0W8PQWJS8vwusq+fDLdJxXS6wmABd59DK7k+KMv/73BNr8
aQotd7/I5uLKMyfuadtbivEaePxIyFKZMh1fJlAA5/8NBrTypVjPXYqF6R1DwM5a
t7Wxw1lmcuYx2zVd4mga+mgGY8gVWFCcGhE39nGnZtT3RmCBF6NwFuwY09nPKcPk
HIHy8tQpgrIu/EDYHFB5t41UNyqZfv6Rw3hT2YhyQOV7Q3kexEg6gs0WOMRKxK3H
F7ZogjmllW7hhOW9ggLd8THKgWKJPzCABgQQj5fOc72OdbBsywiuA1tyu/J/NjDJ
Q+D00+xRbgeFoSBPysUWhCIQFb/BYl6lqPe4VIjZe9dWMSnueptKD53LxG0ZUY3l
z+lPTDE8azpeNEBy0t/yLAxVf8knwoKqiNTdGwdpF0clb+nxoqWzyd96ZShwY2SQ
xnhz/wb1cMtNwEtzqahkOOacxc0rKIWY77+tGeYyC5CsQdL/9iAtCCq35UpXP97Z
wC2eeOxOY61z4jam8vewFegus0oaWwuByB/791aUMFDbyagvntQ+lLNJlIHNEkcM
Ko2vc4Oobk/rk02bDdf7GKbfnekQjz9tVbLnEjamaAWtI2lBGXMehEI8CWVogUB4
vHh5Imk27BcVXYvZAanwSs5duQCUIblMyR/8TJwoSodHeAGPrJnEVvLLAEtivxTk
ts1sSWRUEp9syThHWiq7GOs6oI4eEYtPFp9UZ2e0qnxLaPtHCKR6HggEO13XQQSX
mPZMJRGPIpC0EwLkmIoMkEjV4xrvETPiqYwvxkQpqH+6s+94Nh6vDdZEFIcsceYP
+0EGgcE6J9Ffrg5ygqYT8Fp4XxcCl4qgmuSuQByjTP2R9fvhFv/S65D2LCiUMq8P
OY8mglGKVU9ZOTygur624qVuph1dT+4htmcEMiozOO1OCj2LX5oCD6I/c4V2hStT
lp/7YsEQCWFaJFJQJyYrRYO+CdkPwcwFlmWj/kpLzFN9Snw7Y35WfpL1A/gXmkDF
d3o/xSV27Hyhw1Sx+fWDrYWAH7KN9Cz7WbH9GE44Gwlhgng9zvT4lwsMOLGpEOqN
xWajRKvHBVagaa1z66Fm6KmtoE/qiWcmYJhcDk9PsG85yUFT4N6bCrwLpPgreIy+
FZU317wzdIv2Vx0viIwiLo0LKKhTzEkjTxhnV11zTC5S1Zi52sMqXIQDU+fuzVEG
Vlv8n51M/QG1n3gJPG1eOE/tiJY5BXZk2k9w0YcI2KMZW8lbGVBVN4ydyXkrH0Ed
tWzzfR8oJhHEJefhjvx4+L93q6KGR0AjAg6YJhQZ3uPS5FqtyPdPzZlFn0Wl6fHU
BSjsdOmI1r/CzEBSMOzUwIoiV8hBAg1SGJySN1B1hMJMHQbrT+oa5jF7bJifMzPy
584HlsgjyghdN1nG7lcp6aAD9HwWFXpHVEbz9TW9dCs+qduLRx3ZnJP/Pl6ttqsH
GFdC5IAoO0jDy6KqGvShcJlh53HeRtSaPbD3SB8oZ1d6jKqfRcOCc931BU+u+twE
2p4jfbUlYvNImkAdXomPONzppWaG5WroYUxpqu4Bt1XXKGEskSCV9Jpfn4wTC9qG
jGImnlsPzdXxuhGu5yXxjKwxKYXfO/NEhb5jtzQUy5i0aZ83q8Pp2RoPNaJurdIB
Jr/9zvSrhrclJQi0AlyOYH2K0Su8dwcOl8UQbgC8XA+7M02eYvMvV1qIPfGiT32Q
Yqq0XHCOd3+JyMZ49sxZOPc1sr+aeS1NPLk9sJmybElsnzmJ+BbgyMnCj97LoaEM
O7aftS8DeJPOSQ9yr33sPfMb3eYYFlfS28Iquy9xEH1J2gLod5R7aDjfskTBLJ4Z
gz+3dC6+BMFApzYmZAGb02AJa5glJ/LjTEWX0YUOj0pWy7mSFVXE/C/AOuOuA/Gl
9gul37UbyROsPyEcQiuPltY0+svSUPi9MgUm2VYODwGcq/tejKgVZGYpTX1WApdK
XdeqgD/xqZQUf+bn9sK+L6WBO4XukM73WWzAcWFJJND2HOwy97MJ/IjoMZkKOkWg
jrFpyzfJYayk4mPTCrPVVdb+v2LspVXYULUOc5PvPdPArax9ucE/PwjH1DEXczrM
RuRSYAhjRZMIvwQIDnayxf+9ns7iMSxJTlnBFef2bdmqpeRkzPsPv5MinGWah9gm
E5kIH1xmNwAvvEx543tFMDjIeeWDwKM9td16ncDDSu0QwDjDt0W+N85KBByACUmJ
etVvFCNOTF4xGorOQzfIQpIPnOCKicYDQbjC1fGL0rl2FcsVUfiPuWX+V5udrrWc
fbTI8TkE+vkiE85MI/kg+xyNS/j4TkESNKwWy7rvXY1CCnnQsiDFnE+Ott7eSXyH
tgsDZ31Vkqh8myYn5pxM4EpAXAyfQ7HbErek7zA5COf/FzA6JHSfjtN/sTFyQsss
bJFex9pOfelr/wYouCi19i2yUSyuGKhVr0eJ+YtrXdYGj206VuJ24FXxcpObVIhG
ymSw9OleaRqYM1WsQuJQwr5yols+OUquImNoqfl8kWeteMLyigFd6htwIczCbjec
uvCiTJU3VwOkasYsO53YrGil9LXzo4XEYxaEMqV0oTtB6IlNchk28f10kuNaGntg
07LIHs/7CB1+5SQbhxxr08izPmAHnJoyk9M2SaYu+cS3sBa6ttxXAgNtKMK0hV3c
dn8+E45yvQ7tufmtdcQvWVnrnoyMIrb9iDQqfCQ+YQ/Ohz6PclKsDFvPMjL/OmVL
bODmHpqYKIbHq0A4bqYkGkF4uJKb+3BLj9E0atpFLcyCgmbY/FH3p2rwPvIWqmiS
hPTaAeQY8eDMJFGfYVh83tpw/YDiG7oDdMxEBd0/D2aNBtQCyzMeOo42kAM4y2M0
e8VPvbI6nlqrIuVWHTdChXq9g16uf+bfu/rNUq9qpVh62ptyt5nu3eReOm03XSU0
JC1Z3Wu0sb7gUuwRdbPQXmhkFzIK9EqzjcnYkWvdMvvRcVMLkE+Idy1+4FtvkH1g
NPL+2Ec3P7lalOn9PI79GEkFauzgOf05569EMtTJDOsq2jFPVQw33kLwbd8XosJq
jwlrKjMeTniXcy4DR0s/ebVk+Q5Fu5NNi6yjHmAavcAQhVTTs6O+a4AcEXPzp+KX
tvB3XT5B4uyu2UuP+BrHIuGLvMolk6fvuVFQliH5zGGLBECj1CRW8IpW/Sqha+sb
YNjIBC/Xg40Jrc2/Lgh8Z8GVoZxb4fLNow+/oRtBDgUWR2fD2cWrVw0SrUd3E2Lh
9RJYRnRRQJxYV2r3vvIj6hRt3epNgcl5sGgZvaUcbcvWXsd3SfqODy74R6DaDN0V
S+U+mPZNFYlS3CgltoUiW+FLYqvDlkIGsob5dT3M6x26nwxEHHceJ1b8p/LcyU1z
a+4Xld9ojZQB7cLp1Vy+sztuVii5Wwo6zd8JGvicIJZMKpozMwLsxMO5uT/mnKDd
0rplq7HFPog+lf1uyxKu7td9kHXrl2fEX//o2PjtOxIuTbwLNh0QqasoNuMe6Wgp
qmDLmfdRAl7JRxsmlsYdHZUkVuU5FqZtN33u55Pp86M1fgHA/HE6HzJ945qz4iWR
KHzUHY0qzLQMQMIM4VCxHbI/FIDGzVidg/5do1bVxyNOfJO0AD1ogGSHBb6Rxu+1
OApaDmsmewPgQ6m/yhr48XyXwMhcYtKLJ5FIsmArrF9ZKe36+qKEWQK3/jj7EXu6
xrohYypgBfgS475EL5tKrr6YAVqDsTpRkMWF8djRnem0toX1QjQqpH5CgNVUKUN+
+gkFMgJ4jvNMtoTvhHuuA+pJ9rvBLHyiKoQdmuni8w48TrWp71b0iHSZKq3L2LX0
qdRJ/0Z8z4zqiNWN9jVrnR/anvXHWP7rRA1BsN2o0J5Ep+yGF9rIMe/Xy6yniwP6
sW2g6/SKIBxk+hzHqlZqqs8TxF8y0Ya0w/VV6KwaawhXxTQPTck3JDqM6a744Jtv
Q1oCKbZW9D10RQPXsLCVD6qk15TMYU6IOsZrQ2YTbr2Zgh8rFCSH+LQhMeB3HBgm
BtF842LoUgyJEzPIhUKz7sYylaCyrqc6z5lYisInSKm0ebanm71UYsu3kUYMYpWr
c2XU2hSJo5/+626vuKLMoLrqyWoP/rvYwwdtYeuvUT1CxEwTlXNz5MeZGag+vA3H
B+6baMi9NPaaWNfEdtVQSsAQ1PHRWsVQMuOvLst+3JJTXJ0BcOwpE5pl/Z4x0uDl
pjRYiRqLNnQWc+5CZiqt/OwcEDK4HsQc7Xav9qD+tqFiWFpJQ3OWqY8mN34PFwk7
0nDMF4saZrEfNpWleJcOt7aRXfV3JL+I2zhmtyTw+cUPKgVrg1DiS0Y6xRx28W5F
yjZrjX/yjovA4d/w1KKV31XWWPHUAmrdWmHANs93ON7K9MTec2Ja7NPn9w1/GjzV
X3woQ3xIFZmhFLfFbbhOeMzalJg7y0LMmQn77AtlKihMxMHrpIkVtt/O7tHFwFRx
EGe0NVhrnx+gUmBZIOiNGFZHza5q9ko/iIZhuFIxb7Aq4GmPelmrRJ8QPh17WW03
9nyGSqJvLecEOdh/RsehuZk6EpWeUkHjSeYrqz/uNz6g3MtEO3HNPljqJMUk1kfU
zQzRdOyOMWg4xT6TsScRaVncpeDIZEZOLyoWdOs8iEIrmHtXdDBwLg9ux0ybGnEQ
Xoa+8cjMcEbPfdr1xZXFQvRgu7JPXkUuuqRgLdEY5GUIP6ZRjHJFVGUdO28ccYFT
2kxPaJlux0gDGrSwF+QGQMhQZDz1exKgxxii3cdqdMxct8eKzMRHv14upxk4fHg4
HoS1SVD1ZTUTAGrP5DZryl5jS+ggEGA1q3cRMVSgg3zLBnMN8GRofO+cC9WdNFlz
XR91A8c+I5M1LpJ4Iv1pG9VWDXTIa2okn9GL4CyWVNFLw5zoQ6g8AsagpJBb9cdj
aEoFbfdbTvltaANA09Aozd6EdIVQ4bnLVo0Ns7sGATMouPnasZCzVxGpOxaFL3Bs
hhfc+luMGy/qkQGjtddbUI3WcqJPZeAGWzN0efXczbkShpH5WNU9W3FdfQxVUE0a
eNI7JkBDK+cgU87suPe2imk2r3OgRVwjQInmAf9uERbeDdaP2hQzTwdTTLUQ6dyz
Rf5T8I1+OMHigiNoRmAlh9VSVFr2mTVcMJ6/7bY2veYJzuHyrWe56IBQ65GIBRaU
SqX9hM7Fu5gWKC7t7BkWN6f+NnOsSxIIZcD+lV5KTMCvGb9E3ZkI95O1GE5IA+8U
yPdwKdYs1In1Fj5ucQ+ya5rSLOeNBk7vjmZn03AskpwbcFyE6E+dzanM7mvPz1Kp
VSIVtkxknLEmzS1Z0kQt51sryD+r455/1KiHD2qEEWTQj4cViVElKso2OlYthGSe
aF3xQVdd4EcO6MKJMb83lo6ReFpA5QfnHsAlmM8YEgSPTtxderKtsrtDlFtaX54R
0o+GhzkcPru3jzkbUir6PsyzS64Z4xyyEMmtJNiC7Fcl2J6+pW8kXUSGh1ygy0KM
ALZTQ8TIU0BfMs/Wd9e79CiJQqtEnGW178Q52+I4+HeiaoJO1AbA7eRew2lc4Eao
WGR3yhPzee3tzkVKKNisdH5pOUbbe9p6nYUofKZa6WZCGx+dBBQT8HdSKvJHmzAt
Xc/6Abq9QoyRfXhGyEVzL2QcC6hJCQuwdkKF/3u7yk0mcG9JmD9wQLGgFWjFxpNo
yGWc+TZEclH1M0eoMmqk+d1vuojzTdIu30Bk0pY3XwSZPb4/+dpaa2NcGTTVbn3n
jHck67FcqPiOx/5Jj0FnxtKDupr7cwTpik2W75He/2dhbxVxEPXS5latPiaf5VzP
i1MjpiTVoKrgYaNI4qSas+vzHsFGYCteBCFf7ZdKeyAIu9Wtkk1lHNRFIsRlg5Me
qgn3iWei2SR3o3G2IiBLTPlSx2C71LwWAmzL2/x8zvxd3zIQSLk9D9UiQnIRxDRJ
eC0UCHqMHWuPaXnUjERVgKlttyNzuO2PRuj0NMV+Z6uZTwcaYeitx4FEANoo6Py5
0aBLozjWt9j2mAT+4IMMvf5xQrRGADKhTLTTSMWH90I5VIrFXFQky/N6we3MyZtN
4rqzrvviz1bhhB8oW5ovvFnJqNE3JFp6LtzG+4VhDhjGCZGp5EKxZYODQPihmANs
69EOlkQtvWCX9yEGJ341SlEHB23RztNRUJG4ZABlxvOrSfaIYaEBgKhsuJwZGE1X
2ewt0hYrm+W1sVhtum2vi7g5NnMljvxoNkEaYw8W1isiHLC1M5EIt20UFCQi3XdD
GIFYOhklTN8sGp2COZhhaWMRAo/aj9ga0zj5AzzO/X3e/ba2Qeivis9xXUtlqxAg
gnV2XTAyqYRjkg8+xuYBGV3yf6XV5P4l+midQsr3zJc7yCFsfNCqx2uhTCGEAeLh
F9C6l8hPWNOZTqsSrNaGkmmDNKPclq4x+mA4D6fYIuT6gVJSl+axBVAsj3XFP/Vj
zoCJVWE7RatwDPuzKL4OPxkmicIYSVGYU3uEezqgV0ZVtZu8Bn4H+XOsu1wDNuLt
Z4amAWhH/PaGYajl+GtBd4ky6PLExhJxzHigy7gMMyHvNd0JCUb2HEBTEVL7MkXC
TWl078Ehp5XpgCjYaw1q+60F80j+PoBI936qoS+rtWYqgbySVo0ShrjmB72Cprdg
IWCk45Gp6x3UjZbxj5alelIHfATsSPDtGCag2WiMhdpkW9P5sxQ9Xz6cINSXMMTO
GonWeG6gHlPeg86hX0r43E8VvSqv2RYd1/un7m748A96g2IC0eDIdepl6c3G6taX
2yKwkCgze3X2qPVWqeKtZew/BXwhCBdDO7vDxe5UWZPi8bpz7oBEChzMjUJoGDhQ
brtK9qpOj8fJXObhXvCOKTxED6vLCfBQ3UMq6PCitIodm9ZhwNY5ow9SljqSaHQG
FdMInjV93zJ3y7kMVKi1hAHijz838nDq6pn4TDZcpwytkPCsW2wbQPJu5bI2m6ol
CfuvM4kdR9Ltn0QrcS8OAqfcj3oLaqLO00lhb9p0dnnPHPQpAYUNLndm6A9TBXDa
amJVi4WJ/fSs961TR7MPPyjxm7xW+ZNjO70UjPbOL1YXj7iUuQoPz5MAOs4mQOOs
WSTu3ewXgmS3o2akUvQRnAhJFxvlVZuNgxi9tCP8wuIr2ArmGqh62Vwlajhtnnkg
up4Chd/lrqdPueMR8Aq3SKqMr4AbtzYI5AFblByC0IBEszbRwdkvdMO07AnsNb6d
c2F9/Cyz4PU1X/HtI7eHmzDuFfL19KUrCr/0oLW7ISfib6BFuR4FlpZqAyjKsIFc
pljFHD2Eo2bZ2+KjOAuE3PQeyy6oGpivLeNa6utq0qc7XTOzbZwBoFJ+E3wJ8QB+
Od2ZcL+1UUUEjcAwDNSsETYTCpKFZDYTI6zltigOKkttJHG7OJXlOnAe3tpiO1qU
0XJRBuLjuU4IzFRjKdLOZ/5/j2LxKt7nMk9AzjNiN66zmWAsLpedusKFq3YRfsaN
LeY7gzniSSeBtsyEHMeziU23NwG2/WlWIIfb14LiO8XIrMY90ZcvxE10bZOopowZ
MX1m2j7qQHo+huvhLDyyhNWcxvAA2qZXflbDvdUcbmnFSUeBz1ST+PBt72RWWKz/
PaqzjGtaNG0kEC90zrmRaRKg9mT2dDW2T6voPfQ2csE12LNlqB57TSNgBNeFg7t/
xAF+xHqJ6kNdx7Zcp/zlsqxUEYEJoeEStMklLN0reT12qyhSG1epL8GJ36DFI6UN
NcU8JGqJIX6+VLNDQZaOMTX/Jjdi9SsH8NyxhuKmy7891jZ0LGhLJKWdl7Dc4i9X
f3zcGub9RWpT0ndLwn5UxBvdHtd66WVmE2MrLFSJjXqob6Dw2EWr6sGsOvmEAWAe
BhKNnIjtg+H9nvzYRrPpc09f4y9LDFJXMfupk13Z1gn6EXWvK0eHB4X4cfpBONRy
pZBmQoDN+xpGpSN9+lBbDmiRrYYFDjE0LFn68lDBLjRelpz+QHh0ZkhnM6JYfrwW
JNeeEaQV4uJczs1bsswQD+nonknVH51AZIuIsmf2PDsDBK6skukwsqKMzfaEohJq
x15ASDxpY4/dSMCOwP3lxELT179wmqFGd7Oc6TsgYZO5yQ5LHY82hYgfj3ymgUYO
vEr2xf7GNzp/qHzVlkApSEULuJuvOhd9HLGIobezvTuNxRaBvTOIH+Lz4rbTUCIk
jPU2Y25g4LXYciinaVN3ZlVIfiUjWxQDiyOt6vLA7SR3xWHWi+fgpcc3mXCpG3Ff
FCQq8t8eA3ATeXsrjED6bPsjUItLIQtr+4VV7eAUuWIb+wA0XM1M4i5aZ7Hx1t4z
kCE0vjA+VGD0CkxV9arUduyXgGJoOeDDlMOBx5z2n0YVxnXQPsifmx5+yFw01z1L
2/cOzDDQGX3dvqKTOQGZnTB1mckpPvTTcEt+e6sRFgoujlmAGg6RrX9DaZf7ZUM5
LT9o9+DCc3606c+Utl9grKvyM/eKtGxw66/oaQJd56iowYNEU828uFxmlAEOKbss
1VeZcedY9/KhPv6Voe/5JkHaiRtrVOt27BZHzGZEzp4dHCZ6d7nVeFmJEBt8a3Gg
nG84qV/GipFH2ZN1rUThOAi7y2ttDL/Ww+Hf0t0AwCS8+ik0RCSCGQZ9O+3Kgfnp
LYzm9GzmecUIu5dNrwrts2WAVbyKDBZr6RlpHf5zsLnH3Xz/AZMngfQ3piIHVWTS
Vl+1J8iWU+1wRah74xyn8kgRWkNFnAU4z/gS+WKOwTDHDOhR4oRlOBDddRnHM47L
T71HMi5AIiAg9og0qfqSXLds203RIqA6ZkRgAnw3Arbwxk9YCGwxlWD1kkI5YkpU
/Mm0Ys02kT/3ZvYXv/6eOMkxoCE5ZAt7Zjul0yLTUCGvr8IvN9JTsarOsFO3TUqO
9R1qtSKtHNKjb3XKCy3F+Y5PCb1RvRRE/wQCGx+bCwLZgPqbRdbdYQHGrdaRHKCE
3L87c12mLZQRyKb39vx9yWQAjdSiekuDkgfjJ1yHeG5Lc+iaCEYAL1yOCeiEedbZ
VJ7SJNJh8kdwx90zl/b7dxrTxGyBPJlUoDCuJIGME0aO/GYi9CYtal18igye2pGJ
2YDfnFc7oWQKI4yNrouSNBQR3d6gVzz43HH8qtazFbIFSEnrYoNvCw+brBxb2zAq
6WrsoBJZWz3u4YuNuic8/LgG5q70sXZlAg0ABLT51lt7CfPuUMxuujIxA3g0MRt9
twfOcu+Q35TxjkbYby+sJqkYs8j6iRL4RZGEwW/E4kWsFFjihqnRF9FixrWO7gBa
Ov5hZmpMaxCWLm6uj0CTpmnjlHjZj+0IYDJjCpw9vBF3RUCHVsORNBUOlJ17a5LS
Ir+nyAOq5im2fAZSXuSkgZLN6n7/eQE0DzP1Dk0ZLZOlq2tKgf/nkp9zG8GHY0x/
wEF9YdSXhSrR0g4sp5dnq3M2wzf3POfQWylstyEmL++yObNqS5HWd5jns/rBArpb
KL1Rmch/pNco1rxW29xJoR4mf5GCX3RM2ODMmpXrdLevW47vGwLL3tNQ2WilW/o2
ZetFgr8mxjEbSafb9HQcRaoqU08QC76eURC+v4qyfo1ebaptcWjNfU/xUX2hXKRs
y4rcwRwJH2YeE39xZukUfnLH4i/AUnoXHkdjwAohhOtYz70+m2OFra/N5iLUvhBE
f/RcRarEo806ZzZdjO4kjsDRN0jmCD4k6I+0woxYl9UfEm8lv/cbbZM3qf/AXK0i
skWNo+9+SdP2VnQDmdoOePLsAxtFsfenuzj5EhIpD4w3Cl2jhplsKtvueoai2Iw7
JNnGrmKa9Wr9v2OZCuqugVwtZcHKjkbMC70kBvYc8kz8EXZVwsjxVLr1vMI23eov
9Bu7QaTvLeyxVbIhRBtMX9kC3/Xgrx6dyEFpeMKAKepfSlKc2MfAy0E+dbA6asRH
Jqa5LXsfTiFNW+I5vq04vnGA9qTJH0FQfuQyGF+0IiJfl7nGQn7GbwFJrPlBRVYz
EuLEZmV2EiVMEkTcixIuOFfltU67T99F/luc9BhAUwp0kliFuQl2WaOlCzostlGn
YEB4Hw4A5099/QjqS1HXK/1b6a3jRefsDJMd7V8qjnQVSG3UjiBrDj4aElG4apZF
4cS282uEAMva99MXT0oXDiSkKqIQNxoNyXVwphZShG6R5LF/VOIGRpsO4mr8rEyw
aDNi+CloeD1JLWiahQ/ies5L90yPqiF1B9/LNlwhaKZ2kRO3EfXPBQhO2N6GDLBu
LGesDD54g+kBzWfn4Xg28xjeLoufbnN2RgPXcOmntv+wn8kX2XsCy0wAojsUhnL2
wRQTR+RievmntFm0qpxObXkjYvufwO/N004S2mf0NT7yzd63uVXOnKOnL5ruCW60
A1jLziR4w2Q9zPJUANlP7DMBOYgShsOpWaIpAQX5JiF4iEoiPGe+3YzbfWvTo4dF
ENbFAHlJuVpHupU6jPWOarmtqmj63XO15ezGWaqPNCOqnaSiFTbSXnycDKuUR4zs
3cASP3/wxwYkO179rtLIVYWzRkCRwqxaIZNAKNjrfsvZQrPOo0FiThMlmlrnPWxa
2v+b/YqMLNk9GU1impC5p9Fhe26ETa8QkmVnfCVE9prrDYPBGaRNijKWBH2hiEC0
DtqoAxQh6YyC/I2F/lNr9MZfZdP08utxdTP3JN7iVT0w3JZan0ZEhrQ5CvG37+bW
1fe7LJVs7fYSiuP4qskBOluRe+vxNSCUZmRkq5njwzdCFofUy158Ed7FNCZtLktv
MufCDFJVeymFNfrCMO5zxU58w0T5L6RkB6EG9N5ebBz/wmfaUV2+LwkCGa+St0Tx
Yfv89dozb3ApaLPmdvf0lZgYfbwBwGXVfH+W41/ZJzByF5v8l0kezpnsCD0aL/HD
a6dHRJ5IcZSOhQcYTBMlcRgQ+HsdIWoOcO1OsgG9gZp6ElWvG2fB620YPe9nIWs0
PFv7pd9oLzuP1Mpww5GQLehpX/3MPGJeDgvxio6xXCZ29goR+y376iyLiHXQAg7B
ceuw4yvT1FnqXcKFrVl721S1fSFHxH+8QdCWWojaeDf+gUwGtUuZp0qnpcfmYruC
8aQlnLvQ7KG7/m+DCtytmsSfaRaMVZzsuT8CcI/m8wE+gqnFf5MPtDGyEE1WllAA
SHzG8IruS/pFk7ec6UjGe0ldlwcwwR3kbWKphBdtNMN9UufNkwNV+ueg/dbdG3MJ
kBYssV8IySKRe7Rm5oyw79ulBpz62mO316vUJOWzI2RC01QVJTi1LFI4BTAhnCBU
ITbsD6Fk+pOkv/CqF2qbICLHy9xPdY6goYtxHSRFWlip6MBu6deCtKd53H5XtYEf
mxksrkzRkmXmniX6zHSwFKo88tnFwnG5w/XaB51QJ1ZSS+leevPqZp6Okfsmkc8b
sTIndbyL4i/O6G8vWOWrZrfke/SposcBGrfpcsYCtZsyhJ8N3lhkBAi30aPImqMq
UVKjYYaht+7+wFUuLGFmrzD508ysOzw+XW5+5PKrR3mxYJpwiFEWK3C5iEDSol19
7R3DzUY7EpU5tbos6gW5Br0ubuOs21B74ssALkDdmCvPxJivuj+WYjHUWHxcqDN5
w3KoLRaGshVINwAUsYrDS2CLqXYIjZrw6Obu2aftAwGelFhgBrqQuu+kG6T5swQA
NpsL1vd3Wn0+oasNbpbOFhlOUHbrezW9veduiaDmsp5hEjV/ay0bViq0c+6pkYsT
yZmwlXl7JtXwcODo9uWKBhAHZHrKzjIjm9YZqdQ36x9E/rvferoatGy5iCNQrs3x
odFEruPJIhJ8fw1oXhxrrXJGrsnW5Z/wrZLeh5b2MHqIGnXgI90HIQtADnXZDZOC
1H4Uoxc23wU+9byMyi4ESGhbsoK3MAl0j2JlGxg9dA+ChwIGsoLhqShkC2lso3si
xVywKHNibZ/Paj5vjsVLe3ZaZKWSXcYZ4VDD7s1AHGHRKbxiHYq2n6yfKzhN2DBP
tCbi6tBDLul/iJp1gOPp9Y0tUTLDrx8UjZAt2QQ0OIDWGgKEmplv9XFpyXVAsqV0
DWtsmq7JN3ia0W+OdkR4O46+EqyUy+aL30LnHXDcb2gij0+4GX69GCLVTLN0gYQ1
r1w480xEq3DsxQt6AHYRW3ynJdSRS6A+A59myhFtnXs62uUwcRV4flxl2mlMiEHf
1U3vTVHqAWT5liISOjVyWpQIkoZ2GP+aa/hOYbNuBiLhWmvG98jeUJKNv7EFDDkQ
GqcL0JosXLrGPzkyqeEMidax2BeOL1cVo7bftErJJS7UVVn1bcu3n6fQgs2Druur
agPf8F1dLvoVhYDovj97gBEYwmTV5JctJk2MX7VqirLmjB4SpTfqxkZjucsCby23
og3fwbzcJ88zeWVzzgRdLUE+tbKOpLjYbPCo9EurjkRq+5+adjkxLGM0KD/TvSjd
cFEUsBFy2ZZEeyav9bwjWBanvhcXMJiRg3YGRM625a2p4w8VEOBDvoywfIlPAsQt
XHx4L5aGsC6xxIxeDQpH9FjZaoohIhqbCkZGcK3prALfi87/egjrJA0OYsFNxlA1
b/nADSfLhrpQXkhUkh09K+tF17L3TMQqFlmiv6R4Q1pBh2tkN97A8/tErYzqigCF
Z2aYIb4rrmkFztlNmIyUmp4rL8YwLV+G3caunekm4Cp7s5/wUPOgcEMKoMlMmuC7
53whvw3AnvysZ33zfMAUGCBkP0G86heryxb4r5/Rx/bVgkSPzls794+k8dLj2Ijl
MM2jiaymW/OGEXVdaJnvSkeeSgVNxL2+EOTgWhGl/x8u6AbnKk4oE0ug2tysHlAG
c3Cluf34UaX0vyrd5JaN21Re9Nme8ShnlTJF/DH+9H3UGGjaQNQD6Svv0T5C2Xtp
FOoy5qzHif4ymvwWzclY901DYpGC0pk7ZMegCixvjVBxrH45DoiySTxuNLa2Q2zx
chrHT7J2cN3e7XGUlNYuVuiY/TDvUM2YqY7+nf/0hK0VHWd4R+7oXDgZECGZ8EMR
oretHM8O3UafeBq5pQJWwHjqYIvDg5iXCCT0hAj8HusbZlTLSzxsWdFUCjgcwuOk
RDrEOTj+1qzjW7NVv2DPz/2rWI4UOX8ZzvutQnT2ibw7Ce4+EN+kGzArXo1/t23/
1NfdrBdqU3uxSBp+JDiIOSqZVjB9NhxI6HL7Q0t7sPLlBVIOtVX650KJTt4VjX3w
itqDuEnIaJVhHIHv2qKwTELvZcDVovcjAEv/CDMdILNfIxUbeuk3rnms+GD7YxZT
l5Nf93NWlii4cUBgKFy39jUHj2JgcKaQDl5cMhKyv+5bE3cYqzkxyN0Uv6SM8EA9
H/MlMsfhJGKqqMyPnD9C350ZnVuoghHO1QuNiWp6W0mtRJn9HHmgp1qhvo7y+Uud
6nJLjekryNW7od1cxfHZiVvBH71M0ENmatEMFK2SHchKy4I25XnTuTS6JutzBQz5
0zIYjLbmLk/SFLBeellYBkUc3CgYyvIdiPGNKFAgJoB6/0EuoDMBCWNDhzYbhWvV
VDlqqZ9hsfkOBhjDkbMMK6hx5I++E3zjNrgT96b7gcLOFE7E5jv+/k7L2ACUEAkl
H0D5ZI9O30jvfAd6LLrKghgPbl9qggP7McB6V/aEPmC8J97kH0nJbuf8Sw1r0ChU
CqPZGDKseXFYRsuB6MdvnpDbevkImgmkBoaET5YuKlmkWlyuHucpEq//DdaYc5gn
EeTWocK3bUCGtavSt37oLx3OFArXhFY9Z2cWVL+knR+x31fWqbQ6AoHkZ2vPVYkU
0lFqZMW8P1/wHCe5TF76IMro38ta8YG4q+XPmii5jeGcuT1FEXcETA6zviNEYsGx
cUZ6tOiFM5Z1zlvhA4MpJDUOGt7su3wj3iTRL5FIkNEH4yfBXawKIhHEHnGYduA9
f28vfKiPOkvVA6kxXwp3sAuvZWBTsjmEg9NSnULhpIuysQ/cAL7MYVwIZNb3mngA
1J4vIlnNcOhfRaMKaFSZguViq8CdXsmBTv5yewKUtZZ2MLZAI9cATIf2PL0ZNuX8
mP1NwM6o876hAhrnhCql/Wo+aTQktkvXQEAVlbRvLnEl8wrY7rQZ7ZKl7+eIltBd
xok7KmzJ5RojzaqLtqBYC8mYXGZb5NfL+sRHRWyTGtocLBZFBZigUlStEoo6rUj1
qITFsBZR/3cBi1Ih6mFi97e3G6VVRDy5V6CZBZ3Dm3LI6IR0su/YW00rRReby/rr
Kor3gEKQcdpnymY2eawuck5CL1esfpgz9snp3x695kTqVl5lLajdeJS7CTBEp6Sz
v6fjhGakOqB3j0DFAVCePyQdQKS/ofpNYP9Y/EsYnVBs+W8otZAO1uV/lKNn1+B+
1mZg+z1704s6FltbGy/FXtWzyYtqvZmy4koW01FM5jCcrsuPKALT+AyVTsvV03bm
zXCrTeDQDXXLw+ZD2Az5SnsoqEzska5E6t3GRYnq/3e6gfSVQdHiHsEqN8nJenmq
LsylHbFzPcL6iHsfFkUIfWcpMdQVDZ2JAvBFpTSAF6lIegF89MPJaEpTeP1zVc54
W84PLSRZ2BHafXYAV0dn07wplJzrb3UVVo4TkMoE9xBaAhdN9pVVTICg1ia4zpOP
7drAgBnuSyswIvd2fc2qfbfYHvQRhKOPgPB1WeYV2BEiFgVziLWS4XNYXBe84kzS
ZABvup7JQvFX7vYRv9tXCOd/hLENSXTtbJ2rCMqgu50F5Z2RU8mpnIrkZQXg0J+o
OBuYKtGgyoe4MiDVtgQF83RlqQIHzCWuMHWOIFHJqut1Wrsa4ev87l0Es9kioZP/
FMrEefgOe/CRLj/HYo/4zxURIP+dkuDkeAWRXF3a8aW+TQ69z71zyqmugIg9faMl
OijheOzWqRwasRzX3t96joocTmoIxTpKzS2BQAoOV4vqEot6PrhMd7pxQ45GAMwb
ZvIdKFK+ED7Sef8j2eMsFbqFnE/4ZZpBYTprpUIlr847WJ85BGEVnHR6JJMM1Gh4
y0u46ra3crVns8wV0q0Vv0mkS0K7GiDrp37WrohvpWskQozLezvmbWCul9+7sXgn
1Lv8XwMJMvuqVaAuipLXfoC55KSanZ1shxZpzNXrrJ6tOss3VzKbeBxg0gZeEP/S
BwWnEB3io081zY//aGjgk3v/k6U4nIO2o9rvQZMz1MoazflOqEgO7yNJvixwqGVt
HgCvB/ZM6KduWIJLuF37y7BfNDXXaghfvRCxyD/Uye2+vXaB445zExq1rFne3fGJ
/L9tsvfzTxs7NLCxUYkPyxFIqoNyVqFdW+ZQ6DYgGb1oTWCBmj1rKfzYi1F+vBsR
ePwbN94cHU98QbkB4M+mND/pYV78C8qPDQCIFxrP6s+fY/OZZpZgG32ie40akHGc
52wOjWeWt9eDvtVcaRwqNs85uNGW0JmiQI0PntGKUhgDmnnlxicbYrhFB6OQMovz
/NSFGnC0JQLTUz4ol+C3huj7IU2Aan4jli9lv9M7XWkMXCPDh9WvLtgZymwm12by
BL+DZ0PvxNLC9CWcg2w4VVv/7N9iygRccpdJBkMkiWwOt9SSM3JjAWHvPP6tqVx0
QN6//85av/YrBSKvzT31LJTMSzA9SlN4rg4ohjPUltfI0JDCHn+74nruEL852jyG
rOhndnfxynL7+E3ZCqWLYOFm2gISbq1UAZSqhiiaA42KyOSF2U8HV1fN+SfENDt3
M4rSPJnXz0x5n71X/lFoym3aZ0ZVN4L1+iDstqFACVtIqn/UGHqbqOl+pRDJtl/v
O0kBy5JdBQBWpjwknBfPMqwIswWfIkF+MePEhpj3AYcbIoOFVf53rSKfeER1Eiw7
o95qfNu60QMeIcbTbuu/iHBpx+1LoT5Pye64BI/anA0uMm+scYOEqjhKg6hEQSt0
QsRSHACNtqhG5vK3gYWqzaLUodMQSfDF5Mo8BqHMXDlev4494QvEWh9TKzQWmrKj
YaIzMve3ekg7CiXdStUDhlA8YyGS+2ZmX1cG65DxYfo3IaCw6eCRaxQg5fsy57T+
bMCPFTZireAkqo6tsM2YB1PfIo7osAmXrXDJkvKWzXKBsjR4Yqe0uaCGCyGwBu4n
yaqJh9+VJTOPncGQ4QhzKBrfeQ4Q+AOysHOYP9VqK/KeIgvl2V8celOKR1Me9wZi
ThEvA5D+oYyoXcIHi9P/PVu4hHT+hbLqofFk9lODDD0WHfr7/Y/ZkpithAWM8AzL
4CUBWJJGlTJpxQjjiFDnBGuj8Jn2kOOcTL+ZDzOYj6d/Df8d860RsAy6u3mwRpba
QdHGwSkSQe2/xLO/NKy1dfrYaTOoXTGMP+O71MJU3jOivOOCcxJSa/5/BgRJACpX
EMJ0pMO0pk7mY/gPUGb6WiZ5Qof4QEma0q6A1aFcg5PO0y6RFpbWpI8/jyso/H3R
IImcj1AzcqJwYJIygNwtXdM0JXbOtCZzWwANNYi6shIUxzVPbMltQOCzjXFIPJ/g
iDnRDqGfA5p5dk9Fo348E1XL+TLlWvHftuep1v+LW+byzD7dcMPFUQRxh/lI/Z7p
gHd1vvrGVxl31x9vkjpxvsi0qfd8TR5z/k2pxj9BxKXJoG+O6kZzZ9MFR29E7N8W
+htNZixvDB80o9inyp6jeQJo5abZOJv6uWL2wXCV6HXtDnfcMU9xMxD+3nAgmsqZ
TCLje0ZPMEwzIGaa+SyLnQvH/eaJPaVQH39q8OQe1ZB0GYlRXZGtAfpFZg3R8XfF
diqx4sCuWeX9P0Q+WXSrOo8D6m+9rDC4vb547ofQ7aeElNCJ34fIhufd92jTzc+x
d9FrXQIXrPmdvVD5DD/K8MDCk5yT4v3rIfBLY9oQEjO74GE+EpGUli6DXbGWO5gP
s4voXBzEj2IMxTpyt1wfkThvGJQJT/2XRGmzV9r3713KCmw5ijNJEr18nkf7nnLm
ManNPNyDDdiiU55wrotb8PCXzzVQK6Xbbv4sSAKlCmUi/u9tSbFmJCuametJI8fW
XF1fm5jiYfJZ6VX1zPW3nA9yn7rA/VzCVZKNvIW70W+aF3ib3G+MtkcTlQDWS68i
uGEJtUvAUTFwdX+bEEm4v/UbVPePMgSGwPuCiaCzBu+K3W3qLZFFanW8lrH7pXxA
AzuBPwAfnIjspHQGQEPiw0Jzr6+SkGuqq5n1CXIo4L94o0PLT4h6g+pzdhEdLY0+
erIEdgKgH2HWvQNDuTvERsJLGCV0l1EGargaFSgji/8m/hIxWARptyDv+EIHvVMG
LZyHKXwcOY9bzn287zMTeuQSmTRyqrtM2jzxoiQifYsErE9h9iL6ly5csD/mIfph
QyHIPCdxIFqcxRE13XEGjh91p5cWirA6zGcdkQBPS2EiXC1c6Q1nO4K47lU0q7QU
Ps98mlmQf5pdaRohFDSgE5Yvi91KmVtXhTN+kBzX7R5PeCzkL/lafoOsZUWUWf3W
2tCD6i1UuLuE1ac2wgWFOhK1/v7hegQ+J6LUVFkY4V0P/kuZ3nmBoAwVEqevMK8M
BT8W7gOglFEZainWZgTatu6pYbxSfW21JzVVIquCzmkHhjqKG24Ad5u3J21O+o6F
ZbGGN/bCXZRNmBlueRYE4p7N0T3ElzwJkhFktrPcaVb+wcXRj6NqSNMuX4h+lqgQ
0EMIUCE7Zaf4gBPS1vPqiZfOX3tQ3gu5lx4/e0iafz7mKp+StzTbu1p92F/n13kS
P0/65cXiz004GP1alaSCmn+91gODiP5RIfIa/30ArASRXqMmhLV8fn7IwG9Vq3Fq
BFE9ebyU+s4fvewFskgFuuSdbjMgam9bGOFuVCl6fddBl386yoreyYUlFyNMqLrF
gbMavRkUNj+lPBShBxZplAOhh0hLTX9KnA7tzV7a3l77ernYxmRPGwibAHXnUnRQ
NRTgUh//asiPw/atMY9nWU17PtPMYd7/PODEf+1kf2IcYYPyZu2S/LXRi3GeSvSG
DN3+AXms5fhyb6XpMJApRfrEWA0Tk3aWF5zBP5ERnrvd8G+eJU0HjXY2Fvt3cd8V
59GqJSTVuiif7KXOfQANd6wNlKFXHoEeQH0U+o4vzZBWWgEcVzC9IgEQ8Wh8I5Xv
gFkEAf+wMwoXjsCQ4Dh66cIAHfl1RLidJyqkcLp9hezQxsm7zrxn0UKLqXm9Lb0z
O3lP1AADPrHHb57ZZAVMsfmofSeBJh+Zvn1FsVm4GKrVdOBbzvjAQWBk9d+MCv1Z
dUMAJI8NYh9TCM+jcUsbtHK/w1urqwCaoHs+Onzghj+g8cFEhnStgI/BsEmyL45a
85a4RG7sNTOvbQZ+/K2nQs09VyuxfC4wX3IJ3rLL4+A881LsbMZnhwL32N5wUFQC
9YOVWmIcX12BQKHWydi6YqV46h1zZWjAmKpuNe9dXqZFDeB/Zy320GF4518HZjNv
PIidpsv4Vznj/nTZXLbrujq3uNgtM7R0C3cxFlvvoj7WpdBgFHekc28vpeHAv8bB
pFkALZ9CBpu0LokgDi+iug2I5vltFWnfjINAQpd1ZXz46tAlx16NMYJ6AYhehZg2
rkyjh6w+n0jYv3ozAwqy8m2PQbTLEXJKY10jBk2oQvKU2D+mWBERTdPbYqXnbyhX
ngvpymUyQgKYR7PLGnfurZVnoqUf/eSNqc257lRTozNL8+HKWsxgtoM3tTkoi+AN
XHUnJJGnzkVm8IpqkCNMXlvFs+ITnPq7OsIsmQIJ0y7j25DGDxZfaN79xwcbcxJ5
kTUpqWT68tqUJiNP+zH9eOxEWummuxb3jjUAjtwF1lqcjXMtUqVJZHHs1uJJfdSm
h7Hz2rh8fm7ZhiCqhCKUNI+giXrXRaMmrbbme1RhTx3k6G6y3Pdnoqy49obbBcnz
woHBZnTsv6KJHzDD+LxKjZjFeVZkkmQgJWPCGjtsotW3Nh+euloaEnazF0YKm6jF
235TgBGNQcGlW7yrahIDiXgwJhg0I4IjLhTWr4pd07JH0XSxmLa/CGgfQJH3sOOJ
/7eWBdHNrQ0qNDu77VfnXLozk4HyjM24BfhdaiI2byr26+vZwhGvEpPxGC75Ju7l
Hn4cNwCkvtYXDJymJiQdgFkY7KKh4DvPBVXdDyQLI/u3VRhw2OV9+48InNVUABeg
hNUwYyOmICvz7yaxHci6eGLOzHFcfJuMmZI9CAGfIM/uidNNaHnaGYQqvD+dYNbq
B0X8WW1WuPvrSyMoUpEOWWHVC3qeSpPU1KEjlDX/xNH/fMeUCSb0zmKafyEmLSP7
yu5mIpi/rI/QLDHPhZ4NBqJrfHf10l8uv8pqz1IDcNDhpmItb8Y3zy/41JL2qr7L
QD9NIewwdcVkuZwdBPksNsv0dxyfYdHnDW2eVn+Kw3OvSTMDyqbZrzZ8YRzv7GDb
bXXkqxEPH6jhDCeh0GpyCvaZjdAWE5Jx+WvgyIZyjt7FGso2uQNUTsScKRgEnPCO
SA7h/4GFvYTQlFZn4EUKAHy057ytPfDdr4kCSlBWIOno4rj2ep+7ptAJsSJU1p5l
iKfmlXc6/MOGr+Jx6e6HUmn385iWucQglo/LdYvkT4lTvThsOhkQ8Yk+0stPv31q
50KIqNlznYH5o4YVGlqwhKJ+cVKGrjzPZlIECSN3ibcpDciZtiEK+s9HJynlmpUP
Ej+mGRLoXZRqtilNmJkZhtgDseGNLApLoSDhyEH7Hp2SOP9Spir+0nyPg6VJHciX
Ndlj8UIt5QW7AaVkCQQe5v9LTDlEaz77f2/gf1juwgWw1yUiYdSmrPk921rqsUux
RiZP2NNeLHOLUnQVviNQS80AU4DRaqcDzbbg1EuyXDHHK4hwmLfM6dOTWDqjgRDL
kW7fEqOVdYfHEItvkwKC8qHVFFBwTFsUW2OrtoYcu2C7ndVkKJZOWgO6bs4yODb8
+bsCtZd20MTHmpCIwkjbi9vw1sKcV5VtLPyRpoejNZQJPFV0LMWr2IGzvHSpFYEN
MG0ur+62597QAwarVxRQtlvFWKHOtQUpN5XzltrgN1g/duL9UeYPzTFaEWyYnYr1
7ugXqW1+Qrdw71kBtwcdF+qfB2GfjV3ajn3VyDxo9GLIJD8zrqW+bP2obIco9Etu
of8Tx0pRgMDREnn4JcYVJWWEZIS67+S2NiuvZB2N9bqx6VHaAbPhw1izn8YRGXvk
98nxOEkcg+l0tBnqklReoP11+FjSxkvCB/92uTnOW7QAebMnBbJ9GU2zdd5agZgo
mw/3H1PCjezHzdcJDgojcNHI9963ggaOqD7qLom7EJ+70VwlMPoNBcrKQ82+0wtA
1xDlB3Tw7afn/S8Cu/f+fdwQH/oAPA24Qk4z1p1q3k5dV7kwb+TQtDxdAZexxs/9
24xUQe+8l9NbT/o7nfOTWRgheUGOce6wrMHuULtyvFIsgNL0dIWpr+zmCRU43nul
Uk8fEhaUg2gl+se7xw5TQ3PGVbI2OeDJbNzdvM0xo8u3kTApsDVxQhUvI+6/Kamp
816Z70gwaNwoBrZEsLukEfdz+/tIQgBHF4AbMV0WB6vPh0/TTIoboZmhFt9tk01N
TlgFNVq6iLyhnv2P7G1Ob66kcrlD0pJdqrBVqZW9r9DsiEawsLPrxJDFwvRw5LSD
1OOcV1Ed6gTgcSH8+q9fGSDpXlq8ncRL0pFYB8LLgNv897phgat6peXqb3NE9r8x
GfHSra+pI7nz+CpEFQo7lN0if87y4NXYAkJiWIQ2KkBiMO9YHErR9DrA78Aq3hPG
i2R5dKPcA8MWMuHn+qaoJ93qs6oSahXUgyPJ/ZwSzsMynIph2I+FzYptDDGdy9G3
LWI1dsUhxHV6Ch88eGZuPuFI5SjIdgKy5Ndc704xgtf45Ktauctwbxd9H9RRFdzo
2dXu9QrKvYTcl0pt8zA0ko1U5aiBOy/b/UMVH9/9EuuYACjK55wUmK6cnhydL+uS
sabEyGKB9iC8wjz2Lt70ljbQZDQ2844t9T5qU/Mddqt6WXne8v2mDLCFcKI9kGRs
cpwu6EsNtI6GXHbnPOvPEv45u9fiKJHdF7qkK2vFvXM3UUFkXe7T+yqrv5+AncN8
bg6YAneA6jztm9a0XT6JWAgbsEydlszTOPttaGHYfd3kn5pjwCvza4/7L3C9ykkU
0ZGhlSQJ552lgXUG8PtzwNlwhLdcMK+b1+HELZCCoqTehGPo9yDtLwT0z1LwUwCQ
TmIN9dI+pM6Ll9Y2sAy+q6Z7LzyYJej293pjJqHeL+epaH0x+ycBljb8UHQ2MBlY
XWmkREgDL88pO4Rzbyaq6MBF2QCk0CiiOVp5E63XnA3Cdgff09i6SZQQp5E0DKlQ
3BnYm0hUDpM4RVN+P8Ls6Rmq+p9MghanUe9F+n3F0eXJ6G/QzWtYPCY1iGtSYtvu
z40ckQX9SSxmmf1IRoMIsq4mGoC92ixhtzj/w9jPOBbHuwOMyCjRy1a4bDHLGxzq
rmvkc6Pyzith82Sp7MMo2jFhzJpuWxhA1iVfzpgfpUlwz/nEQCJyVOZw8Ib4RIZv
IgY9tmZ3FIZtqWR7i/e4SqFS6OxDChdPm9tXB06iZTTE/a37Ra9a50wFF8QIE5wX
xk5lwvCxaQtuYQIr1yiqo2DDZ5U/j1rTWweSmeT06JDPYqbSFklkVwy6SYdGBLLW
iLsXjP+8t43E6eVLaDtFxzcqWVn5GtBcLsKtse6/n9B5bQzQ3kdOvJJq9w3x0d5+
upCsRdnkAuJtYZKCX/WSemEpdYIE6sLHATNps6y80wq722l9oSzvc0mWmCBjZLP7
UA+dSGJHawVNYZvcfKZ9inQBEFOTkArdBfaGwS/oUoLmdWChdxrmkvMr7enDgfnm
zMBLiulGpG5XbGEgBcPwJScYSp3dL59RHfhazHi2yMxmn3967+SBOA+Ls/IdzOLO
199Uz63+vp2vrL2iej2+AezC/xYSF3yqMXYt8ADqr2N9BD63vbgFo4dTgDDIqEo0
8IFF4OKrFxx9ipCjan1PsptvTi08SohtPf2AtqtY6DhgdzWA1jk6/LZ9SXyTddY0
K1gGrOewhJ+BOQsnhPis+7DMS5GoFdTuV5BqUm+U7k6PIawuyRqoz2X7iIm9Bv1i
yN1AfKZ/BFo8q8kad7NKUUR5LkjpLLcAZnP2YMzgzIQq2PxRNk4jpU02ptn6wcY6
fQrU75ulqTS/HY7H6QHCoh2pOdzznBTFp0G34jrH/GjDYceFio6i3bO4T5SBjrhT
Ld0yPPZH2qA37MhYIr25D56JZxcrMZMItonZVJDDJQg8XBRDNJbAnsJmN4glWz/u
OVGeURbn+OTOpl5pLhkdygNo8QrHtvViwQ9/u20MeShPxt6NOgJVxivXiUOxxY3/
svuAqv1GncykgyJ0or1k4AC0Wr5HlqKTMEl68uzJUFGKUiO5wY2m6joVJw/S/yrY
M0Z79sAgoF7WtdjL2l7uOsLC/b+NG3oke67ZSkYNyZ1VCXg1kJaPJi5ZLdUgxMge
/GVvnfh9FLI/s8XZuWWmNXmqPKZgwuAwB/q6iqpidsV5vNWIZQ/2ESRSB7+D6W5c
QU+G8XozO7QzPcsKJ4+i7+k/xTyVyS3bAHUaKMZMZtZLn/O2HhfgRzmbVr6sG8Ut
V2aokEUeevoRIwQy9W6UP5FV+i9K+uoLZQq5MMrS37h+Kfazkj/443ip6C8GDl3x
dLLhztYFOHiKRWEjxMpm9I2EuOaa7oVT/WLk7/FdriwIByLrhaErUY4gEFnALMsu
aDDaK6KwNAEFkos6WvdjMc2umk5L01vAQd5f61zcc6LqXBW8VlltcezyGv5mveo8
W2GD0O704pphxfn4jMB5j26h52FzpprLKRYE9Ra4CmM2NuRIkejhWYBpmylbqdo/
rvwDKmsYwjDfnsMCfOJU+I5+HmwheivEr3IoKksmJ1RBhp59QD7jbUwpFoR6hu86
pbGCrGQWgViRAfGWInHOx+VT5xbgp7Bb0CZzI/5LwTPv7su++VdQfs0xuqw1b9wi
fXHGvqfZ68g/ol/EMfoYqjFIqFFRZxY2qMeUCUvYck6xnE+8kIfOaXNVSIBosYun
zZR0iN2+aV0j80NzzrNRnhQ/QFvNipVBvp7IRczXHriQWLYYQkZGq57vHhqKkpeT
j5csxuF/7aBVRp0mGmj/GeBab4z/AUeiLtrGA/Q8LTHBqX5JmeJofB9jxlmtiVAr
EsBcZl2hl+kSU6EKzMk/Hcl+C1u/xTNoWrXdjyMpRCBX4bzFzATbX4dJ1QXrlde6
Sk5VKhmQiPof7rfXcXAMmScnEnl/fmmR51wZpoZXk/CcETzsZZlVADJdDi1aQfA4
QIcXjDokGp/EKjqh4+vpjSEmm9foJJnr+9Q02OmjtB1pl9pXjF2KP8rJSvlvCEsy
76oOFQ6fJ9onjFNbt35TvfkkzJu0ECVVEg0/aQmZ1HbcofhuZqhyLKspqGs8XmFJ
8R2zmxnkDbYAwAWpNLa3X+RU7qnBwHxQeB/zxcHQNUasIr6q2D1P9YwGpThznoaf
PyUgCBpdEDBnAGNp5dFGR2Hs8bx9bTVTlvu2TCGQzmSB5ZcLzOfVRxqlUwK0yl+w
98dN2adXn2b8OBfkdd1TIcV1Ji8THFLi+qFFjw3sYEzap4iuxauNSTUAZUZEginY
ue8TPFx7Bi2l/80MocDrH7Op1hB5RMwHhHkz5X4YfNpIRvqxRLrW7FSmpiAspNL9
vdowqvGEqVOevynks+x9E+NJaDIIvnmcl78AAG0FghYcDYhwyflt507fITc/3aZY
oO+tCT+8o6eLhvPgQbSvVFyNfO+DtklJLc2xlZm2NcYVcLFbHc4WU6FbUxQuWVKj
IcFLNPq1ldeiSPDb07J33qXHzHYYJ/nKyrb7Mm3MbJZQ8AHnaUE+ZQGaAh3uFTev
gjY6mWz+jb0pmm9nAeLm1ihvK4NFyy9LafZyl+SpoeIMOIQJNOvVakF5rPhX5bQO
VOf0al/+ru1bbHFIEKdQJG8xXi+CRUdg+W7pDxFK9IsMMwdE1fy/5cEvZX2C+vnz
SOKPuBWZs19DMCvALSOYjbQhUZaraLS7Ol3zb8D148+l0ATl2Mul2R0k8SJXZFUW
RY1lvkMh7bBjcfExjPVJpGhkFCcVjwI2h9CsXXSHfSFp4txhTcFPch6ZWrHQkPyd
cCBVDyloARfcCPO0qDzSpWkH6JiTbXW9VdIulaTrssstRJHubtkl8tolqo8QkSYC
iUlLiXFqt7aXGjczR3BJ66fk3emt051+M+PlD1dbPy7/lgEJLYNbCcA4bXQjs5L9
qlH79vxbG1quUhRGmHEzJPOE3OOehL6tR6A3Ypthav3orS9GR7FTeiF8ZcEDfuiI
xSus8VmkcDYR5RVKw8CZnTXcH9oD2LnqSt9ZYvcydhwPeixZvizBwr3jM3deBSyM
N4BbnKYZaxYyoQxYXSZHx+Rr5RrItuvSeBmHNWdbliU7k4v8hvKWBah/6B//FAIs
RFM6yPJCfIGg6h571Z+gOlXmMpxjXwkIByTi4eD5oxxNkLvAvsbHPM07zQxoNVD2
kAHCiiy7xhXMwWYFdBYxSpJQaLHTRZ1TEB8U6apdjuGLPIP2qneKGmjgycPdI4T0
pR2QxWqgqCg2kW0xRd0hnv5Qt8I/x02oGY0GgNg8LrhKcgmPQUMexq8CSIONVloX
hzszQmUttSgowrM264xSGoGxfWrs9jikhr43/UKvEqqgu/kh7I4rDOxe34ng6PsA
mGbp1Kr9JmTX+C3aVfkj6Lz8RwC890xfg/kXtVBqPhMWxBIIobDVtAAC3JJi2WUX
zh6bfs8dFhnC6hA85iwnZCLc0r/Ec29bBiNZioNM1BgW8sgQJjMh/mkg7qypmCoi
b/WEnTis/RJKjn70Itj8yzfMfECdPzyZKuOTknHemMh3xMtmg5NUC4Kd7PicRvwd
BVRiYD/msgbS5naLITQwAjDGI0IEORIUjwgO+2uL1lXtvekKLOGClnvBGHW+GV5G
SrlOGOiAlbIRODOB0PCmcDgkFYUxs+XAyCvhge+1Y7NuqCDB5UeTlhSdvlcloYeJ
joZh4O5EYq3IA01/6Seg6AxSOltv9fwJYvHkQ0kXR/oLHDRin91Yq4lEX4RmDt9u
veSbdBsWB5qtlbrBE9JDwq8/TKOWOjtUlusOWH4+zNNv6zBQgTpUrNgYhLJC4haM
HYo4lZskV/7IxT84WGdpV8mYieNmlOM3/KH6IC81H5JtgOb0VnnXQoHpnbg1dnvI
p82d8u/uL36rKcJDcIzpIKE9a7YMS/CDe+kex+6EC7Hh9W7ZpMucxkl3v5tyQEP9
qCQPhq6aN+UW+umkd3J3zNhJIJIwqtJ+FdDPFL3yceXHnW/P80EZVJjPcu0DUIvK
MMb/F56vP2dEZSaR868UaoCQIncI5esT34wgWDr2HDYZ+2dOZDHB+1xl+cOkz6wf
W2iXtOPS8q5BGO/JFGgHYw7xRU69EL4CRkjDzY/KC2ANkTDN5wJaIAYj909Zjfrg
g+pGTXmNgD/pOuJZx9Oksk7m4BI3TMCnWK69NsKC1vNIXcwMVFax/VIGW399AAqM
npKsbV0+xR0HcAn3wqiaHA5W1B95OHwzpuadVzhZpSZ3Eu1q7yTlViIkow7sWYut
29CRk/97UtZY5/pX61WNAgsnFvHk+rRRU7DVisPULstzbGHDLpt1TuJ2ZCWat4gx
ypp4NVhK9piLL/BD58lmy/8x18eV1jeuD+Vw6rbulHerSqcHS7aLdOtbzUxBRGml
lR7B6qOAxFvpCV7Z+BDRtk961lR93LFGAQcnmYxdl0TQKjp3QtFmSW4OSG2bqh/k
fMwOVYQDC0KX2jSyeTJ+nRsCpJxswYsHfjaq23XVMMXpTurstT1sRZsj8z56zuwF
CUxRiS2qSb3p+k3CcuqcAElxoCEMkNW2u5l1HT2wKNKxesWwQroBiCtSb+Y+Vd4P
EmgbgI6lwSJDQzfbkV9YzMHaSju3ZzStFwSKUq3baYWBHzd5p7ul4k43oqDrTyzL
N21DXpMIDNXsFbEeceg3Zfc5mw9D3Qfb0xHkHyOPf86OKvmoPg98DMjIUX13NFBF
WdbFw1RoQeUZ55iD3xngtYgdStbbYJMx3dPiBK1eMdGu8qfVilHHad2dmLIkvbnU
wrn0XCDoxlcK8MD/xoWhJr4rGeMvbJff1+TofD03ycaaebFjeyq0b9ARkRDTJNNT
ikQax0Qkw5e7peoglcaO5d+dFTY13baTVfE6sfQhmdvlcYB0Xv1dQl8VwGbVOduB
xTP/Sh6TBckFsjusiCSpS48AGPCxhDdRBUaWH8kc/AhPzr3ebJpsgxr9W6JixHhu
RAERswnxY7wpckKta6XF99pemE0DIiXeNylxXq2ku+2UNJrJaSkfx16rp0pXWENQ
4moONNbknB327lKWylnvgQ9usvZ5a4Lh7iTMVQzW9gOWnOQJ9urlywBqn8m5wJOT
1K01KSh3i2DmNf2Foq/vMUV87WQZokLsadurkFctBzoItvYEf3YCcLDH3+b3RnpU
qvaN2qqOj173E6FIAFYdui79eMYSrh+ks/6NtFMaf+fyra4u/2QKKBw5gzEc3CrL
+lRhpvM8izAgE4ReGaUZCBx+5eUo5xZu/CpFb6CmUvssQ0B4C8+j3xwuRS+5cmjj
YoxsFMwF3Co1QY4G5upAx1muOa89B6rOLkA5oxPm2uPLcIvM1f+P0znOBY+jiUb+
ML2d6azixWuFh79Fhcr8TQcI+ArH+BK0SBIkt0kNlbK4XyPkjyPsafyDEWQ5oOsP
U9+dAMk8Gz7c3BlU+hmXtArqeKmx7nv/eHdHoK6N/2VteLYr0Z5WyNSJ2+uO9V6q
3HqWZy4E0zPGVEy1+4QTvUEY12EVCvoZS42QwWeTRgXHbqCSeTcFouBvqZt2Dvp8
KCA8Z8VXu4R76IyogmQKW69I11dDxGJfEcwcfefd+xAdfY+36be2ByTPi/qS0X6p
OfHoKE6+ZrSUmcxphcEFfpQGA7pFSAaJYaYZVb5hK/xZV8CA+UoIcPNNG5rqiqvx
qiQQ7sZvBUAsJIRFtErVfEOklXHKx7C80bUnrZnPm5uWHb2Y0AfaJHrmP6oJ4ZgN
BBBJztXvTlVUhLDw4CfpoSaBCrVgP+aewcMkDlysl8YQxqEKFGPCfhukjR8mM1gF
BdjkZ3cXp/ujUxvy1b7UCUqbbONlJamv7fgSw3OSbOEdeOcK5/8yXlrzsPJ8vwBs
Ffqo4DAgl64nATdAtfHEcISXPU0mn+XYON7ZLVpJ0h70IZyHh/yWW6RlBOt7BqLP
9ypd9mN/ogk5x+gClvF8nNYpMbMWz0laMPaA+JlIk5wt8g8rw28jB0coDzpU4XPT
q2Va2bFlvb/5GCBcHQNK7McBMXbYyCq1fE0Eet63SqGE5jaIKRIRKWRWl4MpEtN+
7JppQSATZ6hS14M8VXtQbIFE+AuBOwcHpUpLf8FadHo9d5Z+VSROuQx7Xn/aAqC2
c2vRZ0Bw0X4KS6pEUgKE/aQwFVeNPOUZMN96ykO8l7aRZ3UpPtWJM+rRwy3TE7Oz
tHfAJlbhaJcvMu7zM66OemXXw/6H4lHIjdWMzKOCXRW7ohvwbyf9rkQ+atCVKfnV
w7tLUevKCCxxW8kyWF+HFL5/lcJ/D5AT4C/tY7x2DfVoTQkLXb8FD9c+jamPMWce
lanqpqS5jS3GvtnRZEfTx9+YCNtWqYc4rGxvDyb613JbSjAUmSkq+MOu7pyCSuYs
a/xeNMmM2L6ruuXA2bj2N3ethgRhqwk06+EQfFnXE0w=
`protect END_PROTECTED
