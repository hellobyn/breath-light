`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlNBy4X9/b7aaMv+4hRQbFyGpMlqJR9HPvOHIJ5Uc7Tgjb6hFzBKxt6G+p6aLnLs
SiOR8Lt1myUoKQXBRysesUS1t5cH41GVWsC34fna+VslDKWbGzgyIULIXFi0RCB5
aYu4bpkZZZ75X9+0Fn+GQJV/Eg0L1pwan8P0WI+dRV4uA/S//oMsujSXKyM2d8kT
nQdQdT3nYp60gVtKQyVmvZoPsvjEycMQMvucjfboj1dKlpobSBk8BfYeGVKG4PQK
hXDLe3dJKlU95RDIZSbny8bHBQPwAaduhPf262XMNnJql87pTjslOjrjS3M5xiQh
qTCimU4qSImgP9tq33B7JHOZWdNAvrZMaDFrzG7xAFRPdFwvVJZJZn+5w6EpXE89
2aAlJRxOeb8Wt1/NKdjFf9PhP4qDauLmA15J0u1CVJuumQWLI7D9GGIK1gyPVAIQ
tkzV9If4ZoKff7HaVJBRdzcYmYLsGdgO1Fs20VrAy8bICxqpiZV3CIaxxGvHBXjz
V7lyhjaET4tIdA0vi7+SvcdYT17Vwipe4M+TjCCH/BTSFu6O1Zwh0Mr1hTM4c5BO
x0bDRdi12klP1LC29fzs+8Jla9YWnHvNZ+0YYEKPeoDLnRKfyzyzdaJHPRBJgEWK
S5EGZqV7aopqYdrT6RK76XXYH/a76eFcd3cxN9CiuEsKct/ydcXIc4o0FVYTS3r2
yeRhPpNO2XguvmHh1IGKZD+vfq6dqgUI+tTZzLqxxXzsdmJAREeNLMizlm2SyFDk
9R5Ew77sLaTFRYeirhNOufxcApuiHglKxX+457WzjTg8vFpBQcnMHq8Fz7L2VbQK
oN3MoAXrGlLP3NWI3ckPQStXE+Y0nuY4KC0THDW6z0jYMmNyowBXc3Zd3kw12n3g
D6H936ENboEOaSuN5FXoNuEzkwry5C2cGCzYEVMwlEC688YHx5CZQKGgxNBNBVD1
zo7Q2FmCYI9etd/4G+wMRCCiADF4MzI4qPlxAj0RXsu+th8FGBiePiFtDJZZ6vPZ
S9mwwzfylRtgRV8RvQx9vwzbqg9oT79YbEPV2qugYK8aBJWqdriL1iHjry/x9o4U
3mlWyMG1qXkk5REZmnKar7BfD5GBlNuSt5iGOBaOWD+yQcPekFGKwGF3bZByp2+U
cyEtOhVem2HiaMrz3JG88bn+gWkE6jXR5JZe7qBHQCydU6w7qNg7kpTx78zeaP6t
03sMFWsm5UaYXJbZeUA23SNc/Gv3mFYHbiISLmAqaCoifAXHTygn6gkuJAHhSibM
nJUS0BK4mLvd1hAXMyrRpEA4QmK2mgX+iAPd7DTMLKIOSa2Qa8ztSJTMzwtXsNV7
Y6yjjtIyYO/DG+rSivovkH3A+Cs8jDmaMk+B0sOscsBoYzW3rLnH9+rHJWhPeBIN
I0uIvk/EqeHa+arR67d9h24eVZWFYSHduGAkgnVMKu48UdzzffBO7RmNHMDHpS5h
7le4twR5Q68pgh7jgsKnGQvb/pQXPt/zSp80xEbktfkRtf27Wio77CWl0cyhC6i7
YlaPchp68AXFFcEOrTaZuYxwt1ADLNeXvaTCcBWJjFlDNjRppet29JM1NdnNuGse
tpWkaYXIyXgXUQZNUWDZHChPi+uxXfCN82r85GO1fFsizLuFgiZLGjWN1VphWsIT
GNKfZZ4cI2kc6A8agBghUpHsIOnz+L6ZYPtaJuA0zU2kVPtj75ENgbcyc9Fck2Yt
k4PZptijH2ajNV2ty9UkcGojGE+Olv3a94DBCSJC2hWjpWGl1d0qrvBBIrmI4UBy
4XPqPbDd/A1IF4baxuSYYvsxdP0296tBWygTz4C6lpzY8kedSsPkMTr2Mf2kpf/h
gQx9zdHz69oFcSTztmtjq90/yr0eRP/gG7S+pKc4nkhk9IH+Abxiw9RIs41MCkGi
KumgukKt+zQSHIXZpRsybulj4P6t+XNP1dAX5MJ5Quu3+135lg94FsHQogDWuOwj
bHYJjlCOA/WWUF/7FUqrN+VTLtCnZXDltIqf4dCXz4uRCBe0eMPuReFT8mKmRNuh
PjRmaEJIaJfQUqnux8v+8ikrnBjI2PCBmFqCuLLL37+Q3Yn/sv37q5+7qSW0NFIv
dgidHdLBzJwL718THse+u+MN2dkcV8G9auwWapaW7h/vrlRSl2/ScJVltwOci+CE
4S9Y0uSKE/UXyM5wYZ3cBVsGXUDXTjhP7Q0FYOdEmaKGR1E46M51b2rDaSZiQuyf
YBxgXv6RXC9oTfNbjm3Ah+o54D79KCCbjrEYlyQ/5z4dl1Co2m0a9Z1xNds6NNlT
n27u1IbSnoB3adgdTTWykVCuconCtG/rdSUVVE5wbj/XFHkceo0EM6pu2/8oZ9xm
pBGn7Suvbksdj2weyMNaaHdeoLHNKzKkg1QbdmDsnQvz5GY50kE76KXFvZpJcxpq
wNMPcM5P924UluTuyj/e/A1dp8TkFuCQFkUuIn7czM0I8Z2kHnP6Fuiv+RidS25t
xD2rCD2ILPIAi+6AwGlICT4sCxNps/Jdz0FuYsQfKmn0ITL+AyvsG9FJIio+9aL8
39WOG0/eO1TVO1lrXVt1Cx/g3h7XZrxGd6CulkBmczMZmQ7BKoteONyermeHJUc8
rSJABXIUnOsbsd1eHd8RmiX1Etybm85k0DTRaFsh1ZZIG09FhJ5oD9an9yQOpBoG
2P4dxE/ZRyemUd0mQRoXzHZxJwBU2JLmjqjoEaIPnEhB4IR4Alkof4iG5X9VmM91
dGomRcZ2c8gKy4/6zgHJarquKPisopQjf15ogCdr8l/+ED24i/1//PGgpFANBHsn
vw/vGQQiDWT1gV6jcbh1fYDRTLougyQaYhc+TjQlmQBbphIMUvkduCjh8gNpQ97v
LLWLlj/RZWuTcrMr9LZ4OXMkuuRKfENSLGdcB16o9qK6HpFyPC4N5AG9QePnJon+
XD7rhFDxXBRVmGcApnAcbymes20G33bILcNyqebroiaBbl9tH8JKW1Ldbyn1k6aT
jYbfbdHPt4PWwzaleLUCiUr+tFvRLO8SmvIz9UgPoyr9l5A/XHKRNsWx4dpFO3Cq
1ZihmIlcVskEyIPVqbFg/jt/C4wjtbcyHnEpDNPOo4/NJgJCqDXKo254e+9qjK98
dzDoRysjo4c+e0+DKEl3M5BlJVgkBGmMhj5Ze9jXnMe5oOIftIhiUSb/sfsYfUsF
Ddb81aW967y5uVwiV48+yDpH0q+A6zhT8V3Rucpl8IHtLC1XGzh7rPXHguVeft9g
O7re1d/x0xL6aT51OLwEqN9XfcHS3wLLFwlqngO+AGqYoICtoND1q4F9wD2DcT+V
CcBf6iu6G+7a3ODzbXKFSxjD4Bra+/Huy7yET65eYq3ZTkN1DkOHlZk9/61MQpCW
CFXkNU4wyA9ah5IhLXfVXFNcu6JGeI5DJ9XhIbaq4DxFcA8rugCEg7kS7OtLOk+x
p3R+ZGzzmUIxwa1dCJqDHwgvDVnD/jwIulUQJNCIjd6BsiVjkFODMC0PvkjFcsW+
3C+r5lpsHWI/hJ9+Dh7WfcxLQLa4DAY0F+xwRjpQsgS24oWkO23eHNQtNRQDRBr+
iYCAnZcvhBIE5Y0VvqtUkNkbmWpYbBFt66t46HgQ4qt5lplH+xvn47ziLvNj5LVz
mJ5/S0FVoHKzpcYaF+U8oQdwwZeDyij/YdJXNqDGM1a8k/6ULUQTi/MiLT8zx7Hy
x1QZaLzXjHo87Mgi5fBjR4vaKuz5FsYwM/gyvGsViXBTFIWugVhyQynpQfu5l9J1
6TAyyPJH8+hm98MHbzx2LVNxHPSfZgKCdIyRitnaRN9byRWBzTHChyDko/gYulLE
Rq3bjFyo78J5N/ivCZ3Gf4p+PisTR72dTQa0IUA4OUkHbHdivYACy24+jFFFh+my
+3HRyi87sdTKW6D7bqTv5YONFWy/QZxpKzsoX9t/k1LKSkBPO76zSrs12Op8PYz+
/fkx3yw52IQYvmKLFNmjpmUVP1KBoi79DCJQuDUt3kEm6MLgHiRr5NGATBRMktyA
UOtIo2njg+G6KBDBE0d1kv2zdPmwdYwlYsazHmr22yRm9D25FbkS8aTQQF6UQmog
31f13yHNgjIpGKv98f6Ro6+Du+4c1w3iWnwdOZyRKabnaxLbIA9Ue/PhTlShAW45
3FO7TgSnU8rd18HaZAdgsnvnP/1W4kYv7tJXadEmY9l9kpPhAK2rypq/xQd/CD0u
VPoOcLgmJGYLLbUlNdqTL20tvJizawR6uvQJjCPRXOF9BKvSjfK1ZoeYM6bUULgr
4IGNqHQtAeaCo5deio95fYf4DyUf6wjcrXjHlhe3G2pZwjWT1V0IRyhm/RuObS0P
aT2Hrs8yl+CjLC4YqLEP12JpJLi7jOsTyC8FotHg26Cy71bM5dr3F07ZgwznfGDZ
P8qf8o2nk7W3XHVUhKzIHiraJKeCJx+BPLrDf+DWrm5A/9P+RTjlNOxp51ESUN0H
0TiP3H5NP3AAkm5lJGOxybYhzcIWUFqEX7dm2ATyhlYQrkQZA4hiX792bnAS7Lnt
RxRCAocvmhGwuG+fVdjzEdYL13RXwgihSedSqN+3wwi0aw0uqbIESLnKdDC5LrBo
Ss21zcx5SftFyh0ECQFNXBQp+FvrRH4MlKLWsDCroHvGca7kqL92XEiMeC4HIVr3
GnshjawA4IDpCS16FIIm4VZJRtrMeFS8hkjy4YWp/OYrQHLyGFQJ2ZCxsnoePOfL
4MUCW41Kow62WXeyw0ct9jEvy+qPniNhxbdY6eoFCtDPDcL3+2C6F2x38rYuO5lA
ZfPQmwb6yXeMlNkhvilg7nGo/WMxDSVUgrvhEAtPMeYdxWjPbRcXQOaFPNFweRfP
Nms/Gr6G4AnYHq9qzMkofcfbfTi3+/tlePtt0kocAYFgBqGn0U8ZTzZkXtVdlsCn
rOi89q7dAILmtHOHWCTY07/yZHcaNG2fHxyChif6C/kNfl6LaP70KLluiCySvRqu
xErbrJqYAiugpcR40DfnVbKVqE3487u2kl1A9/dsewr43ssPj5lkIlnTmaZp54d2
ogO8LzQIwwKjkyKhQLK0TPygzjGEaY+Cx9Dq0DJhGXdSXKghvIDgm3ZzUTte7tRK
RhjjY24+/j1+AeHhLFa2FytMgjj3aoQ7A69Q4y7+l+W6H3TV9rVZgTikV0P2j9C0
mwMBPKbObhu9VEQqDaKfYkNF5XcnkkFcsbUJq7Ir1tpgL9eevd6q0Xybhx8YfJK0
RCrOeeUkwemoRTYzDuhE8jZ18B0KqZTYdt5mW+qE7mcfz0Y3v9YFSvGMY7OLIb3G
0ti4qXtbWpbeGGBTErALb2/WiOOLeRaAmJQDAxZ/3x7W0eU2xp3I290dYw9ZRNRG
LPhIDiMKVQIxwDjyKvfld+tTCuo8JckFrbecMjA6LA5HU+XdyC8W5e/y7FfHkCIg
tq4I4X1tI8xCWssNK6GnfO7PjPOkFA5ZHc2GDqZKVJq+Nbf6XA+Ngd7LKRvX8/Wi
9HzZqe7fwhkvapA1kYLC6kJ18V0RiUM3x0UbwtQvKYkn27y/Q5+//5yKewsr1KZk
T5Sh4d2if53+I9mZhDqrIrI+xxi2aIur3dcHMfMVVftdKL+8qZbGCDTRhXnDP1so
W/yDLMm4NQIAEXXesu/hQD4IsItzTpLZMHBo+nGxe3GACMmC1N2SENFezd5Ygkrh
u5G09JKbf7CEHghcTHCHJXacrIO6Unx0DFeTWdHsJy2cxkdVkJDQNx5f4zRuTQjf
KwoPRunsCzbdAxkoo8/ztvriL//U+QTf5RQQD/lj5WtH843KDKglywFOy1Omqbqg
/CPh0Jc9YkFDsSZjfXKkqO0N9+kPoKlPadvM6ELljwcnSne1/SqmOIilHK99C4LU
1poJ8WUz7QQ4QTsHh/UvgqCb7B9xKHIOSlJK/RRIu38TWvwqB79w/aQQ4RpFI5dA
y323huIt4NqCFqCbdu/bWZqjCU2+al9UGcTsTVaE9+RHQ/06Ij2oTOnJheajoZib
AElpI83FavHxMGsakUsMeOa9e6IUKHx4+YU21HWDfE+GUTvypolXZBbHKWe+fo/q
PlG2yUBv75YpGktDk5h0jNP3ARadPnaXFU2Eb65XnMH0R2AS5xlLb2mtklQCtgeI
pEW+iHHdlPnp+6zQ00Jvvv91jAr6s/jqlsm70HV30gpa0zMkr0QWGw4l98v3upj+
nun9e6nwFY/he7KI9LzhJ21AA0YGwRW92vfSxsGPnDYQB+VzpGM1TXkt9eTejQNJ
cZ00URoiaOBd3YcwOASBbCBa8sdHmNmMUXPPg8vH1s18Tir4hSOvD2wiV8fQBM60
qUyhI7FULp7fjSjw+LyYt7nYUAczY37pjt28LMZoeaRDtM5iS7mV7BgOFe2WcK1T
jTMI232Ty+DHyVz+yceFawoEmuD1yWUQNGhj6Kl8dmC7K0BtIO//bMPpJSjnN36p
uTfaUxfYPYLM8DmNZFUjtEhtLWQ52laJiaKspWhK4AIbZ4m8cD4SkrG8ksyx9eYJ
7WCPhAqBKNgcjGWl7vyOu/3Mj8OgW4bHUVTONzogzNsqw511WQdaVQHKGeSzSxZI
nDnSuPHBJGXnCuw2m+vFgk80ttu9srpFBvrlskSi7aFZbkLpgckkAAL+lACUFJgd
0G7T89KgfAYNhBB0ZuzuLUWM4vIjTCilsgX8ehZTOurCoBMWy8uCR5XUQhghOfpr
QKwCq07+DaKESgh0VW8AjQ==
`protect END_PROTECTED
