`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bw10T/2WP3Ez9L7GwCzdwRXU4OMNHChe+XBaL1spoRUeKEqUrZMwDJ4DGKpWh4cV
EGT05ONnzZgCIf/AwsEIx17nL1rVdYMIpxeU/b253LR2X3yaSuRIZkfgObGYrAqm
Gn6vQa4DYrj1EnXxvbO4txykxtQUkvCXIenrGqIn8LHOhdw4wiF5fY4ZC4QFzei5
p6kWOjAHhRjlCz32020sNZ5o5rKEMnEE2IbYeZ0l8J0ZYCRcR61DvlJAb/KwElLk
sjVYv6EGQP6amciz9Q7+Cq8WUPP8Dw4wtiB4wa3ek+pnVWfFLd8VclbCRyzE1Jnm
1/UFOwUcKa5NduEx+Tmy4N9jbJFcB+aBcHki/FMJ8CsW3ajrWaLKjneX5gyvOd6r
cnOVfWy+GM62sevJgwXKEuau7Cn02jUSpxP//70T9uJeZ1AL0fPpao3VrDg2t2Kw
wbe1I35YWIIZGCCUE9iQ80zXFMSwUwvowPZWsahgFqfSr8YLWT4aE0o5/c3JdRE5
AabiUv8b6r5UAVLb66S5PBqQftB2wzZi1q7TAunryKd5LeAPHCMtNdl8GoQHLCA8
Wwxlog5aF8MCiwO641P4DFSrXNkMS64Hu/E3++V/v2Eh+xGGcx28Ye9qC1Qyj94z
gWta1SkkmsNbYnQqelFhh/VnmFjVaZ7o1zxP73z5i2AHELeFwa+FK4VOOo4ZXPy+
9Xt6bfD4WyH6YNSK9Y8sJmEc16tHKOVkVZ80B0CUqGMSZYjnyn4aWTll+Diwz2jd
s92HQVQmA+xo0+jvmaTbHU7Sh9r6VmluHSywTzrX32ahKxd196c60cLd26v3cDmr
bskqdCas/HdhzzMtNw6Sobuyic7oCW2DrBd58xoC4gsy6V7o+q91Pqo1b1HqjIq8
ixvlHoGZzW9cYmRo2hU6NTMBOOQyldoNFn/2gkDzPyAUeB7D0xOgigG37Fctz90y
NwyICVagKl2ntSAimaySiHzok/I4iqO60ubwhJmK/ZIyfna6IDIjQwRvZM3hsoNM
Ar4G/kh872EoFqRdKHxbrsxSfe4lX+MgRPx9XUWnZSPP8VW4WLokNck4qdk2WNS/
Vedj+nTDzqVgcjzzAOjFmZd6jjbIpY5dZcXhz51J7LaZ2GTCN2wvrSEiiAh4N+0V
i+7oAAorzmoGNiQsyD7OK5hnaOUoNz9PmtedyQiN0kjW8ZArMO/H6O0Eaganor/K
2HMoAs1mUBGJChairzYrAOkrTUu/1vG2eCRnkvfZjmo++iVdtEEmdCqbGs0uthrK
AjFFKkaYpskf3dmPmWziTJSKLjnDERCMshhANUoDh4vMuB7sZx4TM6JVhCrBeeNJ
aVldegA6sfsQbc7Qb/SXqjdwcDhW5dJihrBtEPdefFrweY4BKK/Wn84UFKDu2EAs
Uon3JCJ9j9VsJH22T3xJ0LBv0lzVQPPrGCrsBeYnjOxkIbvtreGcaUiEE1m4AzkY
a4iCQ0F4KP08/vr8OwzY+7nEhB0eu3sw1tcxhkcg7f1LcIfQTKqF6UvZige3rXiH
nYysSv9B8SH6HUGogNRNEMTNQ2mF8vIoftSQlyrSlYS6ZySZgNVFhST/UAurNoF+
Tg4veYjOlupd1ak16so8+0SSTW3pnfKsgMy7CxE8F4vvVlydLkXmqVvs3QPhfFpS
5f8il3G8ZAF7Cq5XhJ5KP4siffICRhl1cHrHWaXmOODo8kjAw1JrMlYtN94TrIwU
Tu4dzIjC0xHkisBVDND/ml9uViCOUZV0AjIPkFwUmAyoGCcMnHIL9EqTME2faiBi
HPZFPLz34mdjWZZgb8MLe2zHJ+GjchJfE+hf1X6Wawz9q+X9J/CotyWNsaKB13Je
KoWsCgAGqoOHUWn8RoISdACfIEa0xGbcSHt9vo2Wrk5F2l3DVvzc5ytQk5qDUbZM
oZ7C8OZW1m+qrh4xokmUlx3SYwC3NlhgcJaIMNw0twmnG0XIL8BtpuhsexAsD2Kk
0znAdfmcf2qpqKJAzRCc8v1xu9NPRpgVZ+zmu7GGhS6cxh/aipkfVOappBC1hRqU
lYx9CmRwE0IZuDdJvNvUfMn4whQ5Z1i+VrQj5ERY87qwF2XMNPJBKUVHF8G0z+2H
hsBHQRV+gV4rumQkw8pBPBaCfHATtNfh0W4DkaFoLNr+fqngagjx9ndv4a5iVI+6
5e/nN5mXy2X1gnQMhyO11vO1pHCF3Vkf60oUbB4C8gGyBiNF2vNcxq+YGN2fwcST
TZ+98Zj6ahn2z+FMWbFUTo4arCWMTVmz/mdy9+RJ0y9BEy3kjym2IQDVcoNM2xiz
iejtTPvG0Aqn3+7DrjKlqGRFdfywKM6Pai3BlruHEjKv0Bts4nsZ4ZYRkYoxjmFP
3o1OVYELskxugMXosbFu2p8I+d5uScblBX+AGE276S/WWjdEoAqMrt3bK9iSrGQb
QNvUxmWsnZ8Cjy1zzmuffxmmk79V6WIb1xfeqHNUu97TNgQFi4gIi9oSpvjjanYI
u4I7KVDTETuZQXJpKZo83xFMXaq3gOhOea1cwFbCr1oAydt64+2NvosZCskr+6Kz
G/7xfwk84Sta8csw5WI/EDXK4ZL6xnv7vuu26OzFdzozN/wSPxNxxU1DLeuhZqtm
FeLm5pqMiYLlC0Ro++yY1jo6+38pnR+oc9emk03woPpKpLmTyAqWO86nroSI8pX6
lzO+5O1kc4RHy4bwZpJD8rJ8C8lptC9dI9l8Xn0npsbjh1KbaDfH26wtr7vW+FSO
5GuWRd5hHEMk0VPDgH3cTHxWSNufGR7jaN7+bbCwVZBZwIkIW99mc7t/WddwzYgz
CFzmsespgG6LX7hyzx1GCvSdMJF1gyrB2YXQQVKSvOk7gCpctJ/rF+kmRDd7mJJU
Kut2vosNWzWmALiBlrYiZUpxu7v+ANAI4C929ftmysBy791LE2BHp9goljzuY/fv
NiZR3kfOdE7dAOw6zKOpwsvrfmKt8q8MjaFl5ava16NBqhl8fZmQZN/fkpzHOLO3
lDSEulNWwCz7mO1K1c8FbuEKhg1xDns3heJIQbadN0pYgCt3PSaIv850AeGwL7in
Zi7RkP4q22WusLA7cWCXUNb2pqQVsvhvx9G4OcBcb385PTzPDJ1MXMIXTA03S5GP
Xu6kYr4o11XxQpDPFVVBes4UHkozOiTdeuKaHmbVY0XAw6jPCLvL28pgr4su5w/8
XIxHyprxYGS09OBwk8UZOcBWoeG0wU+cQ0kMv3vI7KX7XEhEnNoFFVkqBMLtnsFA
URbi14EXQ9XNsUh+QF8PUD1J1zwz3aQ19jk5t+sVuKCPU1mO3AB/gYSM0fFDTZ3/
5CYKWQ3QTrTklCw4qeTlwQkQ8Ds1ZZTSAa7Exeu09weEbpr+fXbuEnJ5fABrfaST
F/2UWCZSNXKyko+4nYZuMb6D35v3RhJ2AMLpXX905zOWG4H1wYcXthFC7+Dw3Yy6
XlZ7JLEKwggq8/xV4qxoF8M917gx60CjLEpS4ijmJhd8+5sYof8jQSZqlhHbhfVv
Mk1tndWPwf9utnzjFc17Qmx4E/wvNReUErLEY/KpL5fkuBviEIUpo12By7+elGx1
Zq0ZkntSZhxiWgzNfePgeYFUnYp1W+/2z/2KmLDi/ZYd4BvN3X72zYnjO1E1RTgV
sNsOJUiPgoTQDLogidliaZXroWY+eRbcr2MbEMit/KzNRFGdlekCm+rZbBJpL7Dw
Ih6yQwKY7zrPryJCR5k0QoHJ1SNiZCdqPdb7vthqmZpy3RXm5N41dgIkztYh3J+l
XIT7dkW9PCO5WNsrkCZS2cJJWmCGC/IQ4Wj4vaEYureZQlibpQC/IPHQZUUGp6j9
JmcR9kNqeOAVTqbMfY5u9uEiSRjpzyHvOI/xM2tsM3DPiCfoBg3NopSnP8qBoYvq
MyrABAJ6gsPOAMgIEd6X8xROaU/MdNDWL6KnQ/vTA4UJ2OuvDsVspvSTCPeT6wDw
Q+LFMgG9fH4WODN5Jx5dO33/fczv/DaKPzkya4wY6juKLm7dO/+5KGMiOl9zpCBT
TvAyMTphDvXG2IwK/ZVlf1pPrOC3vns4irkFflMbatsSMqfXW7Xgl7x5ES+8ACeb
4PWaTpVVP5Nquo91Vnc0IGbYq6yKEi0iXpVCMS796MKYDYLBrzgdzAZ8rZygG58p
1JE5tjmOLoYBRwzr0t45oY3S32MMUSCkE7jTewQaIe4m13kzBnVdSUol9SfjdDKc
BMlv6EeNfXXEFKe9oleWLqfoBG57SOaC+l0RRKIWNaSSGoqtbvoat+ShcxW9uKk8
MoA+3dDePaJzzVMDLu7auS8x057sssDobEwurCKuFY5rqgXjZSY7MOhgcAtcRHFH
Qav/pnrCAMyuMMa4ZyhB3XnL8Vkzw3JTWDngexRu5ASAeEm5NRASPNZTaMyg+tvD
W1BWKKGUmFNOqDfMiA8PpyP6u/nwuhxQz8hepf0AEFmesYV1xHKIm1yLgm7k55r1
mguJ6EdjAxbq66r/WIHVoJHhFNOHExpaCrEVw4d2hx6zu0X7v1g1fUNd7VN+G8uq
Gk/gyGpRUqxJAAtzTc3cBU/9xqTWQNZ7KNbOaPLvVlItQv9PLWp90jKjd2dCqX2p
hGLOJHFiizp8ReSoqwEdWLT3Eby8uVd+KuReUzBD0BLd9VWr879ws3T6WTrd77GI
aSOP3lJHgv05+iFyzq0lU9dRDDaiBfg2Mul9jXpsPWZKostXRtgbeGxdWbRfrv9E
7j9Rwg00im+1QD06ys1Q7SmNirkbnkK76v2r8CzjCbaj/v0HEs5Bv4/vLcEi9GZo
tVbnff2F6whXSPzwNGvOcBp1QGVAO5/3/R5W0jCAvevafr1YBm21L4wyImtPyR5M
yAFN9Js9w28n8CL6hJlNJ2rke4dHvlEZwG7b/PlLaseddPLouATKJUmVI5ZlAbNe
9xZnh+YetWw/jTGr7hvKnSRYraytJIPImkoW8+kIHSa2cJdNA9Xrd6u9SUM9+D37
Ig1RnpHvynri3aQO2LFgjryyBD2i0oUbnNtyr31Pvr6CLKq72PxdeXrwQSLruqIL
miQhR7qZJ7NXa35xkNwutw==
`protect END_PROTECTED
