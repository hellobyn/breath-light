`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NDk4y1QIR2vclX530bOaofTnE77h8k1nuuqRXeMRSlH782raU7oSICZhHPqSfiq
NoFYQ154uHi9G02yCnHaCnGEogMl4JG+DVKVv3Wri7UqHj0xsuIfPYPrlILDg38n
D+st3UjcXKBisGNLooBVBlXu9bE5wzML6hCLylRUBx24EqJszbe4xSfFFeE8Fygx
vcUqYhOHBCjJ8eJ5qx4YjvP2BX6jTXa8TXNmlHTg/UiG6jhy5HouVRO/+DfC/44y
b2QidVzamcZcqVDGUBgK3rmqfEQa3t5jiNCXXLXY1EEXT40FUBQL8u2F+JEjwuEX
ihlB6RBrfDVai8wyX2ZuOpUOVsnNGrKmBbDKuJA0/CwRkzYPutFniNsj6rzC3xL8
A2XkpVNmiOedrKWyd/2GOPyLGOxF4o16USHpR7O2B7M29lS6P/7nrrV0oH6ps3ml
Se8pDycp/QZNeRe8265aZzLL2tCF4j0h8J5/M+a0ifJdv4aZBWMXU2kz3cXD0MC1
N6JsHvtBc9Q6ZkqPgXSbbBsButJFmFhYiHrLdlXxcTApDBvRGa1mpDdbrJvXmiMW
/zRmjrm9FXyBrlSXFOEggMZl1mIJUQ083MDK/U79h9SlQh6r9crWTFdvVWVJzPF7
v9qJwuUxIklnhxmwKF02pBtJkLAr8+4AmG6Tb9/cYOcvr2WHUVSUK47PYFxVxUoI
AVQ+xK+ezvrrXfyP8PJRKHi/uUcr58uHgFtFnStox1aEKKVKtv9XschX7n3jOAhu
+YTkWou3FhAH02wdFY/fo6GYsyfJzafkrU6/eczv0h0ybYFGB9wAiaVZBkk/ivqP
VTBQmlR4ERFRBwVzjNdCdPncs0FTuBI9lNevRUCrvz8BrkNrT5GgpKLFfXI2gvg1
79I045na82BeIYgVyWhMVf4dzMPQboTSY0X/+sh6WUO5AxGRRgD2S/k9H4QtAIqy
LM4c2QQaXHEhDT7wEllRXc5lOYmKrbIq4WGKO5DUvGpkN10Ux5Z7yd24KseQcNHl
Mn1Suf5WjOTtoed6jEFNYylCICoTMHLt9hAmai5azO7oJQtWByqggMB9M4Ah67m+
TcNB+49PjKIKqAI7oQ4BJLhcFr1NXEih7i0c3csv8IEznPw2HkVeXMcZKr1EMG/e
vqNFw20ouP4VwoOtMZd79eZ5u1vDmncswVLbFMoCKl7OTJLowGyTLmb/13Bjkwc4
RBmtKuvynpsRpBsI+yGY88UT99pzRL72B73s6EmgCF4X0FD1kDZF+PqmMWNK7XpW
O8jh2QQZrMS3X7XOx+902k2FEZCNN4t4vRGgOxZiOdpLdx6QcjvAOVWQKPKEaWpy
GUD/4+q6dmaNXyqADTodZdD4wyT8P1JHC6XwGRynZakUuM+TEKVG7VIPu33EU9lL
rkT6kQeHI5kZgbTu+Q4BNgrRhNw7JWZ7TxTZQZFuzQafmOeoRUnHDCRw5FwfCuLT
`protect END_PROTECTED
