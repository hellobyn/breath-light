`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjlIdawBNGRNNSVd0qHa+NhY5pgcqhlUKfDAqVRaYvJ6Np3Dd39rBgOS9hbT0cOw
t3npS1VjDHSTtzH+rz1mEMYQ8DKoXcf9z6jgVrzSzf38kIx9wEzpjWDKODNYHm0E
DYS6Fy/pssKIikFxo/PXWm03V0WCwJK+7rYwSA9wIqBQXYevT/5vtMON3NbKV0/x
bObVsBGHPO/DDIVQIFQTOEvsd9lxNp/bjL4BVLXXku9FJiqGbmqwX33QaqbJtO0t
k+A9ytenSKGxa0JhVesQffTwplKVCZwjBrxIHqbmvHffYwzgtYP/U0FrhjRKHra6
4/s206kAF+4ZUcoASoxdfzovDLEeQmuPzG5X7RTRZXPvypdy6GAvPtTnAI0zWE1N
m5IVwSJru3kZnc5povvz1b6UK6YLwmam+oJL04C/GjknDpBLFdwaS5YALnNMKxtH
DPFUjdKAWXhhTBmsHS9arxblALuDF/WuzhV7uRi4ZEWsFHEQapwvyYH2DMv/4KYb
8D2U3xazWKSJFQu5i4d0NWMxv5Or7VxnqJZLSIzU1W4HbqIXDDKM2CmBOQpSHxEs
m3TCLN1EdOQCyKCo/WCVRm9HOe92tS1xbi0mqQn/5RhwgPpNqsVA1/R3t17zaucu
wcyakn+xMbbqreW9DbBnZyCnu5vM36Sh5hTsH1wGN99L9MkQ9SCeaK3aMDa4Iott
4/tOOLYFP0rMTy1ze0ILAl1az50Dqvonca4QpV1FGv3QScR1AkdgzjUT1wtUpEnB
gX0GOUOJu+S/IcF0NT/wMy7wyWAXqXrkOMGiHZhC2QI9Oqw5j5GKa7uXPX3UVROG
2vfPyl4oK8MrYaBejlH+TUnp0PwlgokCVmILSFndqgYkXOwVkyrkF/Cmyz4yPAkc
qNknIe6G0iHHoVezCgVsm3PWNjvSE3XCas02zrVSWS2A2/UxpAOUt6zBSk0spr7z
uKAJ54CHzCr4xon1izdmMoJKItzPuRIxGyNywxaR88E5VyQWD2sa1zvicQDDhicu
O1dlAGrW2s0sCqg/IzHf/aNSi6PtbxmjuCEf7XtU/bju2jOJxnfYxMgr/1w7i5Va
JhFe78vUrNdtDKrAGg2cPzlyQH9f3J3csqd8c7Hvgiemt5JCmzw1o+yE7ZIARkBH
EXvaYoNFY97jDXp5LE5TqTaeYpqhMgQ8rD/EAYOEavJELLd8prBDgt3nyQWEzUFh
4E9ZYLkmRe/U0qlFLmVosGFta1XnWPrL241LqAIBPL0H8DdRHCQtUEc7kcjzgfFV
T5sr0c4gOXSuuayT8AodQOu7tN/F3B5usyDi+F9ek+haJcJt4VZaj71b3JXG6RFG
Ls5W24JEmvxdnG/2NKfLGXmzI82Opm37oWet9RyNx4SHy5sTA1yxKyI4TJeIC192
Lrr/dxSU95LEd1SrE4l8wmSYT1bOdkS4wv9bNGlZTiQ=
`protect END_PROTECTED
