`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jn29J6y8EeF2Ll3wIcMEzqWRNRiz9EJ2tnwHrevMmCdzHl6v1/Fke1sFVoNXi0tk
QZ1BtvmBv7e3FUHvAG1JFCQMQs5L2Gyezpc307CyNFT/+gLG/DYz7L8gRVXiEhti
LBv4QXdOfz45coApbcVFSOsx1lMQZB7Lha/+M2iO0YhycuPu/DTSIXWwDQqnat9k
WIq0FcDWs6zXNgKJFeknbQRnWK4nIQgLrUvrMR3PJAa05k+SBXQtRjefnCci27kA
rmOMw4kboQFXNpzcguSl5DXDBX28gdkaEiq5A0WvhhRmLn4e/XTZFuUa2ESnC/Js
ECjr8HUZ3Gnm6oLn++X1SPJsgsamj1iCEDRP/mroT0DHlcd6EVusuEx7KzIRN2sj
yozA2iKPuhQtzboxZjjhqVB7RJMenylQbHKfqiHy3LBo3n6k3oSMk72gQRfFo+R6
YbNIHa/bRazBaByfBEoAxyPWcH5orjvuDwTJoaakSj0k0RgFxFCZelZCTOjvBFum
nmOcCyvqi4vdofaai9eLvJ0uKTuyMrEe/4JynlFlwTJG6wt5ymsh5m/lE2nqmASp
nIPHLRMwqIN/6cbgvavZfge6AHR/h8pjApyXeVierO7CqFAiGsDA5qtHRwb/H1ZV
0D4r9WPfifJZuIQTQOi/5n53qR/UD6DP6/dj9Dr86bAiGSZkVVXl2DnZqqgH8yvC
NvgttY88dD+8FL/OHFqkWg/pSq/nBrXG68pLtV9guO96Ape79ZWFctFon5I2Yu3r
+dFUSj0U3oZSavFm/Z1YHh9W9Ftjb8jzCKg5UTdYsek8iLEXNrM1WyorLQqxFayc
1bTmJtoC08nxcbfP+KSYIcb9Y0AyipBHn+zB4/TVMPhAQIVQzPwwx0gQ0zIqOjZA
eaIkDM9NJlqC8PzfI8yr9i4AYP3xD5lFesPY65A2AernF/1gh129VEXZtCo+yhHO
WqtczSbA2I3ShnDVHoHnUR6kqQt54jC6TKGc7bueUdJi8SawRlieBEobD4EeYrvK
OT5Dv+YUQNHYkrlKqrvSbTjCU1QbIhJQuuVE7yStzQU2nlxoLTeCNPFR1frNXjUp
hEwB6Ao2wzT+Hf+WNf2TwUY7/PBxfY9s5G6CLtg2GZc6E7WQTW4GqzUZDWO+vcJt
1aDAIQi24oglpqcx53DzaQJA0HYjky0guXKP0DYXv0D98c/jmJ+yqnxD44aFHGoj
JMxQwWy3AwMf+oaPUUo95e9V4no/AtdbwtlODNV2DLnuklMeYJgjIdfRdNRTMsGK
3XYdfCD0awINyvSVFjeOv86+67Xwq9tLAGxrK9riJUnfizP4642H1IS74lfjAfDt
eCK8prEhMubVQW6dZJqWfFw7hazcAXbNvnzpYrdc6TIcgNJ/7ceqpPfG6p4kHROm
klp4uX8vrPH8vXrhQSR4gdiZ0i64eP7INa57Yo/Lkq1Pfl9nE2YmmJcAK6HYgdWi
oPys34hZHz68iU+IU5jw+FMZM/rZfE3+MaxFJVHtyQa+NeaMPDWY4OIfWVvGVI6P
SczB+FastvmGRMftd+7h1306B8jzqzrf/4/vNLVxBzNvinZefpJGEo6GuyV8BwdE
7w7z15A5nSN8QOZvPxJsonEPZGg1x5bASEEQkTNFICzb8ZfFurv5aYOdZ6S5c8y3
8GQiChO22buK8D9OPmBUCUOl8F7mDvXiHaa7iFWvvXoPiGpfK/ObMdO1bI7+TnmS
azqpsxUrfuzmx04lt8cx0ARnexLcJhShLjewIyaOJ1ii0ifdtzv3QDCOBrojiEBb
suulg1MeIXkznPmRuLVt8SUn0gaf0QQuLGwAzlppzrDyQMNUzS8iZG7tNg7PGSuk
lVZ/JnSnh6pYYoidFCYw3ux2ZVNl4R5sB4C0LWjbKcXWTGfcMTV5XEJ2446zOKmp
k65RHL+s3HCb0t5DsCKQB3r9y5XQJgOMxRSAmqgTyVn+oL7GFKfhjJzcYleREIiH
TArEzjNet8F4IkRzqXVKjw6oSyKd9YlpUv5zl8j+A3TdodRC5ULRZi+NvX0mC/js
aJ/wt9x296D6Sk7xfZ6YvJo9Mxv8BcN3LAmmOSGrSBbyAq1bkyBiDqqYSVw8vCls
wOn1qZyyYv/m0i6irXUO3Hdngr1il2GoghkuEU1wHaaLDn+GZzjxzdYBtAVW35/E
tVp2k/DghJ7fuA/9MMzNkUg3ObYR5im6+DznhBeAKGcFeNmwae248AFJ9HWGfWMB
DwY52E2c5O2ppgr8sy6CI9NDzRBh8oJTfcqVQiE+mQhRcFPFhKM74hp7eBua8HF7
sav696DAhnQ0mTQOopsd18Hqa3IntfbDi1MjPr96UpcGfW2XpWkT2JWJobhndWkG
u4KwAsC4K7FQVJmhpNK1CcuP+ed8+Afb/dqkyXFTX8UORWz2DX4zE8icwBA4BSyA
rkBS9yDDl8JSdXg3m+0sbqO5EowLDBUtq8aFSTmj2hXUnSqwul+RFFBYD1iORjUZ
JXs4SU/rS3thwrw161lMEtsxJSvSERYg8ALQbUrbzd052Vzb0CelKhp29HZm8fkT
oCnNZNxgQ7MbUSGu/mKDz6oPIFnI70F/w9/wNhEw38KEbR6nC0IZwrnadDJjgvkj
iQgMSrnlP5mAkdtR/lmPYFXMWxxRLT6df3KzkvQo+/YZuF+y5dAH72snAitbE3mt
1ZBQHghLCLCaEpE6tp89mLgqO1pJY9hvx25E9bm2s4J9y8qvzZjQvji94i4Py/5m
8hPdP2dyFBTW30Iqm3iy0uhxsbp1BStZfFtTYZlPpSbINCY57+8Lg6bTu8fFu3r1
rSu2iulrhgmf1MXUi8yJx4dM1XeJxhWFsxEZAt6sjm4th7wL8b1r59SIYE+yREHs
KvTpV34a817YQxWSNFnQLwSspy2cLFEHm1rvyw8aowc66Ko7G++LKGWwPPdVFQXd
2P9lEwfR9x8c3flkvGBH4B4X26obu5vzwa3kLOJ4xtvUsGABN5UU9jsP+ExcjsWN
Kq1rIo0QvlDzQK7NJ33VFADuHIbg9mk9B077zPb6Ou9/BC025jH/T2lSfCtVe+mX
YxZ3ywMFKY9X02YvPI4ay8JQp2JzySsUmL9USO/Va6ZaQInrjdz1J0IQaDzf5+i8
J+W79Z7cxUmcPP8UCcmoRZm9ymc8MzvVMNYDOEWLZKBOzCcFX//YkJRB5HW8SbWZ
IqiESf0KXy+clTByKHgbTTyUoHk5Tu5hWmfw/qpeWutObRs9ISmwCBXgBMfky5TW
/3F1VFVQq0fJgtMoVIdMPEizAizIWZ7yDWp8p+yu3MOPZAXAfL6jie+3CCY0cEvw
HQr5iHYyNgkqSQRccI/QPAcanCqBDDTDfLhppAiJjSpSDqz8Cz9YrdFs17pR5UMV
79uoCevYO4L8N75X6i6nHhv/MMXBEhgEghBgzgLyBBGsxQROoWnVcnOLVIBmpoJ+
2XaL/9wtWs9aVKvxzSZycstG+AlvTbzSwzhEFOxgZJSNv4n42UWckm33ZLUv7znO
qg5HcJedDKa9iMG4+dPr0201PzFoTFxk5GOVk5kme07YeFUpm9BaCB1E7Q5T6F1Z
swCkNSGHWVrcHEntvi7p5dW60pDtJFXxZAKVIieJjj3EyDxN9GvyZVTFH9kf3M3q
nkSFjizyF54Ty6lcBb3hv7RV39kbhFlwBEj9eBs9fXfXgjdiZMdLALtPdwAy7rpM
IAWia2R9dCUbs27hmm3iT/yX9JjAa0KUr03IYgfFOUr8jX0kgvHnJtTv6opglCL6
dHaUAzpNbTXPWUaG1BDEnXISd1H6Txp1XOvxQ4SzWJAbzJ68YDk6xUQH5ynHxwDH
eJLY99NaAl7lQmKy6xZnd0hNGpr1PspKx53dMcJXwSzDZ2iHgmV/3Pjtx/REUvfS
K2om/RSmxIpqVekCAZkk8R115OaedkTUmUowcupAjJye9ZOSuw2+mPndXLXy0uF7
t9D+GnauRcDL9UshViQS+BsPn1sntbMcRnVPCIWZXYKLgmAOO1B7q6I7h+RqxONe
3/aWQneijNR21tCI0jMwAysp24PmeOimnKRAhGizXQGDa9wEGafkjXJ5kwRjGNFN
bJPCYVwk+qhFYVoCFafQ7Hy3EyPX/HRlKs6JmtosKgZncVGM090POEukBHI+FtDY
w8KMDHH2A0GZDV/iEvZL81cWtTt7ePn17rTz39YaqQZU1z879+xgKkwacyqY1Fse
5dSPmq5s2vKSkcrcq3duztjeRBEpYyLuXelCqa6eNPSWcEtZwJ1XE2IkLWYIRYjF
rqRTx21t0HaoPcsggQuyYpV9llnAQZme9k52St9pvF+Dct/dtVi50ofLBXOJVGNd
zdZ8NMf5fnMQp1AWgwYIf+0mNRvVK4MjIGIsJ/uXKJhEG6IFNNdTVwEA1KvMwc0f
4ZZ1qSxkZjtT8/tioE84oPL/2HdlvTesENdClpreuM7X8Bz90TffslFTpuZblCIa
LLFYAJ8tjfanF4hLcXuA5i+RLE4KRzdnY5Xt7oZsI1aIRYkPhoOajBL9EMkC2E8L
OZk3p+GBUuC+U81+FHNssh5GGh47vlwZCFProhh0FjXVpXwTDGnVmBBMCl9sjLmz
JaxhZBxloUjRcZBx22y29xJYNjI7KtPuoS0zU87KiEYS8yBfuRhy4xmy9kYCAgd+
tbdAj1Y/P46I1whl33+FasY9QyKIOfByyEOAKERMWIVbAG5skBK5O6g/lTHlZbzR
4UFX4ZGEYGF/JYqwBt89JKuuJHmMoXrHSyiIEmb/G2VR/8E9E2M1fZJu+J1Ziglv
Dm6t1fjlD93df1AUt2ObWBgk95jb0y+FIGiTZgGTXLVmGAptsa4x192bjkdjqOHD
KXw5Mf5NOVbCA/qWZkgFFW+zIp80VaU9oklMntqS6tLCAa7gWexe1vrBFtuU45Nx
Njb5XPLasqaqIZhRTIy2p6y8ZHlit2oku41Tgk5QAUMpmCfEqUws2zn/aKP6fhfQ
CjXsujzioiI9Znl+v0zC3Romdq3UXrOTJQfuO4j7QKF46sQAab+jQOP+G/0f+505
YzFXiWhbufahnd9PEliPPlJFphmD35WRjqzgeEAdiUfngdd3dRs/IfqTyZO8RevB
F3xNOezStiNzMNzFWPmyXNuDqpY2BC+H6msd/cSJUvzCx4Kk7Aa03vTpb67SPTRG
XE2oCqTcUp1d+4u55v2K8+cY6DS5Z2pNVkhHB4WhlRsqxbUTN+EZpv9t7eGWTCJZ
G9c/SVor7ibFbucVWSE+2kX3PWB/vZCPqzNP1K2TC3eoC6OhPMXEvbUxinZKUl/j
GbmnX38IXHOlX3aLtkwR+RKj/NaCRcqUZ0PHNAEBpTwj7rwVdoB2TS/aZ0jOvilN
5do/XggDrYkxHtQnEocv/VdpkhPtSze8B4TudlMn1uxoKMln6xqdaGWKYLJFOQWA
ajCPGU2MldyZMYK16Xu6q7SA00H0WmF3n8AygPy1mEqfC4eH42xGBAjVwz2Khyqc
cXgr7CQ8e1me8UXjX+O4PCJ47TyeYMTWogwtgYeHH0tGuhU0Cizw7/6lEf/yyfoG
KLzHetpCr9Wc9EuP6jQJwDnw0j/Qf2ptcfzu8GCVoNnc3df9GUYBy2YxRPtM0Ido
6dwwCWtWuAbnSMufQIHRTmTDE8KYBzQuK8mOt3asCyQPN8xnTkQAb/iQ9cICTYya
t7/Hw4lXyqD/U4OyIk0TJ0oeVHDm9ooDUoNiNbuhOdazygOP/gpTrds7YeLPpThw
KkH3vAZtqK3jvSJ3JdT7YTMCEJA+aD2YfUFQkryRIpsjmZf31tilf1bEAxHurDNa
CQtF33jr18yNOeH7c5AkRrRj7Pw88jLSsz29MYoeNe5kXYT9qDqrX4qNN/j/HkF6
B5CRE60w1fplZgszNKF+T8dOpEQLIBcFDPEhBOaoHrJqkq2to39MBoQ6W0CgxyCd
20KmddlILsqRboGJMnWKQCph+AgR1RNVptg25wyChnqS2WUC2OM661xmPGVimCcM
TQGhb+DFHMB4pnyQmmpxj8MPgRQtur/bIwtV41RPGptJ6kkjuyTLZpwNnUu5n8bV
GC9+6w7pB071t6y7PR2ofSkM7OfoChR0ogXjf0L1CETSsgbMpAQASRbL3ftjyBKM
AgP4U008bDXYz2yBTPZYnn6UBFPUHm6OmkD9W1kvRQXThCB6yFOmok1W0d/VkrhR
yAAPRVwl7X33uc8kstibvAW4qL1pLeAIvpLCsg3OP3XRGDoV8N+CZj9z0sCthMAr
pb+s3vdCgkHr+QXgu1EqnstZjZwtae8wcUpSdM1hhshMy/vDa8gP0vBpi8Sl92sV
AGrUjlZSxrzi+h7tW/j868s6Ga0Gez5fyh9DBwJLvgpdImTv1WNiesO6mChnOrGl
DEna+byCq10S5uZXaAwPy6zQaaVZfxD527ajGRxbljXVXx8oDbAlPkIFdVTnzsQq
/7oIxIT202TK2mp4AigIe6MWBdYT0QvG7en2Onr3d0KkYsRk3GjwpkmLsg/jvnAx
vdLd68Xu+QaClvUDLl4sCb8HiB/vVHK7wTF0jD/5MJSUoFyQkdeYSl68KDbVM5+q
YGvqoF0tNZz24FhgINSrfg0RCHUdFND5e8PTbrIqHX28yrP0zck2tuxYD1M+qyan
iPOe7lmnuX9u/A2JsUOHu1Pkce9TAZ+KExMikVuI6LBq4LPNO5UH6bJf29LWo7IE
d2hvjeEeOpgRmTLqF5svht/JuKnOGD0LcKjbVE0EqCGvlbGwwvSo/XU3yw3H8ltW
kWSeNWzrl3Xo8v8GhbEiP3dCSt/Ce6jKQRzfH57GRzGvr3BIaRtMUW1qtmNhAxFy
xaKsNSqzqrKI1VSvQTRm26YecOQqDR/lYg5QcqNjNTSh8Uyw4E7UC7RDwfdycD2W
OMIfVgJdhXUE/mr+XtI4Kc9xRrJj6KTdL+foD67GHr7X0ZinSOhGliXbkn6a/3Pr
AEDq3NxuKvSYT3T0xel33jnkBawnq+UZS4zy/xX+n84iyDpqFdrWIrH+x3WiqfmO
vo997rHNuuktOGRCpCT4rfiAq0r+iyeP5gtvMDx/dRjaTi2JKndTVM7lL+AgTPgy
a8KI6FlbwRLD2/86ELZPt/uUsn/yul3MDFMX/TkneGgJ7XiFoBPDz1MouyG2rLKY
48fB1A9i1NHHzwu4QpaAShg5DppHMbDnKL94mNKB3XlcI7HyE5VuTBpA4G4A589L
2qeuDzBiz74E/mEi1Y+riS4z/cr4Rn5vdBO2ZPfwF3g+X6wQJZzhjTPGcjnfRp/t
ke+WFI47Xq32BJC42Jx3FDh/lAs3lOtN9iN0kbLM7HbbBYppHvlCYFCdPTvHe/pw
KYnWaiZq++UsO2nEzLBg6DCnS3HG1WBFvhXPHk5sok3vZaWrdqbmMs5wr2TPFMmP
HZU9H78MucrX3i5VCprYbFX/UhKVPYku26tmNYsh60x0ljH2K4zNQWZYzfU+USR8
6UirGFb/4cQBF2mXQ5+f5IYfsdinTs5tm9IwCXZ/xHaRznWM248I5r+bPpw2DKXh
YjYFYyhA/CT1a1Fu57OXVsH+floZPVxKgsM6A84+TArLg9PB4kTTjYKRggwGpmvi
3OH82FK+D30U8xUTZv7BHqXnocLSrtPhbtUMrk0AUfE0BBH4xfi8lGngKP9VU8Sb
8ooAEA/qs6vb0xQz7crg9R58NriGa3yS9kuZ46DKbFqDFeUQ1CUbcleXMr21ri/t
w6Sd1jGXJ8yNmr6M0FGkuagIbOwQdMIs19Sud2QsLdehXjCS+LracNP2z/QVKU2+
bDZ9ETgMjN9EiORekd9oMbXYogourdMGttNCkz2JW7lelPJUH/XJpjKkuUa8AxaK
F6rVqWx14eXlD9qiUa0mJ71AbtDYUcV6KczWbqg9Lv0MGbDxcIFZBMb10BO41Xfp
huTzHhOVcl4uzYcRzcnAejxJS2SxOJ77PrClG3mh//+p8sUmEtlttF6bhKNun4Us
JF8+d3HnlqnFDVPjVpVLrusuuWHhaucD4e6EoL0SyADwhZk8S+CzRZlEcUOZEX6w
tYhmJsVMqFmf58pP9Ns3ktpzVSKkIkPNAOIdhCQ2I2TjmNq/aGFo+Cil4R8mKaaR
MWa75QHINZGtBeRLF+Da/ICrPHaw7bsx4+ZJ3W5utSKsq+llxu309wbN4k0ctsG7
Moi1phShpVw/WeMnK8cCW85HaGaE1CC7fTKqdDD9vjDvMIm5Dh1k6B75SRKibY54
kc+OOtif1YBN8Hza5fUrUiEiTZFE2lwqp1wn5k+AEXlOCGTLsyyh3MQBjVxtg5xB
N76q+GzjHGmYPzwzqyaqkrtP06Mb5mEdD26D4rWuBGo/Aez2inWfj6u6gIfZeLyg
vbsAneRcqxuRa7bvckene+kbfp7ezMFVd2KSs73nlz8cn0pJ1GQH1v8vkhFg+ES0
Vg9AdJRdiNRuyMuTr+/IEXbmTMFhpoV96fXO2ARZtI6M1HQm+Gx9hK3yuLzd3gLe
dpQc6tpEUR0GaggAUIuZcIK8VeuyAHezajN4ffTitER4Lh8kSrUyhhjoAe3xYn5b
vnhtj2Hui5mOs5O06LwhBUWffi616kx9yG2GK1dH4DtQcNMIs4U9neFyn0SZeAja
8GArTvsxqOHbj1FkjoZMXjR88WXYfnid8ItdT3FXtqDJVYj7vrfch9qhk+ECmevG
1gSrvXplWqXS/7txVFKgSbWVQV2ix6yCzoV87iBjzXUEEe5dqu66S2ESdKq7cpL7
5wx/spTKGcaQFQm6kMXjLrlG+pl8nO8q09oSdVgGt2Hfc1p5IZqUMsetscbeD+sE
apcV5+TF9eKOPfSO8Ty18pxSI5CBoljHJ4Ivzjx8y6FWhF8G5lpdRMmHn63mkyNL
TsOohBOTtRXrmh3SSXqbZQy1R/gexo4+BrQPCshmahz4/JbTfR+l1/ehz3luTpsG
qMvzwJ1Hz8RI7rHE/Wl4x4MJZMzDJk7tPF2xYy5sZS8TEFcwtXZhMC8lZHsh8KDC
o1pS06B7EsiMirK2cnJZ17G3Juv82vZ95s6JoI8FvAgPzSCOdbqo1gjHWdlRN2mm
1krrh2voSi63U2IGSYa1wBCEUXclP7kcojZFNU052YdurHTxXB6fyLULYsw/Lqfu
BKaibIFGEHPmFlSwcYLIBVekZbURgLmT2C97d7z6E0z/iu7X0VR6J1mRsINGJ7em
tM769E58rE1wp5Edxqw6pY1VUvyT0zzSsYUauidkk7Aui6bBwwJAA8thWakeKVr4
m6KqA+GrJIzMTYDZZtfHtLzCDrcE9284eHc1Ml//2H6IKZvxXzkBFLxOJb+uVdfR
4C7+etsUtsou6O1HCb6iRA3cNNWDoaVcNzt+enx0SKjoo58JhFEWFOvrmPbPil4B
qovo4zJfFz94AA1DNRQWGBqtbUjt6MK0VRfFVQGxvudmozluioahYk6dJU6kudCG
MgI1Anjyx8xg7CRtC6VDstTjE6iilIM/HEHBn/ex84WzRQisl4k8FIB/pj/3+iOI
RUe18pFWPQGdYJ4yZki5XykbKiDXuKgiy12KqJJGYvDKlm5XtuzKDJToRxXElA4r
/CIJRbDXK3qYD1BoM8ZtyPuM55u+mioQZ6DIhD3qrdzllp4q8siGnApusa0AqV7b
JR4JKBTibktMbEDn6sUP26fBYv3X/r9+/QWi3uS1dnsPlKD5Tnudadj5NhfyztMB
I5T04CBJJVYaGTZ5Hkz6i0p267IhBXQNV8znizq/L2SK/aRlOuF8QZnkQKdunj0P
zM+ux0EGKwgs5YGCUT83WqWg7hUmVG5AwuoTBo347puZZ83Ev03smQhdIrQFsK5/
wltAGZNp4d1yQuS/C5NmZ5t9bF3cpL51PkYFHRSk/82xWpOK4oq56vcMgevhIvSu
tib1S5Qat/06QekLpd9Bkfx+/DFqt5Sl3KPwhDkUcVDA+wEHhvfVcHk2flcN2M9V
fyikozeoG7jnw/0dVuwIuxHvVjhA71MPxvjpZcy/hllQBhTdWosSQXT4fypAWi2a
v1MJRXjXoMlmJ7ekfgZby1jtWolLzSEsLcD7tGtnvQMdKtxZq69dCpuhC6VUawhf
4NTVx3BDGNEiy3KPUxO94SgtMsjnSMyrer7NbfnjUoN86Ld2GeC7pc0E3RXe+6V6
Qj7iE2DcLgR9EwTgbxYPFOBa1CAOAuAfRdX/DrtqjckyZDXFh/oDiPOdeQ3mK7oz
Ai6TTSmoaIigIGcApU4cITt/ha24N6hz2cwBkQM3f2Oq6JENqvkZKVR+MvRtlrtj
sZhow/IdFVsVV+20wxOtcXXZs/CtXDdeSDdCdt4V7fOenfSygR1y0wJWDLojvAwI
V97cXhbqB1OQeWLWVXfAAxx8SyiZY1K172L/E4FTpUuNdcYO1mjtsJIWrz4yfTMS
PsZj1G9CDCy6mpjq4MqLzl1hhGL7hrh8RRqbekl8l/tqlqg45u6VS8BIREqhtP/K
Fi1fCucXZhOydMD9Oi8fd3kG4IMZrGVfoUYH5MPy6COyV5mJ2GGSY783Gm+OWGbn
AKftIr11k406sgsdG7GA6ducShyAsPQlK+KOGAJqD0XIojTGJmLg+m8Znfo10HHw
Svfwxn12OpQCukVrZCQP7ORGKZcVRbNnA69e5XU3l/NVLI2aMaRRAOATn+a99pzk
mzXZJ9Ms06O+eYP3KgT1kD4rS/O19cXz6sAsikV074RvP/e7Iu2UHTnGY59AFk42
3pEfEUWNwMsRYy0DIp3fQyaz4Q0+FEpL21iQH0IzOTfgaZgZiLqtp7jxH8ihutlg
XnbrCRc74Z1/kXg/4XVRsvf0XDsO95PLRXRTIgpyKJcu+WsMRZBKwlB5OVQrWi7c
FkdmDyWRDSpmCXy/pGamih19Be2eMSMuiVP004pfk90c0IQ2Uj8rAHC+Iel+NaVG
TEEK9QW/LulIHBx/QL70I26WdLVMaLE24xu5dUGrgOuQSDPGNa0aNp0H6A2E17i1
hhb19b8uwBK2P5TDJnaBpz6gSvGUT8isY8sZyQK3PPkeube6LU3mEA3l6qxq+p6Z
llVsOdYB3OF35ru3S5ODQSwuhvSbmJtJekb9kjJHOoGXtrm4MyeZrCVuO+JR1K0B
2cHUciKG0WHqiOhu2xEE7kWOTsnUPgeXCXIvlpVLC0SnEpQU4tWFosVqszZgz5hz
9uaChC5ZC8GM9y5oQnJmGcbI/WZYjuaG0XCCJLOcXIDANhflVeGnx2EHYtVTJIeS
OzAoybSkLaT3+R8fUDziaqX6eqfbsjlP0zuNnJa/M4hUik/pd23A2q5tIjphcgte
iGZOyoXgK8442mffWyioPUf/j8/hE38++wE378UF/qGgO65Ren76n7OaaAv+lL46
NCEH+D7hCwtUrqWXLtOadmKXs7A2mggGY7BzXfKG4RnGK4tPbVHNdlHJRBnf/qF2
rvUMlITCeUcA06cUWyK3JIcdMBDFVoGybvCcZllAyZH8bOZxt4EWNiwCh6O00nrK
RKO+YGuw41AwaVmbxlGs7XJkBJh47dS27W2ojYcKqz7AwLJGqce00G4QgT4y51+E
CUeogSo7NIWnUbPEf1SxouAxniW4cSM2sVTATY5fn9j8lZ56ZDxH3/E4Assm74WX
xSqnVQXjCu6SyuBb6APfEggvcWhgSMg8IVUHNgBxZfSHe0ldVXPyFn3/Zvip5U0b
3fsBh3nE5UXESzrHgAd5CI04FvEZ7I/Pjq6ykAWHN8kcgzqQJGQVz1wSMI4Dg6Ow
7LTT//RZfsthMHqUV030WNZpG9HXkNYBpTMludrmVhjZAckmBRWsbqpcmO5ZbAek
dpMVhoUlDcpYHdc/aczRdwFTGgtMhCXP3t6MdyLv0KemKfwz8qLqdPxD+xiVCcU/
KWpU80N9gA+jFdpmsbedMt0O4QN6L2Z6fFdpas6jJYtTHOdTwoLQD/fduF2831Dw
0kEjvdRqq6fHc3QSkgeALhk8ouOGa3Bk+CydI3aqVLeUmPyM5KYv2DXXRIHZrD/Z
0UMrSCFm9f4mPPJ9s1WYhnQvI6DfFMjU12g3hiMep6F1xJrksPpWnEPedioHC1Bi
FPdm2mbkj/QaWCsbmjapruzXTHS+7YWNaEZaiXI0lBS2kute6In+zNJOryxGcvhB
OsOOC5SDH7Riys2sVVtj6nu8box1fRRK8GIUFFhKbj5Sk/8AhC2LoHgnnp828PFw
sbdLO4ezwgDSsjc39nDBMCeSZkKZjhFTaqQnraLeU97XHBrozkU1IV8jkT7HDvfB
esM4hjXmgxA/pntBA383GQi7gXCo1M1Nx3i+fRrUt4yv6JaZ4tPdISS1xx5h2Eig
WZDYFf27neH9LBfo9Bd0iyvrVzKnxYVISpttO3Wk61gICNB/IGNrtzpABwr/Evl1
PYeTxP1kefQNSzNy6T/6wQsi4uiY3Velf2NZdbPwHvZW84rD2/vvhANtGaAtAxjD
INmaYS8ER9F6bhq9eHSvP9cdcxXugmC/J71shzqctcwSEb60FPDgF0uTdJOLw7M5
1r0SMVKS8M02QCesR7pUKDNDgw1C9moYBeXEBOXsfp4fTlMTsNbiw7K3Rufkf16f
6hbhYiuUVWkDDnhtuUVQkpnWcEzlFSaTXKQ4WSdRudfbURrNJMdNJQU5EeFrgYQ3
Lex5TN6rOZRqkPgyhHzxSURcmdBzIxiJMcq06MkzFgk5dbdanWJWgDgU8+H/O6xe
u7HjBNb+tRTrxk3VCGqc7YkZG3JIZJaEgoU0uMt0+Ogprzx6DHZ1XlHBP1FOWhXy
eTLjoTsQKkiyxYU8ND8wlLtTtaGiuBngt3Yp6we8f7aBUsHgAvlTPzgGyduxM7cf
ugjcfFwIeGzBem3jD2gpvfBtSnuxvOoshvSl/AAVyP9E7PtZRc2JqTS64wx1r4Lq
K39YOs17pRhKpZswkc09Xv4z637BPQB4sUZmgB+GOsMyme9+gfglE7D4rcDm0PDS
Fqy8rxFkmuLCBwC08X/JTUcotCFnhqCr06mOBC5uAs6BWcoXgGFTkFb/jEzwXhTi
AmA4G8ioykETPJYrjCESiGCeeRY4gqd5WlIPVZ2NB8G/1jdda6j97Gy/Tsg/Y4CB
h1VT/aO863appWHwwu1BS2gvqD+rplaG3q/tuwCkvRErBGDOJaiRaVsDHEndBBJP
kQXsledfS7ggvEny7nOY+NDQkUNUFdOfz7yypYolSip44h+rP/rhOkOyQ+vnJ+LQ
3gyInvRRRBjH3zDY6C1YdK8alpo4h/VjYZ2+oAunqkURD7llhBJ7337yacpc9W0/
vWd2GGXm04lgn61zA6/LXhZZxq4V2WnjMORhLH0DLwiDFXDSgHjw2kFta6burtMV
U7Mks0mLm7K+FG41hZcMMujfv9lOBBQjaY2T2lppdKFAenyzKx7YXTlpjzVGX9Sq
u2L0drb3v9y8Zntti3BpvhNkZ186xrW9zy948S/q+uyboB87GTVA6nUOP61FoBXG
U6C1RWuxR+cgy7HNfvYLIqV0XDJ1C6QjxbMiI32K3rGv0UL3306JmtLblZls0Zvb
X+blvKaut8tdeYEg+ldhtwqBnzTBU4u2x4DmKptlt+NKkZj2ESIUKDyc8+vL1axp
6+Ma3uw8Lgybk5i8gt+zDzvcxDSSlCSd9emZYGyKvmC77OXqSTlQpMEROdc41072
ORP/wNB0UfuKPQYdY7K8SrqxKNqhoKp5lZvyRkDDCVR7Cf4okDLIeWuEMQ3Wulev
Mn0eWsd9rqyq5GzHh/HplbSnaHFvdION/tvlvYfZcYZ5AT9LjuUpyZeP83Q+0Qut
scbVKQ6t+V1mHISirPL2P97Z7SBUGn4bUqg1p02OWJe0DkAEciFlquqUE8cFJUpn
gaEAAKKJgu2sCjyFCZAOTRuvMJ1IXbLWRGYFFu13HnQQ34Nhq0zE2+CCkKXw7XV+
2LLTpsf/+uWmGdJ2/L+I0rqfToF6703qOMR2goGq3DZRYkFmw9XP+i695FDFYxzk
3mdZE5uka8evDHkLw4JmtdwnmnLEevnzLs7fUUox8+aEZ7oftiYp/stWXPPlZzNU
a5RHc44ZPZxaM365vIPVqZINd2MQUmiAa1dxpVLUJonRum99RrAjuKZaSGuBaNuS
100UsRBc6ETFRMarzCqHTRJ3y7sp23p9TKn83cWzxdvFqHmlJTJRicljxuMQb2aI
s/yNU1JB8LyGbI92257PeSOMXFTHbqBSOXWSTl+kZPFex2xlzU1ZHLCNaLj6f6C+
A+He64BweuTnPHbHS1psKfliqIZt8tZmf2n406UyMR16JE53jdmFzmjZ0IVZf82z
wX3Tih+KKwSLR2lKbZCOW5N6IjAclweliqq1NC282o07nAATkyJMIvVX61AeUuJP
Zu0cUjQr7r05b6lv91RE577zPrU1MXNVsnOPnzTSTSozSgsmWhGApW8yVatQVT/x
e/9y4PJm8/s9jIUAMOcUBHGzikB+uzEzFkO7rL+44ASGlWxGC7u/iFdcJ2ORq3Xy
5Iq7WFWQQ1jTUfbV1T9LNWUHTnfmTDWNP95YYpHaDTwa/UblBE6PwbxlYQvTzCca
MbZ/kEc1TzUcCR3E54FotyK+mr9ImEVKee9jzFI4+nsHFlIwB8b59a/479qH0wI2
HzMNrOLEcLpsuXcYDDXSczk433vsjC7+29gjxpCOhC9f1z3aMrxXMGOme84WysPK
lQTHoV/0Jj4XU4Z6xEskakRjxOWbYLkdRm263R/LR5X8azjvDbXz4GRXWhp9Zv+B
X8885JdrAgNJeC66pXUCA/eLY92glLwbdt92ZKV8nIDi9LDsVKJyJj7w+zjOsEl7
GrE2SvfY5PaAgJzdvqzIFpvzrpRTBc7k6UDxPOgTrjRrVafNn1wQhAYOVGu+K1Uy
9zfuJMzM587cV0op6Zx6FlmpfnKBc9lJczWEW/CssNwFlFpZVJy4J3KXVVIsGop3
iR8DD2ygAJv6TlHJpI4FhgAplNVvIMfzuIqRYJB9k7bKNEUd2nu2AehCaVDFqWHj
EQh0TJWYACLPmUkEurVUmu7uZwFiSnhlo/XCpujg0VNWgOjPWRsvBEfVPPw4l6Ue
6cZ2k9UoRo185edIotdTIMRwOgAAVU8ACQW5VS2CIW65Sc6RgicerohtyCg58J2Y
4UXiuyZlXcjRawGybo5yBld1QRg41/hldYTyy1FPPYgfc8/DA35mvop0xFYN0BxV
meFGfgivxQ/YQr4lxWx2i+5EeWMm4RzJ00qdbZk3PASIdguFaxS8CizbRO9PbGAd
YBUbFBfMvAHh3c8+/EE8JWfedaCmu2gv/YmcEVWzlEdJzuDTm/ikTpgvcOAZ2Drv
/hyHhwXZ1kX+h5W2haOd1xkYluX9t0CBpGI0IfGzaE+gikfcuVjdaClSv4AjXkPl
bsXZh3sy/6Tw2IwsaQYD4MYBICCdST0jqPfyVJM+0JVig3MBQHN4/KsTPyQ0kHMp
JpB1ChlRuw/6QxkuDO/eUB7GgPYrRQFP7MqZswejG2xIrt6yl3gRvyZjrZ3lsVKy
njngFC8k4PwxpzPdw2mETPrSONUg8GKH44vy2y2b9yVrtJ9ownnUcht+VGqbEpnL
Na2PymgBNbYRyc0Gb32kcyVS7smuZRjGjJCNSSzA8kAzan4e9wSqmnZjin9R81nW
Y7HPvA2s3Ba5T+9A/3NsXRIELGOxGukH+vW/2GrBrYbJBJjvcEhBzDTnKt/fR2w4
MuvTMHgHblVXKzgZRFBTHZkt9qgAu6vr6nTWBFmwo66OBP5iKqFSGnzldFUoZPsS
JaPZlbxGb5kg07SrnvXZ1Xg6j9GCyU8BnT23Bq/HTvEl1JCqgmecA1Ken5t1Q6yT
lhZAgQP7kTooI5H+sDxU51HdPMH6YQSVQv4nnK7ylZCxLYVSVvXa7ipFXMU6aa5V
2XuZJDegLVkvUEDjl/ASRRa1AqjIg1SwdIp7s35yJrMyccfMMlKYChY9+vt0R75x
D3mxzH4amdr9b6N2MIIxyPV/EbCR6d0SzbMSjgmunQLFAd3WTOeQm7bScxgtg/dt
dDatIetteO3q91fkxZ2TiXuArYHKk3xl3sNVyju15OFrzlCbHq/dOl8fkUCaamCA
qwZPU8zolu/MaMqPldceIWJGVG72dPW+Em4EExeWkdK2uEM9/c4x5/4spu94lO/Y
0ztKIoio3f12fY82/g/LefzkcJ5neny1fqLgJ4ZrHdzFaaq2OSHn9v9VlWavDdGS
YjXloM1aiulonscgE0uRA+1bVma4J3+NJCx2PXBBqKIMK+EZny01GFYok3KbgnxC
ct6lpg680Xelv1scFXlEu2roK2922g+o0c8C/a+VGc36ECGMC8xNoMuMenOJ1qTz
T2S+O0q0yed0fgLnfqTKLtOjgeM6YLwpNDnWutWTUA8uvod7z3PPkGAxt1+N3vj6
cENhaMuNAnHcQd0G+FZaZPhbWxVzRFhv3b5Zu+OKQGCbPbgrpAgXUE+GpqY/zLTA
opzV529ju/zg/8PunFFu/JYGudmA/aLnP8KfbkdcQLGkEHmU5vM4VFPSbVRNxss5
/9u37OqhbFS1u+Axo0fVWhEgW88Tih9aeYklQ4Ow+UTE+KSipgosQSoJfp3gzGez
d+x5CpFY6PBMr5TKLV9sNRjwGP+0Hk56N3vjGUI6do07kw6ipF0HELWPsD39XBtY
RzPazLIXXmB1NFhke5Zm4tkMOD8J6yGK5EV+GPFFJVJMG3d8bzesGFMbFQ5kujRE
tiI8aOH+XdA8TVM5POpfytiQwBpggyS9f+5dXGLqtinsR+gAJF62SiEnflTr42Om
gJ04Sg15OB9Ucuq7zvZ80KS91xYpXROR9UGRgZ1j/JnYhYb4yGnGJZoJ531ySRZS
l7/fG174uk1xupO0cbuqQiApSbRJCDwBPDtsztt47RGEGJ81cg8ZCKFlqquXA4um
Zw+6gSefuXSTrtHNpyM+ynxzBxlB2dAIRMgJsGVrvPX6kKjsjQYULLUbUN/XFq1B
BSVHp8U7wq3DAlLrC1zMJ0lzVtlai9h+fgSjJo/qPhPVw70l1ry48iBs47TR3VOj
emZE9u85OOSw3qsZZE/BXOKHH1T1H+vVEKozt8J65s0mDtg/b95t4E2PtcK4q8Ng
/PpRoAGa5MrvpxUbBU6zV5iN3DbP6dDhtW17MqeqCQj9R+6uj2GaJQ/tfzilQ6nm
j4jWDqrIiF/vPjmqBTy1aNKvwMzj5ivA8NCzCsifcz7jHGjdLJI1xK+YBr2bP+1F
ZrYDLeCrBKobCXFcCEFSspNEMw7yngUDhcaKQlSfXJEgyQmOw+oo4cRCGiogM7P6
Z/DXArAzL6SGKQcawIyko0sqkDOuf/6B7wH4wpmUZl94wgMc8Ak+iIqPt2+MaHID
Mq4ouyAdi+aLz0mSK0A/8Qz0PvJnCdGROrhdH3ydwiMeBrqdXxBSWCsErpFZD7m1
lm7NZ1IsOi/EjOK8wNqoCDXEyHK0uF/O3JNKvzhaZ78/67mHb3jLKJKwAx845+VQ
dL0MhGEELTdHi/nlFClhRHqGmgu8VBwrFHhcgXfzp6N1jCbIBUMiFF3p7Ueqsk3I
f3OkInL+S6fvHPfiFhV/62rGrCUq3atrtvFuu9I8C5orc32t9M469eUDA0N46FCC
UW6u2RiKG+tA+O4HD53oDrn9Y94UgFAzS6XOoiyugJXRcoZKqfbPAcGYp33PgO5R
t8CYKEe1WNXcWHoPLotqztHfCordfYjm8qVizgv0Vp6gzSgRPAXmnruPu4wz90zB
wCMIh7o7kbS2lHuWrgHeVryowmX0iXCcFE2AayGsJ7y8qHDelsCcfVwek6/XX+Ls
Rwk5q2FFaKCkksNvDFz6nrakmfeoo/ynpFDTx8zWEco2+ksbb+01XLo8eD+6rNNs
GNuY0a6yCx4aRC3kQmPypEYEuxCEPqSqJgVLfa7fheRz6NSQb41dWigmHp+NShcz
12Zkkv1QVcbvmJJvh93Ms/CvzP/J+zGtIs7t6NZZdZjFITHwBxuzdglIws74MP+K
R00KQJpnIwx7Femz0A3DKDvSMnNNBZhvpdDadsE73j3k092rUZ62jQuba2ef1fAi
ifFEjSh4TrYbdc6l3YeHv45OcDPXiC2a0YB8pT3NOOtTSUUlu1DcpNJ//hpskbwj
wmBeSUYS1GThC0Km/EwpXEDbHuFVQOyZpJDkONk0YYJe+dh6jCUJYcqcYAWZ1H9G
gGv+6qR3KAvLcRgjQhCaIHP4cemFeP9sqAbi4VpcpO3ur0Enyy6U4Lx50Xf1bZHL
AdsSAqYjkHj5Jzw1MTcvByYVghzzgTckI1LB6RwYXgqFlFe51ZgzEupM9jw/VPiE
BKWbZ9GA02gyjhLAv5PzSmRUjrs7NlFZnTdtbhGkuHfEpSPmVbiUAl735zNYG3U+
koN1Ce+ffARTAy8vyJy/yTKe7OU1mNiuCeUv+APc9Ni7LusrKscgDdquO7t7mVeF
9HzulnnoJWP9/HBSVNeqel3lXI4juoaqDIna90151Ksbdq/rdqcvsRvF96SNlksj
zYP2ZHDZTwi8vajGXDVq1V7nso3/0+VyXg57opVln7ZBXZ01UsIHWoy5a20hjbB8
PlwbW+Qp56+agljHvZY4yaVIeEnzULgTTpfHL/rZxFAJz4PcxMinfq+9Z0HbelpJ
FRv0RinQxbPJRIPfISd3nHWxYbV/uHlkXaVpt9CaAU3LzbmzV5uysgilE1SC9P4v
gUWM4VLfxqwIb7gyGlRIefSqMxc4G9ev5dZvptU7/lPJ6HH05il1uG9UoDmrgSDV
6XeCcDf6C4TGdakPzX75vdtrzI0tB7n027qQHQSIYlgrsRPaAjJn3cESZ2GIIh0E
J2OK7h7H7arJQDp/KkmqmKiLciWEiAMPjKzw50p71oWTr8qCid4jBdzaRqJHRz4y
M8hpeyx996qTm49gic65eEG3IJpVfIuI+0c/VBUhvW67FT4E002W3hnB9JU/w+KQ
gkLgVkKKxgca6vjEQvnkT7t75uV9s6x66Gv45LRGbbZ+Z9nDfv2bCtKvCSxjMEZ2
y9QLjRPmWQU6gzE4+Z3yE+hg2aleXtDYtYLvVxU1PW3b/xNSDu7JryzwGIPH/2G7
Z6OXogrg1rWIV20B2HVUX1QIXc9kvJ8ioVDeG6jjGEyUkxW+t5qK1PXgg6bC4cXS
jUmk/lqDSbasbZBIlxPS4lYl7WzFK2aLR9gT9XauODy141kXXhra71756S0nve3d
UAzoLzf4JhdX/Cxxr2JLUawoM+dJM2udPEwPDScKQt+VO+vbDZIq92DhivWNuyQb
2NnXQyLhGN8ajT0Oj0H/y/NlN0zN8XdcnEmVua05Xy9VOxVoNOtLZwj+81AQ/Xd4
nA6WygZjUUnM6KZw7CxJj+2N7/tAHuRXGoEh1i8sK7+7iy9d929PdPozBPnT6KqM
CY3ilJG2nYWUaCpSXepChCbp+WbauYM1Qkr0FYfF/stttaeWflaqzaVgmaYZD5jE
b6KJn6vggP4ifpKIGYAvHSOEVhmgrzGA0xzE26P7mD/11/NzDAi8X0Gw595v7/+M
i4/N7HVw3TRDVST5XsKKEuD81aSHX6oZF5SUR3DXKh3iagnBv3yXf4D+O/mgMfeC
vr/Lo5AESXH0mUWekRVbCQlR8xyoudlszneYTYNCcHHnPTlfaK5iDvCxcTRtTGYa
osT4cL1qJqRPGtyjDUox+U8WmxcAPhHaYtoojCLxXNA5HpE1ex4PiPwGmSvm+0U6
reUpO0rtqcRBLjIDGAIs4YTmzHjFo2vpgNZD/9O9ftrBuNp0w1OTX7lgVyn46SMi
ylwouOQbdnBpbvo8f6FdErxE4kxcBFgyxT1asUeacAEFKmvduyEzvhITSi736HuS
GO2tabjY1jabuRRFMTwyQanZ8bQQkFvA5c9QblV7YJJU3FoWU9hfRmpz/CuZ3Y3b
aAVwMc9ZjCpQEF/CjUv3ofDCQO7qlhOVfSMWnI707HFcfIqa9N1VUjId1sx/FQGy
6VhRJuhowNkD+7dkioxauLjxKWLewuubd/Xpue2xfc9LO82vCZsbAqdI5UjGArG5
/UAmSxf2zDhdAYwuRoOp+W3poJBfS+eo/7VU21oa5/B4bK9mphnJVy+GKknpDkcC
gWDX8I1dH5KeEec3kIMLxtMLWD84G8qWWh9R5Ook0Vve4Lpcqnvij30sMRBhMnJ2
39QLZFvytLUbv8tiOqAgAl0B+VPp8fk4mXycdZtDDG+7X0z3LA7Q4IIM2KuSOIyp
/i4o71eL38CEZRblAV+tC6vi7xb0UIEeaOUl6F3FkNnciEvNhJbkB8uo5mIWJBce
BbrtGbFsGExUPqigsy+7N7/uD/kIQevbB0bU94pUFdmXWj6GHUIXuKJwzx+SZP6a
gML51S3r+nCvfjIAs8Ri8LSN0r72LXDOZmPXSJo1IyBSSzkh1SQPtJ4Ae1LrwlJZ
QkJfWpkIp53Tn1zZYJWc0I3hPpdr59EH1OCDZSWBfpslQb2/eGntfunVtm1gCzO9
ESYFkOP0oDig4C9ij+QJa1PLm5W1SoSP4Mu2uRwHdwq12qG/MEwkQ+lbtaA6OOW+
fhFdU+OxhyoFbnj1fx8oE8fbA6UgFqIPSlsetRpC15hek9peFgIK6T75vj+guseG
RElY/xXGPYCHv18md+WSst7/GLerpIWdzZNj3CAAt0xMnU0KJnRfLjd48pmXoiHn
/18R1UHxW2gXZ9be5NGF0B+55ey4yOc+uZPE0BPB8LwoxKTPQFzmDVYdg8dum9Nn
jVd06dzdHWQIpvnAlARttqVCc4cbCUI92f4dWXiTg2f4U6PxHqMzsIAYGKPkx/l9
MTaIlMJ1C16Hdmo5J3/ppqMjjS2IAfede6LQ0/mJ+IiatM1CGAj4ErpGaq7xVX2W
qs4uaUFRlVzYIW3xljtdw2uQaQT7825NHy6M7Nsaj4onFegQ8IuO6+l0lOwIR4A6
zi7fK2/nLxJgxUaYHVfBnlDm9jgUNR/6VQ9TWXycuH+gC8ZKkclqxNAP9Um/JPoM
00FNwmCNmzpYBheVtLwJtCvtdviP1q2MPjDJC1Xse1x9/ADJh9xo0f0+Q6cDumPJ
D1Hwvpxn0VZcb/0jFIml9Jz+XlMNbZ7W3dzHGEqhKI286kjurA4hB1tS9tYg7vl+
NTgEseWBRoxJb3zUjPdjUCes5agoH/mW7KzA+m/+AbxfjzWVnBdURlvn1Jp57PnL
Leksc0DEfw38ifcMxq8IwtwRFFjyzVRh7vDQPYCZGZNCZYfy8Uk18S9CLRgDESP1
BVN67ikmGIleAteGyfE3IIaXgyCDEvXiyYQpXLlWZo5XxH7UsTeDT/cZbc94HHLG
xAKjl7AJiEleoysVtU9g91AT451xkNRjUbt4sXHkeGPBEE+yKO2xBWBYqP635kDQ
ci7qxo5UDvX/XNZ5cC4nYEPZJdvAxIL7GBdw/FUl9CCuJbV4/GROUFE3DRap+uUE
28Nw5Y+ZNCSBN/tPRKIRdj/BRc+xXwdojqcNfEuBCZ3Wd7ZyeojAJOr50Bdwvom6
F5rYSAxzWM/LF+oew+Ygbh1Afu7KyEYa5XohEPCVQ/1pTXxKCYG00Z0n/n5szRks
jCYuHWODW9Ax3PfRXtcngSLjgjfgdApDOlqGVpZMl62avXWOpJ8V+NxSD2H2JSbN
V4M9+2x0r1S/fL3n5Ml20XXUZDVxE4mtE/P0p9nlQX5fo12TyjzM+H/umnsXySWC
KkqfLVX9QH/E/MZkl39zm0OmTZRUTXW5+k9altSX5NX+ADc/MrDt3lqgtu2rNyqF
y5TwTKC3KkAxHbV5M1FnD31PoHq9O+dZPabQhxxbR+IropriRxwrnXkxAzEATf/l
rYlLFarNAr72KFn/DJgeoUUzPCWcRlZAY35vLCzyVCRNrGdiLPnO6qocbfW4Wx/4
YMr0sKsYy/8LFzE6fJ/CW10zGR90JCn4GRALmp0RVmnHIwGHYckYaN/LcDSxzeO1
pZHwlWB3Rtrc3SlN/OEbUqY/p9IQzmGA1wVEAsIlkZyBjnbLTs9fAQhwCX9UaHdb
Q/5ODq4b4wWp3rg2DmTZLIL+PBZV8aItwYF3W8fqsuF3+l3SwkuQxb0bmSrNgbFG
AjzX27hm/8Jgw82jMGN/k3nYOeHMxfwgZD7DIojjPP8nIsszKNajN/Rp2CfWvmy7
sQDwyy0wtXD46KMsMUaZObuSGc3UHN+QelySefjZL/am0DEVzbqjh+fHDN/Yceup
a8YoFDZcrArhQhTiKKZIzZ40+NY2IimFFjmOjTXQp7SSkdYmjNsgnQxYYjOsJ7DT
KPxJzbu59BqyJi6lVoLnCD8tl5Cm72bk7YtwQ72EXTpwaN7qmrAgz1wrAmqyPnqS
xNnCybe9v6kImVNhKHFLNc+WQx8iTZbQVtoVMj3on3e8EIE8krcYj5IFbEDLJbu3
8hMEZlhy6cU/5NzOI+/ghUMK+xsdQKNPDBH17NzZYyMhB+rKZqsksa/KtVD4gzCz
1sPv7L0tMPBow7h36UhQkWcxBLgE66VLF0I5qUB0CFMwZK0UNE/NaOss76dhdm76
IKy6Xyz7VGOxa3jgZGJDaYJo2cajLAxfAvbFS3Kg2cI7JadY8Ss8aohE8WfN4tTQ
d5v54tlqs83GL456s9qM22llHXrgFXQXXwSmSs56J0MiV81G+ndYvjCpSEegF2sf
Pjefx/wAaXiuzxdXjtsTvM4pWfJGwURPSRjOlIINfNSurtPZfUwPdhXdXKK+yph0
h9/AtMpq5t0s/S09Jrkxt7b5W1Xr2zzkqsBFgEjCCYMZCBeOOHO89yDmAt4Ur610
BQcWoC2foDTyPXQ6cmyclIY47v1jUsou3q9ZO3utORLhqRx8YgO96VDh3jgKt3lm
koc+NyRmB92Hd/wvqcNFDy8wq7KAAA663f1AgfnXJsOnIsWIwLEP075PJA7iKqwX
HUvJD5H9xvCDw3CwXzJuB3dOWC27/Qw/3gjoVfIMcGO2kGYfvZFh+fYXIv7Bztkq
WoD6ijsMKUb/4COR8LVttr4yzvgGSL0N2nHacN5fcFk/FK2r4JyAlTjwYUvSKei4
XDgZ5+jNAjj+XpXVj9c74ErMXxDfIYT4tJLcFOpQqT6r9ulRFQjZ5EIFWkt9Ubu3
m8TXyvVSOWIevVCFubj6um32JxJyr4I3Q44EPCM3Ydcc6d7x3VKBfqurViOlHu7X
yJDnYMTYmA7W2YRPKh9Dm8U1oD2XUGyy5bf50Za54QR4aYiOrR1CZV5rJiLyzc8F
uTBr4636oJYaqFXbFDXaIdVzLfvYzuir87/uQyJieJC3o/BRVkui2+vYiL0ph3OU
Ln1DwuY2SDfZ/nY0aQ59iLFEu//XaJQeVzHSPrYH6AaWobwP2efr76ZNKlenLvey
tmBvloW/lyhloEFLmxTh+lsKGZD5jXQUo8bk9tq24unee6Mub/D9WnJWmEqC/GbZ
tjtos/eaQ54etILCY+qk6D+RI7zfZl2ILS1sPB2BzJv/vg6UJEjkX69L+/trv567
QKieYd5C2rjbterqpPR1TeIHFLkUvrjvLARw3FhYFxan5DbxIFwcry/91oMOyXLw
41Fr4uskO2KPDAf1OT/f7yB+tNbFq+7t3EY5B4cRxA/xwUraOBun+IXIrEnIfsz8
2D1D77OI7EsqBtmPDSR3VsXcm8TvCpoM6V9+REAjxugpjPU4VRbHRWpm0GKfs8VP
FhLKITwPLaO3UeJcDHKIUlhRmfeFfd27E5kB0eTGAVm1I04pyuMgO4j2i2JeWabH
OnerxMGozdPyqw6r2dhu+apECmxvsekUimRpZOCecF868QWZY2xLWQPn/YrodK3x
licS4m7oZTU5944HjEN8DcpxmaaIFaSmZ94GdS9O8tN2p6xHYAnDVfZ/tG0G6xjS
wd3Scy7Y2Y8amRBKGQ2FkQtEChSDw5ObTP2Wjn6CoCaL1wkHCFiAb9pNKH/OZ/Oh
C/7Dl36R0Liir/2K5rSXSeM2nOkWivIhXyHwsyn5CY4i5UrS4N5tg6mDAs1TxpZv
POyGGgV4IDaZ3v0TQINtFG+PFvV2P7Hfe691uEWrJfC93XCMlW3Ig1wU+RKX2HHm
t1E9FE+l5AzPxfogOR3jEdaVUqZIaIAHmKh0iNmfx7CV77wamUvcyuxuSfHMgOhf
2xUHRBGPWQWqFFj/5QR3SZpJMCCZ7m8uxD2jrND9sq8h54XQc1koWcj7qhR3OOKL
XoyoG5pYUCndviVdwwe3d/uAXheFf2aCcUIBRWmYD57Z3pspmh8v4sKavo/0AgaE
DLXBT8n1J1/QgRoJwYOKnZkNMCB6iZQK3wlohJz6Hmiz3y9mhZ6dSOv3NP5hu1AD
dAfq0k/+x8uHzMyVBUfFSyw62pMzmIDoM+IlqpWdHlKOfv4B+3gzv12jE90HUzh+
tIojxb0z+P5sYYKR8kXbMrUc1oPQu4LOZ78xvUKj5be49vkwf91w3w71uvXz8jLZ
eJjFzMhuhMARBFOuN/bmPw9TPXnH9owBBpQtgxQCm+Q00Gdkun07SMFnFjI1dDfd
kmvqvfPcJxx6rL1B9Mi4VyTWPKJ44qt4w+/+eEGfpY/5BQ4vrCMnJkziP1SE1M0Y
FeZ1r2GqLsMiVlBvTN5m/mpjWvIs/ye3zgZn3vzAVwQ117Jyw+3sJzvHdpUSajJV
NGlgQrtPMIs3RzCpxz2nLttFejXRkPn/HaIYbEm742J9zYWl7d//VgK2rMlLtI7T
+klFMm7pZBqZ7ZVPpXZJqOAkwDp84/3cbikpQFswe2mDaF5B8b/MAEpQnpm1/88l
ydDkQqijygSjNy47mp0r4cu2CAGf44ojeIJXCOSEVxsGES7Fl6kEVsOnUChumzaR
7U8NfpejrFboi0wWefAv2CWP88WOatPrK4QTxANz8w/E8MsAXi6ZAqF5x5MB20P6
cAyLuvYQz3pGQSrwHu01TD23Hu8SL2ClK+2ODy3DLsLAPdFdmwnsISnGkcTSRlF0
/Zh42dC19YfRZMqrCHUJ1/v8yOTDosa98QVijKFSYnBEHSi1txxlQ1u+jBodacpi
XA9xluJlT1RE6+/NWZH/gll6B2CHbCMgVsonGuGS3J5bIqOlvypm+GizAV39cVro
VXrWsM1SBIQo07Hr181+bidLIGhCqSobjyjMv4ntB6yi+n64MD4s/6UW1gzvhdoG
NhAwEHN387fBPVyDACTVWMOUndgmYxz0JaomepRVoQsQL/sBizshkFpwFvC+sgbp
KBXTkyKKRW0UZjeMtMRIxxaLZR3VCN1WeVIOO+cRyMMVYNnChpYVmkxgMaO61X4L
PSM3sNgx44MpO3QNR1sOwVtcAhmnpVRWS+GM+TQSwouNQqEXaQATqWMtHImOpOR8
nXGGy0SygR60TDgAw78uwF8lo/Mz1AUqt5awNEwxb6TRQhOFdLUM//vwQ9Hmi4wE
XI3uGT7I1p0FbGE23p+knqy+UgV6feql3xigRVYC6aGj7WXcL1WXjQgtOJJCcZFQ
RVTZipbd06lQcU6UYjwZ5jKZNqR1gqzvc4LRDmTTP/J2wpRnYvkHjgaG2por7Rod
R4jrRT6iyiLwqu+TnyntYDQL33SnTpShBGvD3yvIX0r0SuvRG1+PwTBGFF55q9d3
kFchYca8sUcHGuddhhGs8yJOD+54r/vZLCW0Xj7au8ghy3XeVRHyCKrbm0dcUBYM
2vJFYuv2i8rV5X7LoATVpHKtv6FQMxy2eJ1Klgo3LkdQkfr+VYQ+2MUqidb+YYrz
l83fWF/wvOP39fE5CkjVbRALragGlNdBBz2LDRzCT6ezd56l/TvhS7m+PVj0a/eW
g1gdAFRCtEqPaU+6VO9+cdbqJ4w5avPs3Dg7qFiCQV7wVt3/zG/WaDxrNJTyPJx0
n4uix6bv6g0Su9FfeFIqT2q7tjueieIa6TS0gjJB3tGdFlJNwa+yVCYeCPthxtQU
1zNTn3F4oVG6AbCmggavulDrkXUyBSU9yl91VS+RTBh4RcvSNTEVRHQ/VzmN2knj
3sRSlkJnwiVLTMUXyTQsmwClzpjcbAixApv2rMMj7tiocK0uvFOskVXP0F3EKxF6
4oaSUBNwdH9ye8VS2YV0V90C9qE9UgSy3GYWlGqiLGgsMXrV32Ml2gzmaySFx9eJ
nsQYtKfUhqpLfq2jrB8p2pY1VQtGA8whEF14cpO55Q6BBc4eAqOnpSIiusOs1PsG
gatdyM0bY+h04iAfvo3anjSy99Rc9lPi4dIABeaFcKRgGSqOrAv439mxiR45B2sV
Mn/c6Kyi+CFclqUMY6Tjuc2BrOGrYU+47xA7ibcePNyMDjFpXFN0XJwkXmDIo828
RCHLHxhZeRB7l8sW6vUGjvTQz0Q03zJr0xGwISyIz7GMdKded1vjd+KAR/q5Kn4J
R9Bn4M9YAcMnsTBPsXWf3R8jjwTVSVS1dJ2xtRQ3R6s/JFJOcTPfX2ntc0bkTCeE
nE6iBvoqS2glcpux30nnlLXEjsN7mA2UvQOHs6qbDSiPuwm2okb+tza9/GUKYpOS
ZhPjayrkinB5ogPRaI6r3UOGD0HVYHvIOQVZGw8+10jUIvSZGksKunqagNl+0EWZ
SBJLduE535x6DFArxvTz4P3IERraM+RyJeud5HpOPeucTMvYxtkYa8qzlk6kkI5l
1hOEcsje9tJWZM0jWKv9EJV8j+7xU+My/kEznvrD/C8gJM3LgitatxOs9DXiXRH7
n0krBLFIZDqV863ZIF99aNJ2vCVLeWYlNM9ge+FLUOTfMzw3hSdqCQLinFw2HyOW
HwNWFt5Ptsefdwua3jd2mRz6YhlkvXLo7pYxkTZsYGwSf37sTB6RPcBN/ETnWPWw
SaPW6T8xYfAyAC4ZoZGpC+pY6MCX2somDYsCORdWtJyEpC9j8jAiDljZmuY8yPjG
43eADM8obE0ipAIuEbl6NvWXOHM8oC44QEzV7E/iRNb6xxkMSDyDI6U1VT4Srm7b
vJjY6RBOc4+hJ4ZalpYpUdlu46UzzrZCRBGe18XmUni+GgSoAQoJ+ApbY21iAuxx
lmumu+FaD8XM1arBoL0FBQBZIL40Zy3upeB26tVOH62TH+QoE0jhlEndykQ0Yvic
s1yqqwVFLAQn2CJBPeo7eTwU4QDlUpH7fxMBTUv/YuPDukMGuPD48sp8BguufNzE
RiwM2XelVL7NePkWdc6KAn08Qb4T0O01McwPznK5jtB71tVIyLNTRXwELS8VzVqR
WUggmlFB8fAFmrgaLL5B3QUqz/Q5UEmQR9Ef5QAvPXk6laK+JJWmXUsXrlh/Q7iv
uw7quYOEdd3gc9oj4T9zqd3/uqGkwhCyWZWlmsXA1YWgizFY7Friv5i0DGx3TkKU
KpzsWPuppyPOXjiHgwG0Fefnn1JwXElpjikW57d7VeBf/5QGh9bQU11u8TEzsCJF
2+iqFVfsmE9iTJ/EE4OWyJIeaEPBw/6ELL8P2i2CrkwTRpwWzH1E9KRZ/6/CG3HA
OENFDkTXkyVvCCt2PZgnf4eGIATBQLCbiEA+WPfK2ovavkTym3tobErUxxRgcfI0
0M+0mfxxmaWFWr88LRIqX6TPW2Z+Fy6Df599alt2votPyB/b87BOqvcha1FvohxO
fVwtQCimjMs8gThbvu9FV/aN0gsPf1nE3TH63UJN7czSG5PbhSVqmOpKpUHsxUHb
MEZ6aywYZ+Iqlz/XD1uBbtatSx18aGm7uvSX7LoPwLoAUN4EnQRePZEoHJbTqWO5
Yk0DBzaCPPnuf7JFpJpnttiYdyLfgptY7IlRaQjKRBu2WhJ7w9Lw02/5wat4vUmo
+erKS84SDGPAGakRUOoPLV9gcO00kFH47YFXNw09Wz/GEpRqmF/COlxwwn84kMIl
D6QQ7lHfXg5UrhfnMSFCZeOyye4WGA4rN+HkDJSVjksU/Qhx6ak7g4YPS7dfvS14
aqPAAMxbVpYu2C728jWRnxLyWQCA21PaRPx4n70awjMvkyqjMLhkUmKKzFvfG1Qn
w85LrHe1ImaDhGTc2AYNVNscovd+WEd9a5WYeCCUyQpUeDZtc0Pobim51GpwLdUy
CrxxcqyjxT4fwr4O+ZjMBm8ro+I3fZlIdx4k1CWWTvP8Rv2t6qvNK7pH9iMU8Aiq
+s+fVgcji+jxYK7Cl4iIaSXWddYJrkhyxwLqtUBFy8sSE8wXfuj24xz6ZsDQqWne
xMFjORfOUB4aVigMYrqVRm5uKtt40QgGjeh0Tb83WCt8w0cAlZLBwY+x1DIogBHR
GL2HFYntmMNy+SYMWwrGk4CicolSKN7bOY9fZd2Z1htcWA4MbF/o+gLNOl8c731X
kQzpUGgMOIQUboahn2qR5CvhAnCJJZYFq4Nf6tzCVSknLO3Iis46eYTTrVwd+Ujp
kmbhZxdpl2s/G1qt/VncutSvPDD9qXkMKSC4/Xbw9HJhGXQmER9mJwAd9SEoFmuS
6T5g1pQZ3xdm8WCwvH99PfSXP8Y3SUkdqzWjWYBv6U4cCHdeyGLu+n1jlBQt8PPj
VIGkyluikZDYJwktmgIv2Ef8nEZJbHObwyNAGfwAhpqeuK/hyErJgE6NDoIN7Tih
1uMXmU8JJrHQTEjeDmiOgEBnhZ9TEepthg+/zrAx1DA220MCPquYr4dm2YxbMyc5
vp4Sxstfg28ai/hzShM19yhly6Y8rZwqUFSHXACHr1E+VzpQY6Day2wnDcxyL45s
IlNDnrAcklYOPhbgFKClwTEq07cLmtaxgV1Av1sR+j+TQKr9vUSP+gjigEhfTyMA
`protect END_PROTECTED
