`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjMpV9d1Ff1B0EVlXZDbBAAIFk4vigGtcNKcLTqqnfqV/keYZMAkb0l7iT9Z7x9P
K0cOqZ9vKfJDAtIXdaoYOhFJtXaMg8RLguejHxP4tP5hZYcbua5To6msXnWsM3+8
WnFAIclc/9fbsnLb6D0Y0kf6XwA8nL9clAArVB4VcV2xcL0vMveHfnEyeQhtnaN8
xXjuFjA/erq1kAvqJmmunIw5uALiVxDK3GoYB17Zn7HHWXZZ2HAe8VwHO3GRojWH
2e949/ziOutsDyF1+9Sij0ElPgMNQBUDHuhs7TLLQRMGfwG1zyJYeI6QqW6Xl/Zl
QV2Eh8fbjNmUGdZEJQdRfNIFQEG+jFuSgFqasn5OLy9xltZeQjomAvb9WdiaWvER
vbV9qtH9KxeNb9gpcDYPCHm766bbM2uk624lP97AWa/+Rq5Ayjd8nVFKgXPaayVh
`protect END_PROTECTED
