`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QyzSWV7xDpT/k3EsRokfooRc4WsaWR8X/Xe9xkKtWBKp3ENtJRJRfCOTk+UXels
GrP9tj1XMVKUcYHLjJcEOlsoPM0yJJ2P55e8+LQCWAtAivq1PJ21LPmT2L2Q0iaV
PzRdhZJChI+OYQRSiNTJyxINBb/XlvOgIcZxRjuUKhW6ZaKUJh3ALZtfW3zciQ7/
NLWubolXINKsHLLHk6YuEn2Yuwf8q7BY5crHI6mbsojywlNdXWNtP9aSz0jdvkSe
RefXOMskC9CfTh3KCWbCXaP4bfTeP8cP7uPStjVT2w0tj+MwL8YvtsWhHH8FuhIZ
WeqVAG3x6oD+47pqXtHQ3xV113ankhkN3QRBubderi+JEetBHfCjxBlXgngn/g52
uMxNmCZ6m8elhNSBBP8ro3KTqCXm2NIq13uOnrkZzgAHlA6v87IL71bL9PWks1/J
PKskd3cRTuz+QlSka5CaPSOya09UZyyoO76P4sXVLSZMxknFv4xzT3dKCToTTYU/
Hj6i11cRISAlwJNF7JPb7IT1TogRfI7Adpo4W4dUdRux4yl/5jhWrxueDAclCpz7
UQrf8qByTG2j4qDIIjNTNb6bvFurDGxwGzzg9VCdlxVLSoO6FJF7a49IhTLL07Gw
Sm4xzN5jSVDqDbyq2dAgLP7Ry0fVjVLP57GZsZYqiY/GjU9WEnH/OKld2nwJvZ3v
P+ThInmFPUViKQYyWp6ryerkUSAmfXRX6Yk2aRnsHo5Bwh1mcHiw6a0ZS0rLSvZf
c7i0kpNWV5U1xg7E8OKxlwgxlc3TWIK9pSC0X/KafVo1RAVEW3tSBuaqG4WiGEWe
xAlptL6MlWIU1q4fyA+XWs24tpIBq0M4yCyKXw1Nyh+Jf+dwh8WanmDlzgl7rFoi
pwqZv0vfJunxxSiUmCzZtu4RPLgmMJIkH1oFX8q938sHwLZX/GUQcGM7ZNKAOd/5
4w/qH5YUYmcOiQ2TiSXTC1OlrbU1Nn3oWb2nUQ1pCilGKxSTsZMiTizkUzqU8GLd
wjqpwLui8fzYk+t/35Vn+M3nlAtio5uyYCMDb7gJgcD9AhfnjJNTf3ObCeas3mCY
0jLBCyt6XN9zfbwseqqZgP1Sr8CHjoOUDrLeQb2xbh/HHckuJnDbCaHooEV+iZgA
AiPgXw5lzpisShBhTF2FG089sZf6g9yLnQvtAZWJ+RiUe+c6+f06SYTBWjp31HUE
Rpm2kdOMDgUMZs/LR2AHS5qgAoJg0rLkT28KT6boB0LzOUUIiTX8wtes/P+JH/f6
u7t2eIRFt2OGkOYATbjNlV31C6V+eKnOeyzNmQ5f86Hp5JF2bF8eD0rqt+hTxgR4
fi6vLDZTqgeTitvVMcxNNVQ6Fn42w/i8VX6kr9Q3ne0681J7T//5NnJovcO0TOmR
zQIeD4CA3DwP2PWItqTURFpCdHjK7T6Chs9LExdTMfyIQ5ToSAj4VgtloDq04HnG
xZK4qHOmANRowOMSuUVYT9DPm5PCcZXMs2d08BPUBO2w1kQUJ+Llgv34BF2auMej
fpwHif1wqDhFVIftbF4/2FzzZ/UIafEhzgr0g9bIs4rt+P0icWQkCDe47id/p1QY
stHmGj+Mdtg2WHduwd0nY/R400J36EBJsts/rr1WZ7iYkcmHCVhju1mCmAHkCyXa
g/Kvy4JJMrHFu4fMlqN2uKSrj3iEEGHayEvRcv8h4Z2y8Gz93Krttdmv7YOyqLvv
ybOrPQjZQvWvMBohezjN80C0ZTIrPVA63ip+Ea/pVKHcEIVn6vVwZT4181FVpmSQ
0PuxCERj03hyVgODlPi/3L+9xSCXWpM8FxeKWr7ooACbfB1Rx3d/TVaXnpbww61f
2mzAj2pHDbUJDTMq2hfOMnged1Zxyph8+ohZ/6wjLsW+73zel4zajpbW3+pceqeH
3aTZFvYP9DD4nn5PqsA8S+RikUrIxxLReZHFA9D8/rZuv+fXTjmrof6XSaEpbsNI
ByhQVkHnIA5+H92pTagcUmisE8TvrIP4AaCod2slLGIKWOWGv1A1WciKHDtX5rQf
mS5Pa3UJAT3rSV80DkVH9zPSGB9h+jbOY2+os0KWSq087IzlJdFk3k3iZXjqcow1
rE7DDN+sA9Dbld24Qpau1XuFF8MBVNEZNDwiLzPGpPhb+LmdeKu1Tp0qznMvkOBd
500ilzqagBRtwRifH4mPXVHCVUkq+g2/P4PDX2C2WRu2dMpHDcxedwQoHmTIEN6w
CCBun3O5F/U5EQnEhZXOZTkuwtBV3FIQUfrFuvbPouyw9jOwuX6dwYBD3oOt29iL
Fry/3/ebBHZFihCuU7uJ1z7EoVlzs71fwBiHN56hW4PpgqzM0U4ZHacUS2GaLcfD
t+UlQQYUluvvNA+lZJBy6PqpRhwhOyfMF/lwxxioL0LACfM/ix0GJcTP37AR66HR
u48J3Ce7AQwXTTLGbYlHP+i4KZ7WKACW3RQ0W1MdWn8bO7pzc+TfobN1xUVYZ+LX
qGGn3NGu9WSSbEWLAp52WUfw62pxfuek6Jng28L+yen9BRsymiZg1p84NCdphHY1
AqE0Fdl6MbxnIUFgOoy27R/7N9dqzJoOlbkOBeoawk/bC3nHXX4TmDJHL1X+3pT8
5uNC8XNnRsRSuDeRJysfnLnly1LViek9P16sWbydXaGa7kbtsynScTDr3JGObF5x
Irm31Iw89+a278nl3cQjMxgEZcTxwrrmwL1b8udWLk1hS18MZ+2dHfgQ5cYIeQ9p
8WRdDAqtNZFBfch8D2pccSCS9XzSUEvWqZvN4TM5IzXz3/c6hZ30RQA/XM15c29C
6/19DXBaKPAwWwOLtXT/7nk0OtJ7Ly7bFAsaguBUHIcu8zKCHW1Edp54XfxPJiyD
tQ3Wd4M0EVxkYYYsB9hfhMfik9CDPAST/CZ5P1tdmQxQS3wAEHMO5x/fxE9rqCjF
QJ+VuKSJ6QzP1+wlTY1h0Ti1n7vi7XsmRefVCHRLejgAINGS83xc5AOWGa41xNpR
V+Q/LF6B6PZxCeO/mgWqGvsA5hw1/FVYZW0//XBLNXmjP2woVZ85J3/T47oTXL56
iXd6yNp5zIgH7MWecSq4+3MZZLVVo0udQSYS+LrmQfFmtl6voeQcENZjMzTWDFeK
lUGqlI17NFlQQ1+fTgDrjpq5scnJEBxJGEYgXoyWoB+YJbyR7f+V98oRxANZk39q
2hR6oOvfmdhNNosKJgTs7B1mEakH9DgTFD6BzNleyScOmYeb1E0EZ7CT24lIx6NE
UmPZsRd9jlgqPlIPpxOcn6WRqR7Iq33ZZaKnYmSDo+5VDlUTpHx15ihHHnRbGn1d
mrR321k6rzIKc/U6//MZKwoenMJPMoe+/kxQNn18BVHBhya22erqDBXf7PKqo26b
su0+2o48vsy8hn53/inVrk25umzzYQa7r6OjWYzWtQV4ciSYss/4gKIL8FoP5gZD
qOcNjXt23rZ02Z9yW9q2J2fvWoT3vkZoxbqcLyxlqxcBqEbKK265yf5mVl7SajKk
7SGYMvLx9vitKSoxH08WMISdMp+mduozQnFICHkD/spWTzOMXGer1ggcTZWN+OyB
k6X+oyFyxJjgW7zRlaYCT8nUQro9xgA6xLPsbQkbwdf5jyRXaaahnPX3wDPnfJYN
lVklTOUlZ+aUUiFOeHKOpZPlvQrJ6JKKhcLis21KmDhrbcB87NGc2WzQuWbYlSF+
w+tfsxxo7Yek2R2DfY/NsWfIZVU5q8eURzWEEt/RcsRCTbZB7yjIEZl79eLvbe1p
jvLAjbTlXkVjKuH+Ba1eUmHNDJvbBk3QbqqsjoPNWTt8hoxUI4Fj5FO9zUNNN1KU
PisCvtHYO1dtbqubFOuqV7kz3w9hFQh0bmGN/oZCmlg+CR4tcp0eF0IWuQtbIxZF
1deLGdHxqMNdSX8VeATiVRbhlWUOxjPfaKYNMNPQ+EfEsNWr6sn/ubWsEt1pPiyY
yTTy5f8eo9vtMyEGGbXRAmpONVFGX44ZPRY8thZU98vMgYasncoa+gGMOIIQvjbZ
bpWGJaYNeBfY6et5YiuVuwsrJXP1hwPh6RKI1UAhGjAHpQKM1UQEMOt2+nLcQrXB
JgdqfgTYEEjQ7fE2vkCHlhEsVnhna6znHNYGpRU9drNr2oHXHzSRIMaW/wgJsghP
2fhwZgDnDNyjXUF7DaJmKZ5TfiDdfYlVeALrCVduCgAzk6ItwLqGpn3yXrKGnKAi
LNJcpQ/WU32xzEYF31v0UlXKmsnWsbZMjePrLIxtgwpRSYiXjkW1yu+05wkSdJh+
4n0f7LpxGIpfoe9jIgddhyrUuBMk3hCJgcxqZmHmekopXLjbhPZh4IAoBO5c1Pe9
54KHFZch1CWrQWedBPtBTvPGsE24wKbhIb0VbQeaEXZJj44OvWKYJy99+fULVjLx
nwNOfunrZUNyG72f4x8/hAM3/h/W2Rc6vyq/u8bpKSw/GlZhBnahjy1/9WmwatMP
hVTBd8x4ZLAqy3Nfs3j5S7Z2rPRcWYTHifnSBoQA4IrgH20sJF66cQ67I8XkFyGQ
9PFDi55d4xaUgX7Uc8b4rxxfi1CiGPDPl5combhDtBNZCRFVvMbCQKkUQB8V8h0l
iYaUED7OvdQezPoSFYxPP3lBWKi8U4nARMhruWldPYoxKkk7nfzFYPLPPufP/0T9
WT0+MkF8t3WvNWZNyBfIY7W+SsaQkRC7zcctwe29DZxDjQYlRRaKSbA7UkYSgefF
I5uue4B+LHzPkjDdeCClujBp5qdAQR2nj70XHTI0SFs71JUOlBTRhNvOzlUV2sMn
kmCWPvyfMJQydxyoSFgb4ZmBh2IL8Kyec3sb5iLo+EIrCwVETsWAu+sMAo/dD1OY
/QmboCv7ACvI1WdN8Zy1StVyOU8WkhL9gP3vyQBfBEpU5pZFQucUWElDZEuX59GF
2RIpulEQW8R3k3eVsZfiwxzXXlBntOfeGemBFmqD/OpU+HAHnjrBbZ4fPEL4Eayu
zVtGOrOWiKrdM8KFr7cAp2678kLPTh4DKaIW78MYQ9ELoZ9eBxhGs6dvncXECEmK
rzxr/6/zzfB+GF6x57BtaoVlm39/jztpZpm3gX77SPSTMIG0LvCpmciK2fOcVvHe
4sNEiHUWOlt38Xg+RhuHgVIg3LeEU6koRhKsgZNfoCYrh/7OaGpMzYrYh1r1o19j
RH8ec/izZiMc7RTdUBJ9AAvJdfZo9eTKIWGZrcpWMKFdD2AubukHFIsJHI3ElowJ
sXHAwuCOmjx1tbOvOwCekp6QxZGNoFuJlqo3a3HUapxF9bmpr7R4f+Slkiusfkaz
xPKTL6X2KjsPAR5HTMiQAQJBaLcqCZm98Z/8GeFkB2DBl7gg8FKKDHildikyljre
74LQ7Kz5lZ6ggwhbjxX9c8OUc4rkVcCPi5LWvH1jN1VCk51GNgcote3skitWarew
YPYn6wi+dGCJHVGB3LS6SsQZYmjboGS8pfQKI9BShrPHwOPmhKVY0klpgF4oRnFU
KiNh6dKs4D4L6pbOK1pUfia3djOTkqUagzc0IlzBZVpRrX8lxjZEk8Vg5Qef74Lo
qhZWOzbY9V3lE4EKdnmckCsQ7LNA36aJqgOzIPomryu7pEBfpTDrv9gzKHG3gbtL
v5iJFsvT2FcrpnXtiB1PpdTm0EGVhXPlTVwut8hRHZIHpU5/fVxjMLvVoMUJklUb
ahluGOX3zQIAjOyxrz/oTlK9gsedWmA8f1PEU2S6hDOqpk7ZgPki+GyTpiROJNUl
QET1jxTb7f33btEtCrhL4EE2+swCeO8n3Zle+NFhoPZ5agFivDbTyTV7Ab4gYzwt
OO/O2jdVbMryNS8uhgSGj6nE7/w8L4zSPFaADqpIMFA4Q3TFGXkUEGwCC7aeoeap
hWS1MAVTUc/4g+DiSCXtMEWuuy9LcpONNEixYi28ptDND1Jlic5TqhaSU4uAktvU
DDeb/rn/O/i/5mSLvMelqwQQi+I5ZZRPwLKeZad4JJYNCZ1c/tOckBgt9R7Em99j
kPUoRHkCZ4ouNcJJHWcdnVWNviQcCFHTGzuFoJ2uiUhOEpQSy05ZOMewTZZiBzIZ
NbJzPa5YioIBAsSRMhoC+QSOq8TjGXPD4WRz1eeJdTZrrx2jzfo31OAy0oGHww5w
JZyAzfvCpW9SGXMnjVfAuonWNjLqSkb8D7rg/+uKrZ2VVEmz4GodIHsA5E9hOaDh
qZLma+nonixUjCdnKED1duCJzesvzvVOfdaL9svbQOeRzLsCLPzx4qFsJyYvzKOM
6GkvpGJRfbbDD3cy2yvwvBI/p5X/OVe9ogPpJSxCtWccD4FfKs+TWgxnxcKLgHPE
gF8l2HKPinn9hCCSsIg0hX5ZDKD3IDLkrSbvBCg1e7RRTJUaGJXUHWM7dv9Jm/AH
Zn4bU4O+9u/YU8kbXs3MRXfHiOH8YfTq4zpyje9CxTJYT1FxB5Iflr0r3LB25cmP
th66rX21BbHArCwnuVu7IJfNKSDYMArpjEizikJ5da62AEP+RSoMEKlNXYlDa1zT
7vGJ988RjZGfvp49irYLBkf1ScmQZL9rFdcjv+G9McJEDkzj1peh5Fk/gB/A7CFU
zbFNlNhzYoWluzzD6v7DewFqsnLQj0A82R/xy4144YSxquddXVZJ2n1flQhh2Zaf
j4qlvny0Szs7zE7P6khTTUHcvUdDKoCzo13ps5FFUsfzJ7YONXHTyYooLmTAjq9s
qch17mGwCCqTxCgTAZttwVjujL5H7fut1Qzmfp2bw7IsawJClcfUcgOhwPH/E4tw
kWve2RAcOT0frIQQxWq9TeLMp/1PeIOsAYpaaKodqvotyuOJF0+e/lZqbrk5wa21
BWxHYpq39ourhajvJ+A1LudH8+5dgHmqsvL/2l9zuMpiNzqkafd+WzrxunOxrVrP
rFU8o2hcMb8QIuHhNqjaKROR/Si6s0LOkcPXS1F9eMpLGJmj3yL9nYUpdDqy+wDJ
iZ+IHUG57cULNyGGam5IODowTKfkd+cquWAZl96PHZpcE14+BOcdcuII1FYozxOU
fytkegBK6yi3Bb5MyFXlIp9BSZUQacKRpnaeVDnRPHYA//Zbrdg3SYQ9dA3Qewgp
T0cHGSUypwutKHEihK+cRyOXg6GXeRDwB6b32lGw+IBTvyMO5qHqJHIW3E+2YPc3
44BRFrS4baYdvUcoKcKXhk+Vke1OCudfg111TNbcyXsLFwfR5dxr1Ly4fqzts7MG
Fg+lmDdmRbh6KkurhVCzA+tSf7LQQzoWZopxmZOrMw8imp/eQIQ5HVVbHgp+NNjL
8xq3oqjDk0MZMn1b6qQ6N9pQ2vDw5u6K56NlljbRcwOFTn4WaJeaEoPBmL0AZ5ey
FIoZkFAM3z/gqFrxIHosqtYnJqLZH5RK8Ixt7oJXGWSe03ozVRkMddQUM92AlAqj
28fCTp7psIS3t0allkKMMvb1hcT7rXD3fr2j4etdcLsOg1dsJZwwi/NOlSx+d/wo
TFZnSmccVqSWVPPNyj3HZ4sibJzw4BjJ0wdFPDN0DMjYxf3bXFgMBKJhK9rALXZ9
HPuX1wbwi1W/MG2RBkFIaCy/rFCZqKR8J3VTPqI92sk1zfp26uj9uM+o71gdXQFv
1pH5bgz7yV+lsr2D3zfg9HqC7140zJEOAjH8zS908UAUvodvDl7G77uAPG+W1tAq
tTH7ban2RX89S/0A3pYU+pqe3xEUc787yJXSvf/ImichcSqNO8MOj1PscjyEw9sE
VOMqYC5adpR3EfxqaqekQLnPZCdcEopII5RBpPhcV9CY/vjExRYTZz8W67wUlkRX
GnJH5Givz56QVpkLGjOcH1lJyxc0IXY0jnm1ZGqopr9DkIYtoCcOEcMESdlo/PCx
SMX03fCs3YAGXk3wwUhndXpskWs/cfQ+mdkdOhPzWmx6zy98T7BrtMPU+3uEyshe
8Y7o6MP0ncJpr/nDkbqCA0uxdBne/JJWff+A0KtwaaBLN8e2F79hRofzegoxtenT
lT+KdfUaqPrrG+FbV+Yay9DXR+U2K+vZ2htm3wQjRYqe+7n+ih5C7+Yw75xTYSfg
B1uLXWpouOAU7icB516p+ml1NrqOaINmSqaknYWs6Al0LDq2GOXvBUUbmsNLPkY3
yEDErHZNToMFMIPi/Ny4gwUqPn1joC/E6kkNuHoe5fnOSzeR+GfzxY/FvvapzWyb
2f9xCaabgR23MkPufcLo/9MZIMQkSbzj7wi8c2ItDvNQb0X18qTGLwKaCV9g1ZpU
r8Yr9zmIOGth8eUZbTsNffILXrCAu9F0pUjIE2ATMuqhisGnbd/H0zTA+mi8XdbW
eNny2f8urhEk255t8g5Dr2gVUxw+9AcA9hFXBbp+t/L1BAfrGizmDrJ0Qxh5VZca
aG29QuAYYBshkgSJhdOP6InU8D35MyN8z1FrnfNTfWlN8Aj59YKiJhXQ3jT/lr0r
M18/TUmkAN6kT9fnycGTHnMc9uZyUT1urOTH6/VbirAxrScF2wJqBODtCjDK18nU
qVid5kKArIpOqlJwAUo3TRkWpRUjWZJ2kNxKCQFkrBZANjZq+LxuxY+luX5mSPaA
XxK3H3yDXfMOtvooBPT81nWfjWAeIsQbtH1OWMXlDqg1twTbmw1ySDVTTzfWtae3
4jCdJPGgVfQ2B67WR7hnDm18tanLsJWt1eJjIHFkboZ3WhGE2Z3lK3aEMlX5Lvtw
xoVujtvbYMyN+YeW2CoTY+n22ro10lyYiqwutTnespbKmwlFTtLGCURWYFOBC3Tv
S96wmOF+L1eJym4luUSHc7ecWQ/eeVmpDWbkr/7pSMuq5U8EQ91pfVJuxkwLshBp
MuiM+I3AZSukevyTsDU401VwoRzRFUpIOyz0fEkEM30xEZNBV3V7kggT4JTE9mhD
GZD4lDWZ931I7ufThLqyMLM2Z6i5VfLU4hDjrEda2sLE5ev/v3i3V4IVzyHPIEbZ
8oTYvDyWAva1Xd9sGrfx5eNyTJvSFwHmQHpgJLqNcMN3O22ffT6u77LBYZ3ZAmdP
QocdgdpceeqjjWZxM6KEPmPNgIkVpWeGU1UcQL+/3vEuMkGLDtezq7k1guOybALN
vzvlH5LCsgZ3Ff5jJ25CQZKq/d3Mitnoj9aPW3zJRji3zdtjAC1SPZbbSveJKSOI
i/uHmkSpo8Pkgl2TX0h2CpRxXXyYtyVPRDz0GIRAuVeLhtVAZ1psfTYO74YIB2dX
1eC+l7a5ToSfA7uEgkgvEDclqROmly3c7lGRTdnAcAZG7iUcaT2kkEop94CEbReS
3EA8dZe25XHMXIDOCf7ekrBzIjvJ2JK7xbLDo6Y3R4AX2Gsm442EsitLRgrrvydz
GBo3YGwJUMWWQM6aJ01E7K1LuqN1y7rCjU+HmjYxVGXzX3FCYZWhT+9M9MNXvlbC
BH7y4aSxsNGkD595q4MlPAzdyzkWra+eNCyB56Z3e3fvM+p/TB9fPOXggAdmHWpV
rxOSYsq+5tDhHVJLMt1mQRt9RtBhOLq5JSgqfe1H+NcC+Z+u+kx7yPe/cABwW2l0
S+HZ3eF9JSCx1FRayWlsGqV4aRpnqgwSy6IBuw67OnbM8Rp52VBtzrTux12Ezs9Z
/h5cNBl7VNqfp0QdmoMYcLybrh3mrgUMQNoVRhG7j+PFVYU9S9Mz/tzmXuDllEG5
mO9zgJnlfIHeH2rTvm9x/AzH+IXs3AXLVYOy/6rmf3a7Zj4DWPsHRwSS11J3kF3r
kPn/WP09nAjeSphGrjTka50tI0phqoUKbsAbRXcoPL0rrztOPjw8aT+l62bstd7H
D1635B4JfJ1lIQnTcHO1sZyvCJIBLf9V0kl3TtCM0+J8C6DMGxTCvlQKxeVx89qY
4P7TupWFTRolyNTq/hfn5VhA180eH51ydiUdhWd+/R87ijuuq3kDfOgov7yBinik
PDaybQGbavSu9XQfPSU/3AmvFgsu9aQkpRCC0mSo8Fzi+ZdXVycZermT55lFPwrl
TYp11B/jsprS9niLuZ5oiIJFNU6tSoXMgZvq4FsPVyP4YIB2XpcCgoxU+64uswXs
TBof9hX6P5VwJ57NPRaUso1kfHmr7bBaWahWVcl761NCWv3WbgUgMibkRwGqSyGd
ADO/PqvMop5qXaA6f6KIwpRGSvolUnwiMTbHpnxHL6R9GzYVfYusMdSpYH/XNvks
RhXP4QiNBENNWxieUDmwx1fGf5o/relk/KOOIZIZSHyIMrPG9eIB6OpuQneHkdTC
5yItYFxK4vzQUDPsQrJClwqM03JWYR5XZCCH7/QY7NibwRqZOOjp5y1izsJiKDra
bwJvyT03bnvrKbdw6LTHqRjsxLY8xNrmfBb63XYh+G6dV0uck6NCw3ONICxxzYgA
ttx5eJ3c2dfq1Rt005bQTYKG04FZWWgnN8BZhlWFrSUL3J0AInwSOM0LUoiWWl5l
5TSgTtBuZrupXUQITFr2E6QwLpiILrtMS45reqtiJGltdstjWduQ5J2Xs0e8uTML
2oVb5un0B0GyRyIVs1zElc5ASn5/TDerjOUFoZ+KzBWRdxgxnkWWZEcp1RsJpRip
rH7lsNdzewFZ+julubIvwsXlppI5Q7InO9bXreNz96fc5DHitrSRegRdSvEqY/Hp
0aBIU4PffDPeAv4COINYrgWDVdLntMzepR0N3oNXn+9PmTAQSwpsA59PS13nNx6L
7gDWe+vXmuPrT4XRiiW6dMVtLGagF2GoKNCed5NNP9m0qWFuosmfOFNQNKKkudJp
0G2S+L6k17oFjD/94eMN9lhdV2vq5F9Mf29gxusSeszxk0jMyNPWNluLFpwC1UrS
w048UDPBo4bf7ZylBlYQmcJ+RUBVkqKz0yNsDRPis9L3eBth0Gu/zkbhDZB5fPTo
tSEBhhjdDjVHGzquY2ei53v76iPeWFA0xO/77goVN5A05M/ykH4QDeMXaf6BgQxf
FQzjW8OYfufgcDhYk+qhQI9oj/I+zjdZyVgg1rYbPhGN26yXUXgfFwPHMnTxtUPU
rGlIpyUuTFAXz9NY9lALsh6Y03zqdzp0RyyXr+MGXBDK8bWXmphAgGVWIeDBGBls
1iV3ojiMlVay+YLGQqe21uHm/VRgNivTDaxvplDEXJqUTgMLNxdnuKJKtfG/eb80
ydrfXg+T5dYmJMBDu5i9C7v1NgHc+OjQnKsYyvIqaDDjzEj/LJBR5h7zWpfiMfDw
Z8PZtQUp/FgFgyjZCrsw6fHdGdrHHY0KScmQSftrkH0r3JaYAPEX8TncciQxU7dX
LMvr5Fp9CTHdbZdIutW99S6iWwNcJI/i4j68nctgIL7b1PKC+2/NOR5vdp59wtne
Ic+W5AwvC0XKkFrxMVezEM/02nFAaPbTKDg0RxOmpnKllfLgisNCy5n+Yu7iNUj6
f24aNL0EXcTUs1CUoQgAJmKleASnZk/53xikwI8SA9QrGfRy9XKt41I5waW2N8PQ
2ceishdPmQv6YTkV4uoKZeE9H+UGSWJ7eelZA9b/EI6cx/iARgseA2oXerlJHfRv
4zS+doqOGx5ot+VIcRqVH19G8jhrvDCuhuWnCsQDo8r0jd7DF3I6FLyXVBfYgM1G
0DwqHX9fPA5vWHjSRz9rmAmsgsPnKH4dg8kzbaj8V0IfyX94FD7RpouyoQcQcX14
pNVqsEkom2ZF30zItEZAGvUpvcDXZPDEKvuRRLKnEvLUDiPYKWvfhKEQhd2dcg5J
/fLKO5/rbmZmgoQW40PPIkLWLDpawCEGKTynV5TANjiA5te3C2hyjZ5PYyXp6EiG
zhSne/gsfx+f0GgkHH6ZvLmD4S4agg+xjBNvbvsL434aps3U/W7wJyOJ+YWYjqrd
pFqOp78xK6ZrqD2zau97Bd/IxXvS16+J96XXc5ekBs70u+DAA2+wLXqF8AvdyKIr
kcYmdVV3poW3OhLeGlu06deEKv1iLqTtvAZRsdIPikJksYqAYf+i23pb2D9ouQBK
wifS1KdSMrH2p8fvaErev+6UM6MAkQ+yliCRj8WMgAoY47mhXXVZ0jb5R4iqUp8E
cXF3mckHtopYleGYurFpkdo5SvX6IqDvm+cGpOvMGS2M+YrebazZ3gKnMk50qWwc
FcqrsrNhebdgsK6wV0ueO4Rp2HVHPrRZPvoRbVH4MsbMXS4GagyR+yBwkVYE+Y6h
a+HiOwj7PI4O90yjiHglzV9W8A86kkT1Z6OaK3kh9BlJqYhRkAUIX1/0HDSF9w95
YJqsXjqPinxQynQ17/pcoLG7hX3iipYFY1XG9he9yJebjgeE83OqzODNHZqbrRzp
cgvmSc84CobrjqUt+IQTAN8JaKZT5NKHwUaiqfiqTacIUL3kA5aepCyz4YbpMOpq
OYNlKTdSoCjGWWVsKnMD1/j7sSIO9lwI0kh0H6pemw2obKkzWWziTkSQTaTfZ0Y+
YzEZTZFIo09xM/6KgfxZeqMxNlLmCnNuy8Rnxnc29XZczjIm8MCdxjZgRslEN5Pg
HOSg4Eh/kyyHodqnRmwAjUxwdHaBhX/4Aiit5bKf8uGY6Bl697P0gJ3RGT8i7gqD
QmyTp4Nd9GKCv6dyyD6lI0WNLTLuXcXL9fB0VN3A15r6gjS6rMrB9Wg8DRpYayng
uD5mPpgNfcOpXUf1ktU0Ex77XLJML+Bzib7WPIMiuE/awyn6DHxWGpGTy6knyXx3
K8u5ebkEdwpZl0vboCEYGbTKKRf9GJ+2oXWfCDxsyaRgSF1xApFByoV65y9wjb4q
NdSWWbbyhy67FoLBYidLBM78hOZL204EJtg2oxOU2bGox1HmJPiq9ZvplroMLohy
SL5fZsrWuzYLL5jo8k5a3A1YUjG54XEmPOWCyU/va9EnX8lPI9H0PT6KXrrImvf7
vQYCTfgUayz5bgMVS0DH+bUeqFHriOxhRREhb5XEpWp0oLxzAlaUes312YsCO+Jh
CJhohS4F9vjdaVKYC8eDgWVSrhSVj2kqbns19CZpqxApiNdyyKkw9N44eChvOYjl
nTgqsepNg7j5zByz/Lnl3Iijk0MNLXJe6Np4KdB1sdcEhRUbpuAb8vScxMftP8ir
m4VQP2iWcoDKsh7xuP4rfweM3oqHLvNyMFk9h7S/oD43al/DD5y2Gc81I4t6AP5p
atTrFkroXWbUs8WQoFxcz45Gits4LvZUPyS6ygvrhJQYAsdySdBRCe2bzc+EawrS
`protect END_PROTECTED
