`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ev7rkaR6ev25VcdHvJJGIErLbZ+HytcdRNKhwWBXtEIcLYCOuRgU1DkwoLMpI01B
T0ySHDTMA1m8Hx0p4sepEBxSj2JmQrqYWo+MwOs6bv4gu3DdDnODqzcZn8g1T85d
xmO8wR6JNqMt1KYDayrlg71TcjucHwHrXo8mTNUvZQgT8tQ5WKK1Uq55GUDjisqk
ZSHfxTMkd7juJA6yxVBqOY+bFAQckyqs8GNxkDG5lHDDocMysKIbCbHRvz4xrkFq
R2e3jW4t6BWBPZwYpmn6srIOHhFzW9wg4F6QMjjdjECbDyd1CYwgpNZrwD04bDyW
LlfkZDpaRotU6L7ppLIpbQCjkp2gCMeInlMx88N8XTHY+ktanQ/qkJ1XNL0UxmYS
wb5SHiXSZCPawz6ctk4TtQTQXbgJAltPXcSplyMAfnTx+C/nyNlbTOSioXkLmwln
nf10pZWFRrgdHS8/zpUyLehGNXul75O5lQ4tg5kSMSrWMO7BdbPHdauIdMqGiK3t
O6suLgWwAC4jwTVidUj9gXk/wKPiTgLpXNsfGfg+HNY5xEyUdCGa7jSfjDueTUrb
4L/21FcFjDmVk74mDF0iWnZ4zhau1Xf6E/A47HLDXVvxnwYYgqtD37RmWEJ7TdMS
FFLrG+2oPD4EGg5qS/eKPA==
`protect END_PROTECTED
