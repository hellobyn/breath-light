`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFMr35U7Bztz1YQdeNeBoChyBN4NI6z/aSl7qsumy4veN5Lul4iSV2pv471Zaki8
w6rhF3VYRRsgdt4+BOeMFjtgFiN3wSEB8pNZ08WgDG8A1Y7/fo7WU/GEFteQl0t3
yob4CYLkMH+CFZFLiHFqxU8wMt4n+AljdXrPs5CUyi2ZL4PUDcdlT33kuLJLJa8b
6AyTsgXKB4rxwTBK/Qo0wziuayJeIE/iwLEpne0VsK6FWUdbp/k47FemZYAjU90C
gEY3SSzsz+DpY72n9no2lypSgiKW6CtsOhvDXLegCgeEiKHa1b/SuRje46lLus3G
RI43DEalYxPiDzdl6i1s0nlc08XcVzmEZz5cJ1Jk0qWblPqzORYHy+zOEVqtdgJY
paIia8g8k94HlGRy73/7G+mEoBCVE1Dq2qJfVWk6IajQ4YqrfbcKodORCrEkVxXe
Zd+RW3xD30FuIJPW5sHwvKzpdHdx7nBCe34MlqJ4G8GVp0TOf6bvwAK/AgTuIoe+
C17nR/LsFx5SJRuELmzaDdTSh8TqMAeKAyxZAwXmQnQItWPbHMSHOk50izGA4ErN
c3kE5DzBTG71TUUV1lPtGlNpHFBdlL1he9rHVbzyWEr9CrLJpL5rhkBcrgAQ3dYI
g6cUbDAJ9rsFA6tRAabt+dh87585p4z/l/8AzJEIi39DWWQ/n+ygdnb3aLGwnsKe
6dEyuVEIFXI/FrQKxVDNCtrXG3Rx272JpViVYLN8gwU+kQd4h4vNkjGN+UQlFY3e
9Kt55cMiRwH16nDUu7e7232triFXqUJzKQRSL/7FfSPhKdmZua4Kd+AOVapxfnqh
jfuoHGnfG/0vD4o1ckMeoT66dS+cHdc8srN4gn9HjTPGlFK6KyWr7uYkkaBnkrqV
NtQRFexggKe78zAGbRu1+nkOrOAP5A3R3sveN1EFMJGLZOqIvTZGO3upfX/cmpR6
QfS4kP9BlqPiV7TDhRTBtwArECqYN8UPUyZD4ewoWklXWrqKlTR3xoGM8l1y5Zd6
lTL5RFylLwuk/HDSuJTRHPjHcO9hoMGc4Xynp25TypeM1gI0XILtD8cED85UEiMQ
NheiRIhvr0D3RCerpF+ApwWhWnlCerdNB39TPrPEBxwhFXoNrTH9EjTEC1/E+anH
2W+Ux2dVI8a5oUz9HAD+rTttO8YBHEmeJPjam6wPjQcnFBC5RZBdIaBcc0GAQOCL
MCrlYxtJvD3cDQWOsFA793DlZcwRmxa4ecYlw7OYDUcNpqS8Orz75LfBpUJN7xAA
BB1MqE5C4B6cRySUEu91NP/Tn2MeY5ekhLAo3ju93dxhruzwEshsyfLFTu5PBu6N
NSDLNPAgo3UtIvW65MGtuZIbKbQvKbLpLTSKZF4Ctyd0VgGF+XznxIBcHEQGZZKS
FNGEA8G07rblJy9K1BbVwAktEM+TLVA5jIT/2/NYSrRLqF/IUubVtoONLt+pYg5X
PJ9vSrQICNo6snqkj9nVLGbkPLOO/FAaF1sPmJNKwPz7TdNFGxN8ywz8xobecYh2
b7RP6cV+4L/UEVPJfuBPiUCSMQD0DPWLdxKS+TlewPQLG02RoH0f7ScXnfYd/esc
44S9gJwP1FBoQdG8cGx1HCcvvX7qH9wLOu5CtiijhDr66GinRi8aNiYh7MWpJGZh
Hs+asmefbhuzG/ErUcFMxwoAHy80VObiBngTsrVUaOJGj1g732p2qMDwr6DF5Rl7
MwdbY4wjSSPBW7EnsocAyWJeGT050yqT4hWIgXpDA6r8ynoDNqEAWspGAwfNUFnD
0KXI91vF6H/CII5PlBnJyLX0ekW3OYxEDZlvoj3gOInIoC2+Cwr49mIzCL1HHsMJ
lhf2Q7boGVMh8WiU2Lgz1IkSiIYEw4id2vwE/dByUCvf3iuofF89xIg0db9j8zEd
4IBqFldTbBFD6Tden4AgG57eHt8UY0+FcOjl1NF842hz5tEAAS1DHqI3jM3yoi1b
byIi1OpKV0FSuOacbUiZlR87313/O7HlpanDXdlFFqYIbY4PYTln8XJaCFeWJKC4
a/qyN3zS/t+u0E4Rii5jXQg8u6wlTN7z+DvvrBGPZbLHxw9E6qFkGmF2yFn5U2o7
XbQLCX+9MEeq+BQweQ4AdKBpMsp1e86NZlAl3pi4pqkLmV6KX6L7Sgr1DWBolGNr
xyZ/rSFwajExi3//P4FggZCNWCprS7ToXbIXiZIrUicCtVPGhpiN8hIL+JXItaxi
THKO+xHSEgk0IwYRle7bmb5EZRuLmU8sBN0xwiVVheEmwzjkjHWXmDHd5nieC8nf
sKk7I6TLAO4OZNXiHdvEfxDqu+Xxua8onVhUGCUlIk2ejXoe8AijDmOYTFAvOYPA
oEX4bkNHF81gE1TE991C2x0nlQlu5Q6fISZpoHzaCdQYeykM75EkJ1UYSpcQg1BB
8F/CVSyuRJZ/I+lju1qVQAR6Jf7xpXscT+/jkBww6lRjAjXCoj5IcYnDi4KRpjZh
hJmGhsiRgzJjm+jhXx9ealND2qGYYhM4doo/9I3Tf4PtiEbM/KRc5enT/ORIQRZm
4BQwZViFgfrIPse3V9D8a+B6WIljwMvvdChhrxFzdW7qPwKWjiMeEo8ZQIxhEF0W
jiF5BPpl7B83ggTRojoJilQdDQAQR1+tf0raeMMVCnHyytc9f4JY8YQrI+vrOmAd
+XpLIbGLn+ZJVZf61NidUEetW2m2JSxYlaJvHaP4ErRDkJpehwzdo3GJiSCopvp5
zQ3SJ1Lzvqh8D5LdO6xdJKUuCxe6uBIE2AjQDi60rka6y/K+nIrXARWlSYEi5/za
RiKIbWhE7nUDSw/rDeCPsOWvMkKah7ctLckoldLp+bjp7RHNoqzUvud5l4xZio5L
x1i+jAl06PKzlvWlGcPeilZk3HIGEph9UnI0odnXguNxl60coSNsP7sV2HC8Sc3n
fUxHvkN1B4t2lR0+sQqJvra6ElLvZ7Sxp2w1cZNtLHykwKOobO6pyBR26nF8sLG7
W6eaqgZGQdizsYOSNupYpybnWQt4h7jmV19njthawGndsZ/cNcgvr4eArjg9KJ+G
VCz4EXna9xnZ1Ed7XV3zv4Yl8at6SVavL4aMX11XK36tN1XVgpM/agsVd9xh6OPX
1X7LH+vsKIeZGopKnqqtm31oEkdF6TnlYZTAXkmmIsIWpm8GE8//GBMUzzqZOFcH
5NIguhJVXhtunhVBmy2dNrtGyPFJzCzK+1brbhHA8K/X7U0i6g1vpJaL4zlee5J1
2b0y9CmYhqDDKRQQOG9fc7YCB4XawNm/5QYgMkZU4XIYWFEnnK/lTcssmSUzOlY9
GmaTTXbCd+x5vdI4UeU1/84Sij1kCbhK+7Ypb8Do9v7lkdymNWJXphJvcS4DULuW
7ZsfkXEKgMtskiW6rzWZgPDLl1mRkYnwyw5ORc1KgI5jOVfmTdOs58NIL81zq7OZ
jjSdPfC3A5838dPLa+vhXXInbT3QqMLSimYdLAlNJ4McjRrbZiovbyLDB3uwj6T7
BWuSom8zXOXjVTFJZbnCifBo8ssZavAM7z49fEpNmAArxO2HiGAliRU4UsGcoa7j
VrHlxon6lmuwV4bTQ8ahPyZEMZaQRix5HPVFUimg/tlf/QVHO4R/hKqEOBskV3T3
O+cYBxa19cd2SF7gjXwCwPjBauZyzZbWwfbEFmQq9UoFZcNCbcbQHIYAl6psSIhv
3LyU2s2aV2ajXPz4nFws+CUnGGaipgfA5anR8k6ks51d7M2IAEZu++RgfO7pKlF+
q7Fh/OupaILuw9A9+dtEaPEVIbJBob5ZEmOK1vHoocZsFoB5RynBh12dRwzQ5jOC
gdAy8Ifbk1+95jt/Aio49jowoBnoo0q6cvyS2EuMR289uIeGL9u5X0OJ7KCpXhVH
1iQy6FRYaXKbfQe1t+L8zf1Nr13jYESs8uRJiFCnFGpq7hegE0LhMQSxPw3IXMT+
YbE6G94gv/5RFlSEbkcDVuwaVBdByI5199OpczFb8wyM57kX6uS23RskchlY6oeB
XnuHO/wGKl+rGPFYQYrpZI7JYldB2rslz2atPXTG7jfH+bpy5G4Bk3cPvBf1OkMk
NyDiAuJjXTrDt5QxaKVdzzZBIPSFy+4VTB0s25n/6oaGSRHc/sosEoVBmvQ5ZdcA
84shJ36kKb4EDTByxD8estDTZpK6+zYEV7+CayOxdxFYxnizxCOaL3lnEnRD3vMW
9RJvN4jc6BP34uf23zHdCtBBnjU7xT7NruqGC+VsHdD8/bxMiBHOqg/Ho8CNPdM3
7V4ldfyXjp0aSoAkomFx9oA/MX9AEiWSQFN9sq1P2wVRSxlBbDujKflYnmQaRhow
u/uNdw1ZZAW5Mue/a+KJSsZnzcq7iBwy/e/5OVNCCkgJ4jHIJHe9DI3Oen6TW6ZN
TRd/6IQIbTOCtAcN1DTu8iX5L3Pfe+PrV0cqcWofrLBOlt9AtsZUM3ixz7BEPFFQ
AAtnrBet4a9B9YFc0wb39zZE3NA/10lpA6rXgLspLh8dXsgA9r44pkA/SRqnyVqh
/ifXhWNwmZX3J7Gxn5CPfWjVlvUm/qtt8oZ5fFJIkxO4HduTevAEGvdIUVbnBybZ
33visVU+DNjRf3V+gb3caw1sIpH3lXvu0LkSDPT7ely8P3/8G6N2VG/PLM713Rbg
qfoY6KR2oG9Ln9jaA5fYFbNfrMRjsXdTNad0xC53mtC3CTAhgZMFmhwVT5T/OIYW
xv7sgrozfI+VtPsedJS7hMDFz3mCK/7LNGUpIkHM/OKlYQ6OwMejziAsnXQjQUTb
9RcwEph0VK3GGMNG+eg3C6/rp30y7h/3hJgBpcOAAsWAMSUZdZl4syv9tqAIN31X
M5fKii2BGQKVJvGYJzuHTjoZ8Zfx0TXSrCyu6SqpZR2jcOHAQ25FYOtcbNicC7T2
9ChEFkEjXwaCkhJ0BhWvB0/0fgLY3NlJeIFduSdMKTwjXzjA1DdZlJ5+gfDxdmtY
m8434l8m2IdcU06ZO05f/SdI8ERhxZsH+ObSdtmFxzvN9z88SktKQ+yPGT68CPbH
GPDVj1XdJNxsBx7PKG0843iJRV68AXYUl9RywyXMWuZBhfP04pKAS4e0/Ln5rlIs
C52lKVtPGG/5BXrdPw1gfDfFBB+OGwBrp5MAOr45OrWhee+kzzkk4jI/b7M9PHUK
mDLPoOqbePemgdFaU2Ct7gHhoLfLHX3F+Ge6VmOfkRtaE71RaRi9dGjv/nUhwT8G
Xdi4WyUyCj/CIQzAWMH0aUsJXmsAJ+dLKMiy2XyEDSJG0zSzWMLelgRqbKxHrb8z
h8qGvrToHiJZJeTLkQL8NLJrUcuQv8cVXp5BpnSf87MXBCfj5gR9f95V6Eqyu5cF
QcH5D38F4hhvBSQPYv5W9xP+g2+eiKKksJ+FH5DH88LhPEvjRJjX4gFSO0IknFbM
eh5NHcv9ZFdIvlNJA0TQCydKq/UmFW/UHJT7Zm0yWTAa9Ua3kp0+dXA4MylPD9AB
aksO8o484FvXwurjhsNba+2bv1w+lXy5arvEL04m5FlagIQVESaCm51/LVhSGi4q
LsEIRFzv4VeZmJF0/Snc/so9UYNxmoGxZOvEP4sO2nLtkiKmWoe32dW6MObrCPo6
9ofXR2DVdDLA6LWgVyxU7FiiOFKuKQR8DKwjM1bFhoawMGBbX1v+5eI9tvlN9iv/
sDMNrq5W1ytwZo29loHtluJLZ3ObMEqs9Wl13uF2C0HtisY8WgyzFu+IADtrehgJ
1JOaJV4QRCpruB2Z5F6dLcBPds94oXRuqEiWNpcBfESTe/JmCUfrC59WDuRpQ7Z1
3qxdccPxySl5unetT9vRjQn8rPy8+mw7oBivGV75kqLXAZlhOvbxVteqojPsxw96
HuOBShf/cl1Dq0rWj4cnsf0tpqtFiS2PE460fX7A+27qQon5IZMaKcib6KMHWK+t
OpCj1CswxLCMPIDf2v4mYfRruTBV0squhgvCE8k84SVt8Eq7QvS2HYcn55mkVuno
dYGUfYj6hJvR0YZkMTOjwJruIEBEt3gF7Zlh/+kE2vBwvFV6hWgl8AMy7cN1htv7
bZccuXFVAqnllhcKhTAKZEawNsHaTkg4tysZil7QyUbC8RviFatb7EMroDkuB4LC
F8wvYaiob4qEbUhsSIf7vTTqeyxj696j3fMLwiUymSTFF8vMDElBSBeT5KQFf9CL
bDIc8RdbM9T0xGSqTFrbUYjHXDuuYq8pmCvv29iZ5CLilzJDGlrQZ9agYHrSCFaf
S0tGSV+98D9VrAugfpkwZCLmAtbyZZ0KHIAv5PmCIvFAdMj4cgC/SXotvMVN/OvG
LNjwkRlOZwpK6AuFxOH/Ng==
`protect END_PROTECTED
