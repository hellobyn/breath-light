`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UK//HL8etuYkvylieFpFDOBbojiLiSEq4UnANEDM217OsbOJWsTWGBGr8QSE2Y1j
z831dL5LXpzocd+OBh0uoZJLuR+2n/cDm8+44Vj/t6NFQJ1gW7UqpROLZFWl1YFO
cTcPnwihYcRWBZPsTw3/7REt6NMTiqFiGmdIyqV3aLiPeB22XaeI/GbPm5e+TF6J
Ogd9M+Og3ASp3PE3gAA//ny7sme7YEWJi/6Hb2WTjrO96b8h0pTolda4RSb+3k69
SKJqI0Fn5IJfJ0NYomzWD/yLQp3fP9iXZi7Oa1Q71qHPP3ekhagTe/Ht9wR55VZa
n/2xVk/nbBMmnDJOIbjJv/Ifl+SvQHuFyHl/1SukXsQ5XoCRbVwElsn94mIjb+Mr
HGahVfW/HwoTJQd0sdcvsrvYv7Qz8SCA+iZr2rh5jrS6xNdnMrTgGcoSku701elK
j92mcEa5paE58ryLMvevUjxVsxqLujV8cNmqs2+6+LdRmfob3b00+YTSjH/DVSE/
yE1IDr85S3r9PmuWpS3uc91gMEVtRfJQKiu+HJRQsNQ+ozWQMyzl6zFPe7oQF23F
j5N+glHX2dk8k30puPkDXS8iw9p7k/Alk2e1vyYK4N0i2ciJeljAlMXIDBRUV3I3
z2RzhJSy1IDQnlpye4rHcry1+YFeBpHG09Oz+UmhnKyGwl5coaFXrPbIQuiKty+m
F845zcpS9aA6hTGGaWT0jaNP4lt1MeSbESX3lz90mMs7zw40PhEME9rc/sXwJWe5
yBR3jfmp4oEMVeILcOAeeuF5nRzlCkSw7oZDANmlpIueWzofcNkOgqqp8wXg9is5
94DElBm2+dsngWJQjU55ibtQh0K8GPyMmCKWzWkGBCWe3syALaz5EsfuH1/5WE7F
0ORHvraTTbThupdXxMZPVmTOSAmBA6vjh45cbpX/T53RBZHEjMeowrZIt7jmccVr
T6JvEn+2BvjJIirS6SKSjVS3fbmYjNvRWa2FWFYlFZ/n+hAaVIv5uM6H0ev5rC2t
/ZmIIGYCNaUPCZURJN9Q5Vry2YwvKLKiF46pzoWf2NA=
`protect END_PROTECTED
