`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZCUJCE+axlVAe2U+po6zrzKg0XpFP/mBNtPeKizr6B9ltScA0b9UhtLvyteVKPn
caA6Qsp3U3/iRKqUNmWcwjdk+GFFz9Evl68oGooDGUi7VGNlTuxXngyPUOmqQGrp
h6Ke010KC9A6wx4ynchZcQsZzyfhN7iaQAN7j+/OFUcfJ3Xvr9S+MpDG8L6Dpfd1
pKczrePNE3oHcO/oIxihOp45wTZ5Qx5e2glm/os0cdWTQboAVVrKnks2Bl/hxOZ4
4fqc3BNxrSvIWExae5xOm4Ro7KM0FLSC5JLDhqcVa3vbwWhthDnMiOvAZ60aKKOE
/+QGgcszs2h6LlpGSpJuRNzieui6MwC6iCV5yM6JcS6A7AMSrdits4fA1ZGuF6Kp
QV/udE288h5j8pRe++IhEHaVD+yOCrVnikKDeSd7cwawsnQ44LXr9ELn5Io3ryZb
Ty6XijWYgpZxrDv7pECNJr4HbG/iNnRJC1IVg3iScAUlRbsbcxVd2KRIT2lbYxiK
bqDLpnAPPaodxV6MPPndSpXAQIkufL0GzJcn4WE5mvJsWlH0ghf1m/zAQWUll7EH
H6I8sM9WAUY5C+Pr+txu+sD5Ij4gjrh0iQVkAM1SfXenlVZxg6O10iAuLjc3WEI4
VmGlpndizLBs8TEN9nkGE1iaIkmNm1SbVn6E91QA4U9As+yww1k88+Ht25pKBcVW
cJum9bOqa4U2mX5278hu2UDjaJqx8YDNLpat3drsM/xNshKI8kIfvAJJ4S9WG+yS
ECIhps3h1cu1Efuk0DoGH8Df4vmDSY/LWgWc5JSE60AFcWap9bWKFVBJJ5pOqymo
iukBlSuMHxDjSa8psoYugvg44Bst49v1yoLQXF8fo70+RoKMibNH+a59zWmHs0Y2
3EVJqij0mRd01yD4qj0LMNWLHwLTfqBS3gZsIqqPrbQV3RykEHfNDTuaSYh/D8um
nMHCQ8yz8xW35g4lGS+PrlsymiIWBYfjizYRDF5p2h/vPlAVqw9f3CPwKNJlqpAD
2EMk9KpL21mnqZ6jhVd48EKaXcTmDlk5Bc+rCEHwYs0Y22ZTvo0+dz9T0PpGhziN
JdOYunoH9W8MHmxVUEEm154Ckioq+CwsJAVfjxYoW7ceQMaIiOP/oy7tJ5GQXSNc
9eZcHgA8h5iisM61C505Y2P+mKbcYa5Lkj0jsP75heYJiGEtcOGl/dzeZQ4tXuWu
GymQWOaMkDEuD2dYWUFLcC5Bjt/jOpBAT68qYv6JuJInylvVRJ2nBWkaYXyCEQ6O
G7Gqfek6VYjHmYb1qsPn0CVkHEF1lM+kqmdRKbWf4IyvG3AhsTg1KA9dJgkxkYEr
+aO8MXwdI7ujkYPEv7Cv/+BeJeHhkOxYSKzP1TRdINMnwpE+kh2ZtLNcRpsjl8rj
TshOKE/EI53UYDkfLL+aehJSqwegAwVqTrYBB3zIFRHqvcGpS5P/i04HTdVT9AaR
mRGTpS1hEUaTPDMR1h1X/d9MViUqOXyVFeaGkF6OC6BpUUianho8XG1L/si1BNDl
mCEb9M1AFlwzt7XI4Y6AWVySa6/twyWSdxaHc/rcI3p1LklO1AwB++GupobZBCGH
e/759/cQzypzbf/sj9YS/tL3rUiTGrnT1Po7UADPakKYm3rWLh9OtuqIix9gx2Ef
z3/e/75fJ6vOmQRIOxgQyz5YJeKJTh+cIE7PjAQCeRmLje/bch+Tcg8rwlzVSw9O
RDjlCNXfwXlI7Cz5TpfErXUTj8+lAeoRq2GkPUVMNqZ+sRcC3vH1rNF8VUfz+ppe
pBE1LwHmOkQuQG43a71I4HoM8rqkYQsAFirpn7iu+jTkEOoAn/UPJALMdOrBNy2Z
8yGJUu7UhopJoWv6trCjR1zcn7ELWEa5QjKQHAc5041le01qebgsM99u+qSTNbMb
kfepgYHxCsUCicEiGMe2d1n0HvAHfowaU4j0CkV10rdZqRHW1igC/94e1qRGwZ4e
hR6VIxo1PUJlFAsSDqb1/YA21GWXaPfeTf47v0+yFfHeP071+FiO1Zim/SbpNpEb
YpznWPq02g/mJwv4PsyLKfosTA26ER92D1tKTzyFEp9AgWK2qPqxPtICpuUMsUHu
71f17QMn23nXcorHd/jsENWjsmCb8syMvJ4EMYJZX6vI5fXj41uhSlRx7I3wUpN/
Vc1pstE7advTMv/+VyMToakItiZ+5O9I3VIP0dQVx7fgx7JvQyPEd1l4FbDnj3t7
6feQVo9T7qxkhfmc5Yu3QhUwYy2JZWHIICD9Uik/RivXq7RACzcJIAFss87ROHwq
jDPJYlO465RL3MuFdpCtUxsLfXAUQuPQvq1toEAg+Zr9QDLWLjrkvzOMFPu3we/c
Z8kZoVbM9QQQYvmOm9HRP67TYWuj7HCKh2+C48xfeWw7JlkWtaQIAhP8GglCcA62
Qs1O6+KuNAUatAmboRFnjFk8MZahB3jQvcWi0Ca+IcveFYmN+Pf1QBkswLD0M9kg
a+po7BPRZrZK7jf0v2aC2qpbjtVS+TVkZK+DkSBLpomXlfFnc06TlHmpI0u5m28D
dr0vHSyABLnnG9fBzOyT+dWtyLlFVXZxEJjbPVx+3R/3DpnqxW9vLD9K0Y8oSheD
krtxyrH+aw63bNeYcnlrnwublBi7J5V9AMybsBYdqLipm0zi9CZWJJX5bmDjOpr7
p9q2WlrT263SN3mfmVBnHlaMLS2piiNT07O17vdwKu9SZZnc+of2zr7vTbvqjtnQ
+1FgwtH7kacgAE3E9eaAvt4ywKtiZlT61c0RVrvuhtHObvUitx/ZfdWsyQUzlJrR
uV8kSQCizqUQk9zu0gahFAwsgS524EaJDPnD8E9XyXyDqp0I1KDinit2WB16W/H2
WeiYuYOrTifLNjh16mzn4Ep7Kcp3G38HsjuoGHC5Hn1gEU5/NAUBsmvGeirHnq18
deoprMLdfMwSrEz2kcQTR+95iEL3DajOQ8RFCBEjTMyhjMD/Cn6pV7zw3oZLc3bs
`protect END_PROTECTED
