`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ujon4InQX+tixQpLjDAHO6+6hj0l5Wt2BXiTk/9Bp+AN2ebHcdzhyENOGqNUXefT
2MtBJjo3G4xtQPJszeFB9VLABse4HK/9mRyMrlI5h86xMQPaugEGBbM1PnVY8Zg/
IgT8KEIGbOShJWxxxNUJJH2/GQkQeYGyWfrkZfWHYv9k8yF0yQZmt+rky+vObzeJ
tVMi3GTfq98cMEDKZc2D+D3gmUVYbsvMQNDdJqvVqY8kg8ub3/DyHeJNtdVqqahK
37KqP9Q436dACxM5RyJtEu1sCMhh8TK4tv7/nbv5vm1xUSNVs0LpRVdP/LSRefbd
5JU7bezJqTHmywabzvVa0AcyENTbGX4yKJrVT0EdID91BlDm0LQYpp3gECeZFqqs
je4+3/qN+YfmfCg/VvZ038GCuPmw9tNV+huL/U4ntV4Fw1paUMkoV7UR/kk/3sZu
8pATkHqKUzjlCDfQb3Tz8PrF5MQb25tt+reRuDEINyVx2yBXxWlqb6tPxToF2v3g
Xh4i+V3c/N6avtlcNjUQRj09ZFxzANboYAZ+uJkn3DJCqhpODIOBiRhdXwK0lHLD
8xKd9oDr6BxL9ZWFzB1fkzcWUIS8/f7+DEmyDDGNvf2MyKYkw1++pvCrwMgbEfx4
df5NuiDKn/PvEne9H9E6O1RRfrnmPHu5fakmTHMQOHriUOpgPkIO02BpdUtQgS+Z
h+Ox2RI+K59k8Y97/9QYRfmVrPCA5wU3k/bSjJf18Czjv+5WsHSUaVRhv6hipAod
zOE8Zgz6WlYCyhOCudm9zzYpyLWqufSq3L26jd998VZjMJDvq40FO0HCPgG4WO18
Igwz8dQVcGXg/QjjuJNEaldb/js55E04CoxuuKTbVoIJvMjldd2uFY4Mt0Mlj6tl
EYvp7si4IIs4FzY9Y552P5M+pocjMd400tJj7eVYzPHkTbVhZli/QsxYYDCXe2Qo
4XC1eNpdKUZgqSgIPWoBdeZiXirWxE+zMNah39UEPmn3dlPBDvqW+bHRKZOGkpJ2
2xpsH/MtXx+2M5ZVvQVie7V2HPENofSqvTORiPUKBYQOzId6gvRTReJvU2a7GuSN
kOVF35CRoIbwmL9f889ejvRy33ThoGMCQuIuNl6O5gA0QnQGnwPg1Y4NzQzUSuq5
wD/XJtSrekL8ptTqb79CLd3JRI2him2HZEnWaCG1ZH2OsJ861u8AeUn7rCRRt2X8
GqDeSkNTDNuXcNroVYaKcv2fetl04HrjUMgI+SwQBKZFs8DM2M4dEibxmKoNWI9v
ElCHjCR+ZQRxMfSyD19uDVYu0da7EdMBtnN93WTGteRiK0lPAqGoQUlBS10rL1Kr
/lsVYaEPyxmvzC6LqRwcLTvBxAk0GXnNctuDlBFbNqka6AVjLbkjDCMTU8oQ/s2/
Nbn/h2OLF3NOyhiBndJVTzg743mIkQLQloi/ztSddF5lIjZfbP8SRdnP/zOr2Yxf
oM7EZzD1/C6+jf91aKUSL4zFPPrHocDRFEabBl8gVEUlEf8Um7jTF/qtCueSiXHf
TASXVWNgAIgfG+Wz2qrf8igCcvN1Jj1EsLjDHdt/86+/RDUYI36Ad2nPS6zksuUc
pqK/WgBOzFtSd98G8jdmRla0f1Q8c5tDrzp/xqqryyebqugJpZzdJ1BxoCURqHMU
eyk7OgUe3d7CxQE39QBF4yij2/1KSJF8tPIXHF3ecL0uV1fkndAaCAtfyII14BgQ
6C9oOlsdns0Gy3sR6zNie7XqScqqQ4Y66uGLG4oKBo4UgBo+iMqpA41oMXxwfq6s
e4IhkKkw+rJ4XQzAOY/i1SFg5HpzW0vSyRQ2MPykm7JyHppMl6mVpvuXW2yyKNB6
9Ut/Bx8et8Ybsa80d+mhk9doxVGLi6anffNzAH6Ryiuz2/cVpxmn1uj0ErVo4pt0
KDHKt/nP4QmYo6Tlv7paaGQanyKnUfnVG1mcbms9SgS3ke6df/0OcRvAXjHdrxYO
++2uzlF81DDQsVDzWMXWUOvHQ9O9MH83TFTg+yuXLhJjFLolNJA/lDBaRx34a8Pw
lbpEK6xX0o+kllwmyQHU/XXNcal4CucfDl6RM76TXI4AE2E//29VziDNwQSOA7up
Nfoq4zmW3S6HD2IYrbF13K1GFc+V0Eufg1qZe1x9i6pd23qcPYnzll6LE8pX7qgh
a8c4g4toAn09xzWDXwnMJ4tDb62/LL3UjbUKgddyeNDdpFn98m+encQ2acAWCg8b
8GdVz3Minb74KfhRXDrpn4CxNp6rlGpuvYlQfX+HoB3M9CI+T2mctcnXyPFMJOfH
xLnGE/rDt6vtiwmQq0phtY77aQVYlTyMKAzzr1s5sLyxtidJabiThcUiP4yMdaBz
j6Dgnnc1sYA93dcvy9v3LLAese9UA/2V2ZXUzqnMdJ2hTbE/bva8kCNsh8yVqVaU
JaJYywuDLS0AAbiku/d1gw+JiCQZ2Ob1WOnICO7RZh0GNp8dwH2nD2XCcb4dMXGq
ZJeak8aPHO7gPk47IZWZkOSZR7FNt+YjhJSwDIaYNsf3w2sSECy/bAzbA0E39Grk
HYdA+52xti0++r8fH5bL/+pDVSRt+RAzXDIEWjNv1JtZMilr1EZyd6XkoYt2NweU
YZVi5rMtTA/yL/cUp6qCW6R/f6BkeKrq72QYo/OJljT6xgO0NXxYI3MXnJoQintM
plu70MRPJ4d3xf3gNGGaKwbbZ2eMlQV/bYCPxBYez9JYd9tcmHZpBz3S7IJ4HjVB
U/gWOx22mnmWWq8GfLPTJsart1a1/gWhAQAd1mX9I6YN938MveqE92rWOJ/y90r6
FOCpi+wep9hVOooOeA6STZ+rQAvQntogLsaKgmLAwzdo6jPYfVM34axoDb037w0e
1GgxYoSKberex6yf/inp8rXcgV1A9SqJ2p0rbpzyikbtnAZDzm5T9+Ko5qTdSGdO
Rk+6+bte7r3jipGsuiyUX/TysH+6hrfra/AAcmmOhWpukNUnmgZiNt8f03DNK0B8
K/8C+8qlPEGpgVPrz+7KRB0sfAmpz3IOFkbmxqOyxGpaEJXHQuCFMTayVy0rLiWo
0UUG+riX3T0obhvfNERJxOp8lcJ0W2QCEzfUBgILe+DJ5hRYLnZg3LtQTlUJQ3lL
m3uFUiY9cuwqM2QINlyzOcsIUER1cDTHLBnTpGOxHKdEU7/OiutOAHeenNgCEJ9n
V35ETZsMGoLfIqf3+JYGgg5Yy85xhlCKVf9XA9NZFR3bVnueKOrMj+gyjD2NKN5g
E86ouSjjbYpWQI5kMF/0KR4XDuFwnygftS47uE+vtOMbtiboTs2mZ9NrsCOE4pfj
/DjO7j+6dLBaHv856XHd4UA/Ay5M8y3LDy+wPKJ/7VCSGK0C8w6Em4FHtTU+J8rC
pDB0fxra7KpS5fqNZjR6fqzs5hpwgDorGpZW2gXdD8nwekxTQ9Jv5cBvkA2aR/1l
T+DrA0NWjYj0/7CSFBlYBAwyNBcDiifw2nfJVAE2ZW75nh8JDeJRy4O6S7EWTEJf
CnxqsqDAt+co5fNF9LcCaY5SGyJBgOWHuYbTRpWZnheSDqG8G+qyKYBixQop/G3G
kduWIRB7wol/HF2QjSZ7fCOGsxScBzSmP/t9Gk1/6p0ynn7pf7jWHjtxgdF32rwS
6uFTV26kyzUGdO3ndnCEYcWzndahIRYNv/tPLcWjRcEn2/UdyDQQdbb13x6zLIna
DL4GRuCwvoMJ++z7FxNyll9sK23RPsIMdb9yVlPLfxo4j5uubytD3uZBBAEKlAEx
GbAkFDuoxEGgqyn+ZDaN/3DPNdmsKFzGGlEl1fYskja5KfIFW+xlKPutPo9WL93C
+B4YfyYQclzaWS1wQn28eSpOi1NT7eW8jVeH0F1G8rcBbu4feg86m0hP3sYVJnb/
WIRtHx7PXT1xYeYfKiS3XV2PqoyF+s2NdRP154uJG5hvdVTOUg7B2gs9t9oZWrcn
yBoJNfuST2aIAHC03oPkOMD7KIX9eZxIBN6QDIZutpDnRGippBC+qIm7YtWct9I3
O2RD6+Bf7Mn/RxExen2bODZf4matXE5HG1Em901YMgGAp4VUWE3HGT9EUnlOBIUu
X2Z7IoHWHRbM8TtkAvp/eSJgf46NsLOuNoShg0N7FkxtcujkhYzL4ezh4AfoLVFV
zJtGLGtCZJYzOMOlUgk9qNsyKqCBQHGeUB4MtG+1e2BJwYN3+oOS1NNPuhudUD1V
FxmVGedAiLOPYWXV97tfIQ==
`protect END_PROTECTED
