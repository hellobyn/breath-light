`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXSXqQpmqnkwQ+Vm+2D6d9ZSKTUph9nxByrxs6ArsijpwzKq8BpoR/dabjgBz/zQ
HnnmO91YnYmD3fNlUGfp/beUzPc90AnTPJ58fN3TzsQW95muWvHoyL4rxN5ekERt
7r5LsjhanOABgfknY+GBxesrJYJGMFWUB965A4/jobFttULDyk3/hq1ycUi0VcGE
rxgu/cj7rfP3pvwZVATjCqBnsWxXY+bRXnJYiOkuCu+ZqnqhL8KHZvUEek6JCm+x
vJWlZ39sillEuGxm/bDtcBMvrAPYyqCWqgzmAnXG6aboBrdAPisLkIOMMmIEqT8V
DgH1dc74ckVWydPlqfuYfjHTPhXQ3IgcS57yjcZWLRUFmA3lkqWRKHl3EpCPJKsL
Ls6WMR05xIfSAaDokdzpDaXm1riMdXdtWdUemxMZgJxt1d2QDYTwVxKFDJCg0yjw
r4MRqL/Lv1FQqlE+P6u1C5u/AM5dFhh+vfsttOoxjZNerKiMxnNTM5N/TpXEEjkN
1Bem4bAzjWvznqZe+xcTHQhuCb+jjrjFm8apm/WYqKTe+Rrp2EuRcTIFZQ+799uq
uATJor3BNXKlFHD0R4504S+K0WDleOQ7q6RbJGS7m/70RDrklSUGgiKDOn5FSCai
YGTyrPSR9dU9Gr0Z+jtxcPqMHLaJtsbJw/79cQSyD8i05WCeSD8gGkk1QcKU3XSv
zbFzwMFSk6QQJcpH0oxz0psdeB+QDxbtAdLfd5bzeatfZ80GJAGwJ/s94mVwX9UP
HndghYJ6jI64XCyjnIzJmXzEigB/45xnHOJDDj0bzLgryQ6FXC05jOS3UH8ruWOZ
H6D11fw2B8LvJwUz4T/EHh71xhGHLHepZmgBB2FuYTXjLkbqG+V0JnJtwSIMeT54
3Ba0tryWL04rnW6s7QDtLUFtLwaGGssM46ZvFgteFkIxMys0Yl/sC9TELSK/UPMC
7lp49OBEi35kYtivq/dwVr2uuMB/HNJQVd3pbrvrpaYvXukYysw+fGONHdS+tRlj
t4raPUv70WK3tRKfIA8dlvz1LQgw9jH+xWOnX2pXeBkM08NuJTGJXSy6Y5jRSrIi
XhV+DY9JlCH6Et5Vrx4oBaDMEJQBeyCdUp7pavcT6o5Ik5OGYQ8E/6C+8OIk15ZD
ex+UsyDiF8XYe55ho8l6DxOSN6Z4yRoSmxXOm43OVlghrIoTjDwcDJr9tXKig7Ow
cLXn8bCfjuGZmjanOCaaD97h15JS74vEy1O+eHgpZa+N7e4K+L3/ty/X2826N7PV
PTD+dBE6prO0z2NFuyuerORPQlh2/Ptv8Xg2WeFtKD8yQfu13oYpwTcdIddF3w7N
1TS6Pc8CbYv/xWlWJjoEF+DLrYFq3gUBbseVkAoG/aYV1Y82jH4TxKCztHzr8wge
22RZ4z2T2lW1GYzC0WLEpG2NRlsoSNHwuvSgiMp4sKoWMycp1Zy6izDVdVeZKMd5
8x7hmtvA3kr0dUu4W+MX8jpBHR+So7nYcBBAjnZ+wLshfpKdajNkMzOfLnTw7plJ
lODWR/p0AwUkBirl5XePYoVdMNNUO1Kbh5GcjztFxrZbj8nO05x6UVvIyjvvTaFB
c1dfqP1LDsl8hZ7SPeoXUO9LgIruhO6s8yARpEexCZjYW0YOe1FWxhfM0E8E/bxi
Lmmyt1fr9WB7owvU2mR4XGenbXtQgmilkLI2hJQ4GfdDHS7K+u8CxO+p75O9waqY
8ZVjFQR28MRkPhM+g1mqAjK5SOylnPmUgKj0nlU1ScDYqHaZTaa2Pla3WNj9vUE2
ytBQ2VSA1Xr/6nUhpthOb2457B7StjHMcAhM+G+I8xqJ2RCrlH8zvnrj5iKQuC7I
BpU1/AuQhQczDq4W+xeOOmcGNYPgkhkLi9Zm69YX8W9SLHdZdm3OKXTIXZ2D/wqJ
kx8wHY7bB0r+zFM5VnqovowEbsnaiSuZ0Sm1JQdmMeMoTYgTtH2eIJp2VH46irhT
FynuPk1T1fEn/S2L2akYKAVTnDBjlpxczj+CWbP02EjEfnV5dMki7i+K6usTF/6P
5I82cf/De4NEEX5dKx9rOOPlrrQyOeiOMBAPzPYqrVb2chW2OQ+Hon2kOkb5kPOe
FcAV3S74kNGcZE0RbvUP3xIwb1rmIp9hddVcTr1moctGvsIVvdqGn58tcrGW2Scz
20ky47yniOq5Cqjz0XGMzn0dEmBviioOfcUcq3hSUj/rudChVEez3Nz8z5zqHwHL
wxk5BBPM9Kkyhn4/o5xs3VikCwiQmVBSWl8Patphqpyd+yhJGsx7g4qnnDLqeuyJ
9rlY9NGEKT0G9CWpOStY2liK+WLAtLBswIcXRUBCGUvSlHBfYk78RKbmA/KT0cmA
DjHkJWtljP47Yykpvl1R/jqGS2BCgMteQ9BSRrYCPfnOMyMiFuFIm4jzAJfjwwZr
o6bzkXpsQVZwBs03MMT54YQbe1RhLPhiYPKzfQU71h2smpHXdl6dOUaTbUP6Y9R1
YJqS4NideER69xQhVaOp6klxhZgJ0HQx6voRrGQnoII40QR8bcAo3g1lJd19r4bi
Mn88Dc/4Gj4/aG/gWkOF3J7FgcVgaXwWGZ0HcOEX/gvYifPGyKJoEFKePBNxWF4Y
7Pqjt9GnU/bMo75kQNGD9nI3zouDq2has273w5bEMP1OtM5Y507p+tpthFNzOBou
ZVenZPJZ0BuFXRcHZ9a1c6PpZ0VOfz9svoMNimg2ksUjHlOmGqic2uTukpoFMIDz
nJnBHtaZyDOVqvEOvuoWZzjONV/QLuxucm39wb9u4xAHCtBuI8ByVs3LPTZjuMV0
g2Yyqmi6nUDS3Cxx/dGcSut6K6brac+riXIA8Zg/S6+yeiD50DmnYvHIlsSBGnhO
xoiIrw1Nf9B80SNopVAwSBOnBbOKzo466ypHGrhbwcZWV5r5bQSHzqZV7lROUr8B
POgmFRh++gtCIfNxaONC7RRFpgWMwGwGIDDD5jKYB97NoDucPGtyO/3OaI1AGbYs
cIUYD32iL36FhFn3M7rDJjOrYryDHqVDf3fXFe7RKHcBzwHkws1AmhFC2RB3yRgm
/H3HP29Klc9fhuR3I+YYE4Zil7OwVGLPIecr43a0BJS1JRqiVDAMLx+gNDiLVwVT
JnwqN7X3iMriD3ke4vx9ZbkSTy15LVS87Tyuck1/E7QN5UcYkycspVZPsMvHbEjy
/GQnaNDJKpEObmPHhL7wtfeZ867mZwjI0fAoiR7Qoq9dsVrZyNm+S14MZi1JemM3
hRY1YNfeyxaHKCr68JS9BOyvzweiA1JYO5+7hf0yvSxcQmxIi6AhxS1+WCIsIkI9
J/uuMhcQt3OhzxF5PL1qrJ6zuETyRN+6NJWKDfjFJqPOFr0icSAvU62EzIr0oV38
K4JqyPr+I7dnzVRXr1ICW8X7xzR6UcX+AbqnmIFez3fZ4xCt+edoPWi903wrOfPc
C7zoXuC6qF5EVYNrA1j0GEv9Pdpr0ggkkCnJ+/gF9VsWxz8AWtEVY6piXoF5TwZb
BEwDZWqrXx5fCddtLQmIftjxvnV+GARZt6eJLp2IESu2ojLpQrGAjlfCmIuaMa3D
OQO01fhHTysieF/BjT0Hb5ysdLGQKFZoVDeMyPqls5XFNIgjMFb6kOC6jW/z9G/b
wwzfgVG/yzK0kg9XagrSGO4UOdIazzA5GYsEZmLU2bU3+4jodMg044mFW5pROv3f
N1ngAhm5li8P0p4R+7LPJOBhTtl35cOK4mO8ujl6EB6iPhIvL/n6y9Q5e+WKy4UG
bWnhkdcfyUlFXyD9SSuoytAntROBkwI2q89VThyKNeHa74aPN2PF3lMm+ul/ooPD
cdJLxzxx1yrUXnM/CPMMjE3f40Zc8SB13/QGLHjFl95TmuR68JaFOKSGRSA0g3XT
9SshPQGQYPUVGD87HW08plQQSa6yalCAnS0DpjORt81CG9y0jSqTTaPNvNH1mR0V
X3a2dgm+ZLaUJFtbaX5FYzZTz2dGs48rUujNJAiIjWMDeMfr1WITSMMN0ArCwVkf
aXW+aEC9DoxrOjiM/SLcYvOCWHd8OkJ1rWKjwqJGv8aRfBLsDb2delmEvJ/c/vIZ
/H9Ctu+Pxdbk0SGGPaFYf3601VryZ+aBjnn2IdnBJ8j5qCRwVBTUL63n9v4vcFMO
9fJRB6su9TpIIC2lC+tvG02N32YioMcBTSYH+se+tdK25Ta1qP3RjSb6jBi0PSTq
hmLbibc7MiYCzKUQWPRix/+7u5//jo5SC8NwHYcxEiiahDH0EYoP/h4PA2SKRwPY
SKnL6GrE2pveWZz2UK2b1cZRHynBZz9DO1oWRvqG729Ds4ePqkt0d+PEfebfHnbo
ALL5hQAqRG8FDfHJ4WXO4Ft+DPeg5MbOC/NK5wcJDnAS1/LSddbbDwOFlRPglNcz
jcP50lffojCsugQKFkEKHtLZ/BJUJ/2/BZaTnH0nOwkidVwQzEKCMP6RKXqf00LZ
blK27KEnD/g62xC1vLAr02TRpSnREiq9JiMN3pMtXSChUYPLwfxsray5tKAV/GjW
asnu/kPpo2tTx1TI48TCaYeMtYqIwYCKebOKo1qewy/NqcFcbgLKckOoFZQEeeUP
Bz8ek8eiazrPAF0BWcyx4FXc2wZgNtFXTvlOeW3sna/ZE9OMZ+Y12ZjE107Qa6Bn
ZE04wEq36Da6ZTPmAyY/StwnLZGApHcbaKrbyDBNVLFfsuTe68bxH3bkuOSX9/qg
E/3h5fubAR5/IqWt7DnHMMziFnrRaZRKOWJGd/99G3uM4NCxBXtPtPzsJhKTV5jL
91LKeu2BYn78R49TfbrteZnLYMW3MRL8V9zCPhoY6YzECxMvkyPR6Swi8ERWP86S
DcIP4hW8hXqwKVZa9JFzoHfdILUlNZBQZu921uVZY/Kd6f4epsRiCwY5LK59XaDz
urxCZ7v/R4/LRcQljBplvK1nARLH9jYn1XNJnSKxZPtCUIajyNb0dTbafzb4Y5i+
xo8KUj1N+tYx/kgKMJzfDExNBADzGKfUPGWN6pwk/1mnMStPG/OJIq28bfR6O+J2
reFsqb9TPwwHnuJgJ0VTWQCIdbacQZ9jeYHlmMRJ+ZD0YREuxWb35rCSgnUXnooo
a3KYD5DZWU+uU3SdnWgd171E1+mzKII2XebGrNaxDEgaZoVPJiKpTfjjy74PkvWX
HAYqAezbUXN2opHRC1khda4z0mMn8IPw6bo+ZW/iwZCxRXb4yFktqS2emWDxKsBl
J3DPK3ppE5whkep5YSnKUMTiXTTEpG5DU2hEdBA49ZoJqsyWrIaEW1AEPAv0yqBc
S5qL01m+MOQiB7Iql8Y/Lx7pCoAt3s7A1Js+7RG+xtE+34+C/9PoBtDuD7Ff5mA2
WkW7mbfF/soycLYGeHNCTNiJ/rxEppgAefa5V2J0dkSAltGUhlG6xG9CF36d689w
fAcK8ym9S+JRIj4gTBY98zcLOA9SPRy8oe6JtpZvDvL/RZvO24Djfn9AaOkuBWrD
J5GLHLoQ9VeAQRBxWbg1KxACzLWc6WFAaI/sDtsen4mX3Mz618GcjgfD4S7omRG7
AMwYX1FFgqrXofOur9X+EqqpL9cLAcwdzPkoFCk6RfU0G8MsReRkGMRX4KEsC+PV
ADMwsmKNklXytl2JdyumjuLPS1J6zKs9/qgqMT3z/Y235kGkBwgKbtz88//5qgcJ
gQZ/pXoZvBhifJIeaTPEGVG/DVEqJMqNMdBpoxKpN+sN4SPS1c0LixhFDkNidphs
2n9uqyVBU23JMpaRSumExNr3FZa69nvoJ+fBrhg4+fFjK8H3MYaYebw0vOOf/0Yg
EAuqB2LzyC4PbE5bOHFqh/slFLeRAKQnSjN66W4Gd8SKN4+h4N8Rr719GOTwIj9e
I433mNId9GLuWM8m3Xjoqo8ea6tfJZogt3tlxByfb9aMLLVl7PjbAcldai6bL5LB
Ga602hV0GDh/NODLQjTqtYN8O2PoRgHQ1FcMhzsK8OsVRSypcbJMXOJyu7HpI0Fn
urqvRzuHpxwn18VU9or1HBdY1x+8W+CeqoXsx/kpaHpyQxywYZLqhmeFi0i1nhyN
EGgsX6G8C2tuopngt3olVYxa/hhEIz6iBuAaYZTQaGUxTDiTYWqa0pIfXFKrwWGn
LltwfCkBDFdb69DG/dWeiddMuVZcwRIj/zg1qgXrxV4HhTmaPrU0d0ZeAOUPbvJB
5dCiS3/+RrZ9wtjOpZi2yTzZHTQHERP3UtoX6kUhLpVaMkV6ffmPFhle6uXB4eIR
VXMKVtlkXlfSVU4ehg3DcfYi844mJg0QUaoke8zl2Shbwu7gCh2QJ3KdvQFiszSa
8Vj6fDF4SPIMYwXB2f0pRP90yV/MMo6eu/zG6jhQdDlLNNa1nsSy0sJPyGDE4Jbg
fpJ1iceShh4n21wfRKK9ivMg3a1l4JOMxmiVSn/9kjobmUFRICOax+szSJXAgW5H
cWkWkoJeqycdI8bD5pmTtG+jFBsRMTrcrvY1AhCrmGx34Gk91yYl0dFygNSMtGPi
V4XWT20UIbkauAMswJQRHqpXK7xYHaMDV6ZUIRn1LxV9j1lhCNjrzK58G82wCYqd
CFXlCNBOWBwU0jnfSWBMimoEektgVGAvIx7n7tyYA2w5Ra8tq2pbWhRrero1K38p
zPuPM1uwftjG+rrQYhdP/LD5PnmfFYTIq0tophnzGLH0wo8itbFueSTPanrK0w5t
xMh6y+3ZW9qfjqR9g65F7ShB86mNPY3E7qFHXqPgo/lc5+VrF0XNfHU2yVmBhzY3
RUiwSUPjNJ/vxlCMJk2kyuLrO/Gnkyx1AkFcqe/actGoR7RmzsbQBSERBCLqZO7+
eYO6wKoX+6Td2QpDvpxo/7liBtp8njGLEDmddY02SM/2+E8nOVb0qrJJTu2tOeHW
Y2p4KQz45vzmRzadnUM13gwOgOW40mdVjZbmnvxPAMKX78bb0CjdARsxY/3WvzCB
6ZAzV1XZ94yatSonp68vn7yCk4zgfrRPa645vsBsjeEzQ4M3zo8mng8+qsbHyvGP
aSw0I5OZPw7yyT7xZIFVVd1RP8bydFV4RReuFQ5R4UeH49Qz6OLK6vu7kpcItUeU
hZTNWkgUwsKQ/JMds7+oIaJmwPBfiyKtd6qcboXBNXjH/SgtZOMQsr+xb+iFaPqK
8oybC2CiC++KuFM1NFUv1x5faVhuD+xz8voKafnnaWwg8XiJe5GxrMFa/rMn5hSf
VggcsJTmxXyD5/00R6mwoFVAu0yCAGnBUHZmDLKnQtp5dBjjLJc7qlsjyVDb9iX3
HNUsSUjBRlNVmIHAiiDKwBlfBmK/6H6mqW/40XojG20oYdg3QIooxfhhvZXRYUY5
+ps84iW/R1j2bi5LjYxdgy60DXQbDPBD4Go49NBU8q4G+IdiAnN7AmqRQVCbj92i
OExULuIBIuQZ0t+oiBWxrnvlYHHkG9Nk756FVnLVho3eM5yCG2WFcq+TzY2Yl31R
cz/0ziycvx19DMaDdm96issJT5SDd47iVsIacshrzoAoZ7kX9OVLwNXcZ7YvLIxv
kJZjQMy/mZXgSIGtoBeY8S8NshbVMNc1zppr/nG+dtkp7Qpjues1vf0qCllNAjtA
3iy0qbsFwNcaSLNeNQGy2uo+A1WG2At/BUGJCFrCx/jFNMb+ld2wqiptb0OKUg0S
Bh4wCXG258I5R/ki3wtigoj+xspBeI4XFq4denrBu/4uzp1o3Z61Qw16l8b2lT5Y
5ylzK5q/7B78weJXigsfEPe7QKaWgZ2ZM+UNH5Kw/JSlq+lkAHGIAmp+UMxCyYDC
xFP8oM9MmAD11YT+V8izgb5sYhknB0WGg0PfKGOa6O0yzH1jMKOl1mYybk/KCRIo
JGBFQ4JWxDY1EI+6gNNxDfVUaRZqIBR5xv0yf2DxulCeYIpkSc/b/NjqlZjcjcTG
9DcPkTE4JZHVfCleVKD+W01BlRio1bZ+RsHdnMpJG9VoPg8Wi+ut8bqETc94wQAD
3ZtvaRqoz7APp5NSHd0NI5eVQ3GH9Qgs+FX/olA4NeTJYjmN1IO2c5djtd4t6tdU
rrmruJa4ZOT/CQmRQIKrWxPlngBTy3i3ODMYTPrS6/2XSPUS4OwpVliQa0SqLKOQ
jqvC9xsMqmERiWLj1NwNl4JASmdFn9wKqkjAKuf2ihkbwgqZbJDdkwD5eYqw/iRs
+Z81We3N0YsfbJRzcjA1yZ5qgIklrEHWeYyX+9Z//3pebf2QSlr7P3rqjfHwgo99
+coZRXZHu2+cxgSJOUDAT+mxdn+uDcR4ZS9Nca+AEKHzmhDFSvTt8BUIUdO2G1Bo
6O78hcBxw9aMeEKR7FDK57FaKl8uDlaTeVtYTP9xhJaMPLx3JtmHEQ9U565E1dBL
zcIwxFV4+uHYyPBd3b9oIIHVDf9m1Hhkp9i84EDFmboSQyQmpUQFcnlWb1UohyqB
5aL4Ct5WoBf9Na1DXkSefWns74RHW3mww+ywNtpoDd2qyi73apUv8YLCV3d1Jt18
txFgyY7gLejVdBXOLTnErwqZZmDTT5di9wgYuTXMwxCM/f9x11AHIFVcUskbfyeh
p1v4FAT8O1+eMF4I0nHKo588cnKMu6FVoXeB0BNkmdFu7YxWyIVl1tHJhx23wGcY
CJZT/i2sF7ymscFs4QXMHVe5PFdTyr4IehkL4i0ezhxRvom+2XsJvkcLxEMF2oIj
MlyPXKCed9y/fPqbcC0dKE1M9RkKXRMoKC1hdtHuazHIy33nD7cCC3TJdeN9P12w
ImZ2NrcOQ1llNIhiSfkq+C57ozcySvjzGIeK8kAhCsPdqEvQcETaxBIJaEYQ1i86
JDYIo+rYUNLgKA4OhAdUJsCyY9afeJhcBAz8BmgXyru+DVL2D0INGwNCyuXk6s/h
rQDRJtEOUpTPxLxRWqnKXf9fYwK9dMBRpQZs16G7fKNEHA4ZASHZC9tCAnqrwIQI
eL9tEe94FZxx208NLMXOSDnOSwixuyFTO8WNEXNUhBP3oZ9g0sdhvCWvWdMFGSBY
+7E8oguH0L3hiKGoAa7m6QvT3ikgRqJfhFY2JcrP9gUVjgAmacEJX/1KCtDjoD2g
tPf7gMAe7Cj2NH9MlWjE8OuCd/z1xPyA+CQE55tk5GfyIRhybd1hyG12s2sD5LIC
ciLbiCbL9IhyPjk8f4T/w+A03Px45/W4P43H/mrNJcBDNc5Yea7dGr2eaxM4iYBJ
pjTTdhzqGBh7ANiPN6gtIPMh43or6nCQ4K1EkOx7sGbanScsriT/vJW4D6wC1ob5
Oek7wVy8gfT3fRoPCtzUZNErKh4/XmZeJz/TIjCvT6VkvE0TDtId2GIJgOaa/DIe
Xf3dbwm/Vmf2w45yMCVBMctzWLMYG1P4tY5/3ZxOPIzHOqx2GqZ4BfAB0ptt2kfR
S+Lqq0zZ4XSomV8GGBIs7K+buLhqMaJiOZva6Ydx+H8IL6asKNdCPuA53lgq5RIc
pieKmhmypOnAjD4Tm3HHkoZ3EuFGU3c5EK6myVmBHzT+1KsFyrCz5DX5BcS2aUVS
ehFWWzHqrxvODM3BrbrTH/4Ffcjn4jPl61GRszi0fNgnGocY7raH/iAMrOFP9/tp
7XRyP5pK5WQIRjHfnGcpyS4cHGgUPIKIbPlqb8d7OuileinoQD7h4YSLgS33LFNQ
wc8rRww0oiTpyHBJbSRmD9TjCpScSWsPnkC806JGbuW8cpQzIUqQ18IcqLhTi7VN
H/uprfe7jZdySGhBN5UaGyJ4jg+RluahjxMLpKgIC1Z7F5t/FWbKaYTN8NblwET6
H298/HaNCYqrak2atrw5Y2AmMZBPPxw76oUKLkoAS/y54Q1106+ckuUniLmfSyaY
TiGZrrNwQcGvFX1dkpj//Q7lqqEhBFUW5c0lUd1T79RfHQT/YTG+OWuuYAx5+55w
aiRNzrJMxJ7Yb53rmozJnJ89q+Wj6ABN/eACJY80CbE1q0sEdBDBKh6n0sVp5FAe
rCf2mtbUnrbhN18zYgB1ag6ah3fa+Oii+3Dses2qS4/vMF196VaZVbHhUP1TiOHE
8hK6C6FTNwppxSBgt/0gLizXcMeJSbvNnCdJ++oMfFR2hHkTxyMzxeXQfCVapHvZ
9mtZ46wgY9Ja52JQrDH7uVWj2df7EgibopyDQEagPAPj8J3O6Dp4AU269JfCdk7g
DnKYHKPOtMoXG2XyO7UtOFrf6KCG7nKQDY0M9kwiUZW6gTqn4//Y+VNTBDZ5cYOw
E9WU72e27FZ+EPHgCPDBXimOat7B2tx1+8MctDbjdZgTv1i+4befJfXgium+WgRy
WUpcGweCPv5lcy7Ew6S84Ff1F7YY1MJzXhTlmSSSD+w9DK/BpzcpPAyk/HopgIgh
Jh2/6JqYdgaOv0gC7TQ3VVxplwXisPHvP0MnQHx/hwKw1GB9DEtPV5ggkWJHbcvA
2R2mlbqXYDVzhtctgvMqkC9E31X6/nJwOkSFJ/hX68RVykJsfH/owAYneeRhRZgo
y3UUQIJ/Zczd/k2shtqiyA==
`protect END_PROTECTED
