`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vIAo0nJCvGdA1MzNPJTIEAAXFMco6XFVwDcl4QmAvUcOJQEiGU8oTywvc4p0mnh
doQ0GIP7erVJ77c0OI0Nljw7qKtld2KZDLnRU6luNByQkAyu1UWy6YQ+ft9e1Ti5
8EhzNt4HVqpoyVG86hr+kwo2dI+PBkEt4BuoFVqq7KC2ci9BYyHo3k1vWpw+7eJe
/uV2K337n9uS2GT12vH3epc2yAQwpwv0oDM7TU986/HRCZ4lF/V9P86ZUxIv01+7
IONOidEr6xQ4vYqOdea77acHzE8fFOlkZpn2vbtNtJika31kseu4UC2qYtVO+6jv
qYS5oRWQG9TfGFHiWdJR+Oz4KmCbxgI04y1bRcrQHcLUbn/89MC9wlP0/SCSnVE7
XzH5wFlF3LHiK+TtPJk1t9qj7E2m1+ChYprp6+76grypwR7+CoAg5sqorVFq+4qR
th+2f2/YNskEFD74DIB7asR9mbljxHnoA7yuLoIFi5yAf5nw4F0sAZyiKblLPjKg
xD4/+0vQ2hanDH+itvg9piopv+GyvDPT7zjSuVjHH8fo1HFYwO71N9WWsz82Lzt/
WQbY34dtJh0LGbLfOKFwiUcNoMtQRxWrKKnlubWOsRxv1p6usuY35DpxuiG59bbG
ZyTA6w0gA0zP3/+682ow0LkXRkI0B7qaM6dl24LfcgBVh/EW6n050DQG8K9+k+7m
b2IB4VHxlErQaJZfpOZXW2RNoBYGBjRy35T8spxOQUy6qdKO5gUVsj7A0zSU6Jfw
EIjzdGbtgGh1h0aF9mnu1M9+rdZwTe23mOkJVFolzCns52JGQQlvh5WTXq+9JtS8
odXX3bgdh8fIsukyKUnmVRuyHDDNRcC0lNGD1bAKyF/UCvjNnpUCcbF5AYGgGyF6
Bje6SB2lSVxhL7x03BQq70+rLKjdMBG18Jry3qLu8x4Ylm74DG3rWBoIquBjuRfT
djVBVOLsFI9V0IowljwsctTXPFwJafkYM5c/QCm62fhUaf7Q0SzWPDvJDztmIUnK
AnJXrp+FnXxn7FyQG9KT0wVan9ptANkZX63593yqtkQLK2XbcZJkrtAuT3VA/ADl
oLCY8OQ3Rm3GA49hKkgCdHV71gMy3eAlDzly7yrFPCzoOa9a9BCD++GEEGAte/Tu
klimnKxME+GBJfKLhIa6KnmK5w7BDW2MFXJ64gaV8TqdgemkA3q0yH/dV2gM7xi7
ehnysUy8IVbHd09Uv+Cm2YOBcrh8bZA33H+YXywkKXc9TiRcmcbNLZ5SZn48NFmV
i9TxW4iydUt711rwfH7M2PgwJRiPj+9/vNlXa+T0F6PSltvxUKjYMKXfHG5nxreD
8bVWXyEJ0l/gw/YQ22dkBA==
`protect END_PROTECTED
