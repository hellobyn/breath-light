`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LAyZrl5+Y+a7N4TTl8mB4l1Una9TOc3H6y5S4G5rDe7KmzL7aWowrfXXGOD2EvFV
/rfMw8MlHkLup3eCJi0MuQwGxJNs9QOA4mIzAIIGAJ3qg0lP70o1N6DFaV6PUuId
a4fXc7MA4M63Hn6tcDEIO0s7aOasS8yFJ7pKjK9AyLL4PoCh+wuwpCKFkurW8PRv
pIRv2uv7bs70cqUUpShsumgj6OjqvaaAMJicH641uUCWxB6MhvTNwX+sYuitUe+g
1mOLvqj4rIM/gGqKJlSmiNmlZofvc4mPZGEjjlB/LouErnkVXuhvhTPyPpqXtgg5
nme3U/Af8/pFSBSJBvAWNo5/yQlSddJxK2R9wmlahtURz6DrANvoDrW0OJpREo3k
`protect END_PROTECTED
