`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tk4dVgfrC6EmeIqD19y5uy1+My4dsED/s+kmXbOrva4nUf8vhjyyqL6zieCFDUq3
XB9GJymokJgfK/6waJVJO9cLCu7F1CFu+Mw5AITgeTsPG2siJWYI4dwFkgRB4DX2
bmGjeXKMgN05Ms37oBd1UVbGoAOwmwOxgM0jGiDfV0tsO+HjOXVt6zSi9DZXocSi
gwfx07GgPoKlzb9u5Ot7uMtPO6hvk056F5GT9ldoFAK9N3D6epxC20rDcrJsJ+4K
O5frsRn/rcrSQAKMBlZn3lzyRzbLCEuTYtatpdNrRvqaUbfgyAA7M/eS83YYTWcw
GSrRLyPT4YUjWjNepUBKJAtzdpnrM2eIc4h2PaSrCSmL6ZhGjr3+dA12+Rqqebzv
deMK4FdixGbSKWsUw9gzJjAYzOs5h6IEtGBYQKJygJhZs837nLk7EsukPVWsU/S/
7PgUyFdq7EDmKYWL/Ym+O8Xp5tlF5/RPAqecMHdwTCTiIxhM4U8o6CqoXX+1aSRc
lV6F4Z3uUvk421bP/XTDKVEjT9hElQnYaNDVX8WceiyGsDLLfWOCnlUyb3HA4QNS
FuAa7AOIiF5PxqjWcgSeuo7xhQBFUtk9sskNvxfrfisZTkNSq8gDOK8Im0Mf977U
5f7A7vhBCnHXyhM4UmX0c+MvnXgebgOzZrFW6W5Vd+JG8a/c/FVu/9X9o4IlXZd1
EDgY3exMViHDEOTV/+G4IBok8jZvaqR4jIh7Uvc7pUJ4kWRgdZFxyv5eXX0yg0Hd
Wr5Mb2x2fOu8ly7WFImE3I6iaE9o3qteRYuTfmtcS8JHMF+ZN+yEmnLuZzlKZtkb
Ow/qAYHtd34YiXt53fzV+uTPyTUed6p7mxSYNthAsTYYFZmQlQOOzMLWeesR0ZNb
ApCyPRcAVmrLLfZ2YiK+Rly4ELwDPCbFhzn1uPOvOnNSt36w/8YBhrqCYg+LRIxd
CNakC0CSoC6VPth7cAKFYMMp7ij6ZqG2lXL6iYDyYXBsUbBA5M6qGLPhw3Sit6pb
Iwo2D0wer8QkEM8k7ZTj95aoOhKq3XYfTLVAIrv9YCT4QC0TPIubrzgKj/ekMyOc
`protect END_PROTECTED
