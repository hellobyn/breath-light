`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7DSFzqpP0WtZeGdk26yvGPH7n+mEvrke1uAPqtAD5acCVPjamj6WVQI64f95UDK
zEuI4s3z82jZnkJ+SuvAiEQILm7PvtWwGfC/V3oEZwicEC6VBuF5pfxlRQqFHKax
EckXlNjmJk995h2Ve0SUof2qGFoG+En4XIBQViSVK2rwuBmfKHgJC0VWX6BvvBxV
ZDmvUpA33MpRVPBVJfEyCewVCrrUUm3kZSiZATNoic3sSKTcfuAxvWBjsicUFZ4+
vRVRlvO6Z6pbFKqcBwOUA7j0LDx/GL5fDXrF/5urbo5Rch0MOsH6VqGPzLxUnBRf
yR6BxN+jfGyCEc0eQh5FU9LU1BNny2SywUEvbzwG4ihM8hxg7FkOfft702/czSAE
AJrMOSQWWaVIF95aHaHm8vUVuwOG2hl0aNGTO922xrcGDnIJ3c13bjbYGLz8qqjy
mv18VSAHVHtGH2dfVLCJdr0Wb8bVvpk2EtWRRLBgxyG/NaaQK+wiYmi6GosgA69I
uRgcfPfm4WJVq+nIKoX0FutbsjwkE6HkRZVWXbaYgzeEY/6bTd4neWX5mMwLFQjy
duceh1XTipGCBway3sbLEPAxW6p5MDeFp+Vg/RAorzpk80irenHv83o4Heewj0yr
CIXhNwFRKBcdNXl/U2SYcs2yyr4hkklYOZ3dtxJDVh70owGe21VrwDVhrMtNM4Tx
F+ELQTWxoO8HVVol8YbBbninXNl/A/sZ9eFHHmakKbnn7yc5f+XNfjzp0ZzUzWL2
BFyb7Ga27LckdRFsRhtxTu+uE5FyaNzOVA3i6RA4h3S3zJsReRCeaUZRq7zFXm0A
6Djn/DJAGQ7YM92+VUY44xM2A2W+7Idigm6hyblwKSvx4ur3zclvisMLQyIj9+xZ
njsP/EMm8iqgHgFvIM5ouxo2MvgeUt8QZWWpc3hGn5+t2BToFpHKnjNTlvSC4u0D
HiBNB9L44a20PGGi5sy7/bPGexrtqWeImkao/UxfsRBVP1l5jVNmPD/rSPbVwQnS
MxanNyRbEeDxBJMIOJ5UPjaBc7i9NHyhGU1eWLB6k5oxHG7FNP7oOPJvWOWsQLqT
7dyB5TwdF57XHXTfl3k7s/XO3fGnuWETB2s//eoN18aaaQo1WTSdLxONC9rq2AKX
xIfGUTa4jP3pykJ2A04Bc4DMuveVmBuHxMYAXh3OvFDHZ0dvH9o5/81JT3dQL3Jz
Xiz1KU9CGgTCEXaEWbF0H3lgMcN8tqR8FmcLtukuRx7x3Yu53EN/HpQ/hcmWK4I8
vcJEmrUAAwOw9aau37j8VQWLQaWW/4ZOUxLC4ziTBgsrwBIrXL8zqxMh44G47Xf6
pU7eNXw/FFFpI9iVhCQaeal+sh5oUQXaxtLx8HndzttphZHcAqQfAJN9uFROCm14
rwOl/IaxuwCikjFWKaI0CsxpbCjSApuc+Yq7aBKAVpXYJBDEOmUn+cVfUYcIf6+d
1CNljUkBuLw2OFij0+ZK2Typ//GKN/ZoGfNysyr9bmYdgt/H/9/PORXRjpEz3Y+S
5IUuY0iwEkQCzVbNylcDauFT5dUUUc217ZDCfB9003gRogFs0IFPlbtRbInYWXe5
FGdQaTOt73mW2j65YHUhnsm6x4oTIUWt7S6+9JQOJM3WPHB4CxXsxZea5m9EOGKb
OGKtzhMXpaXGhKjg1tSd+UjiQyjISGk1pjBOWsfILpcqy7mB4DyckY8cObgCOJwu
EWux/q/8GUO+LlMaY3WOydIiqSzYPENonKQIEMyRmFXeCN1Ph9ugGbUofWIZ15CU
mZSRe0AG2pO+HHtCZi9eppOFCM2w1eizdDJOlupQ7qTdpHf8o0fnwH9KrsSAjuQk
HSkBAAyHWQKBZWK58b1pG5ENscrgSg2x4U7BHEnc5TwmaLYyDiqdYg0DA7Dd3wYg
Nncl2+tSrLSJpe4NGK2J/kJULqhWfdi4zvpLEhayN/OLriYZXGfpYFBuFdO7y5Zw
I9gkHzA3UWjhzuDFGTDY1ZqfGpIuNdBLFNNkFz3u887XI5b54sBAOi6/NysqTosT
atavfgjmCEQgOwJh8b78xkijj48gWCKI8zCc5z5UkbX1zNmc27BFbOxOLffahmAp
YzNTkPUM2/CbnhwR1GnIP97deTUCcL5WMidBI2gJapJ9scDIq5l5qzXk99Y4D9Eo
So4IBQnioPx3ZvCOYcOMdkPwh3fPkyG1cAd2Jqn0S7MMSk/lJ5LLt/TW/D9qsDqk
c1EIAgtuu0m4s0cvzc8wIo+NUyoijTSVS5Evo5XEfi1EeuER+KqFIaa8/Mmx2nTW
gGguHkb8Z4GDzWqtOxvkTwrtvGINtEVNI1NXniwatZWyb/Wo+O2A5AFCRDIF9oXB
9b4BQFp+GyO6Ee4PguYHKM4jWSKs6/iXSzegca5mAIJJAwQa6W/olWlzeI3NxpHe
JHNyjOhmTYQveARQeBcdYQz4LQZfyWa3fbuDv5zgvU3qTU4DCXGM5P7CaNb/DKnr
EaluxEqLFh0XJYqk0KWDZK5BKDkiXQVeOewtskQuhmy56RvtUKvxwUe0BDzAv0Xm
SbqZTtW6EMEkj+IveEQBBpds60Tz4SZQy2igQiPCYWA+4teJZxHtvQTjSGBNilX9
W65oxwDbyEUmVgqBOJyidGJ2ATNcfdCuE5I2fFs8N6PZn89Qn4cLLeCBfMVA+Cdg
EZfJPTTENi7+tjy+fTB+JM7ToGqBCtNzaX167D5m6zYvdEtgxap46Z7wZ9bcIggp
KDWyoK6KJ5zja2CMMyrHQQHO0Nnf2IYxGIgb3cbQcKQ6/D/RN+hZHVhI6DX+/88i
FVAbKUzYyLLbOtACMnafJE63wp5IYeDpr2rxpNqBW+W/RoEBTgnhTOWV8nIvjeH3
`protect END_PROTECTED
