`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qVoHP59x3cfsUz7VMJbfruPzGWShqc/5vW9wkoqYBmSO5edUVbH45kEEzH6UOLi
rFFAXtiPQcmXI644yaAc4xsECOor0rrqSF24eHiw1/HY+IINmt4GETwm5nu4oGMo
gyE+cqbVHzX3fc34Z5fVUWqHoqAqfdwyljpRGxQiICTMqPFyAouV7X2qwEcMAcMx
4crHqeT60tANtBabe1I+MdWMK9E1+VkNYzWbhbwLzcHwEDmltNlnxxdoyuVbNvzz
hjCbq8Ey3hrBnnU70Dne419sWtxNj944eqyWXxIpmv/FGY6ldvqG1ixqNOMlaNnC
/XiuwZoOGGcVPwRnvLR0oXKgSE7a2sXX8ezOvPbWHGUftYUgILqVz983zaTG7MzI
VQhrVJ5zmR0IfzoeV7AxJ3dEhSz1DaRhSwAblUdk6s3talA9HQDMJoeJeyDMTpxq
i53U4mTBVHJYhKteYEvLsLwRmBb5g/M8q2rgDugpWMGiA+HVuT48rCSMYKbSoL80
o93Xj1OG/gfhQ0SFxNtFKmm2YlHtt8lpC9VSOcKWHpNetyNoE52i9KC1GxBuVr2g
uPU0idT2q+7UQGvk1vgO60fqf5lJQB17cZcoRnBz3mmGqsg7VVUjgkAfFRrqMQHY
D3URL4/bHu4bTDVLN/cvlHQh2l2oBf0dAxVWxqzWrAtlG3ZdxtdtdcQzXuzAf/Co
2QrZ2w5GLKpw0kpNuko6eJ4S/LF3lYXpLHsX6HXPsg042x4Qzsq41zqWTEpBrKMD
c2bWgVGgWhWBLndXJuhn3SMiqOWzHsTJYdQLBUs8Lnjt8K1gjeDz15QroFjZJlFF
yqvpvkyP9eAundiLSHipA9CbAgHlH5VbHgeHaCRydIx9aCd2udMl7yD19by8HHLd
32j+jnNTFfDU9xgl+agD+Qvdv9jz2e9rwYoACFK4mDJb9sFRMD9jY897WIGw75Ub
DmpRHZOqfgJ8LaMVtTbhrfzSXRgjVta3QAGUTasfAnVUF8b2SrU0NN+aiTKaK0AG
5F7RQZfGVI4D8+W3mvz0/KiNwADMTMCytuPDiJdW/PkmYG1WzwJuIzsKii6VGl6Z
`protect END_PROTECTED
