`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mgtq9UG8JsOH1Fj25DPraugIR4aM57Al1dEbUHRFzoz/DWJp7WxtE0l5iMflBoH
oqIVYte6EMwUHE/hvZvQjUpIju1ZT8rkhJh5bD5hgYmE4YlXTt7GMSXsF6xrxRLZ
sT58M87daCKhGeWVSV6fvoyGIzdzz1aO4k1UAskmZ6ulzdWKAOvtqJEhfVU9JbN+
TT21C7m0ADoCCvQ5Y4AtNmPKi50QwAcSEZN3nmxc/wCOmJt4yAcx9P2tvnW0sDnT
CaUSX5LhuvnrjJgzRevAyXCGn8zUBxIgVhw+tX5DeNxZC+39WPgT5aOdQYKg0b5M
Hd5DfOGz5snEeZdRrU5KrMGK2oWaVep96c5uXvb5wkH+t5uFuqQj0+pnMKpGN2I9
5dENSuIupsSeWV04XygPDrSxNua13RPXoIQ7Bng0myzKNmYx+M77RSCgHVmR/By3
TLQZNtXEbbaL946Lla1gKTwm0mETPe4j7NfGodDGhoA8Q6KX2iCTWdaQnPqjUQwK
Jz8SLffmdF+WK6MRHO+JUWoVKGTJ8OtCuMR3tC+aS6r3Cu6DDkePhU2nCRtVTxWt
UPliO3gpbybs6dbBZ4VU+HdL6ZouFyjL3LKuTa5xO4qJ+SOkzs+m12SKKdZ9oHfK
hF+iFdFDFHZscK3wVjThsADOR52OK16F6MnY6IP1zOGz3wuuXBcBCUfVtjR2tpAU
3reQ1wJLw0FMg0DtvIUQy3vYi7WqV0wWIPJgxhaz15ivMOUabgBERppaaCi9ivU+
eRLenAGtkSHvofGM5CdhNA/zCuFxzgr16nmQJuuF0IqJO/fiWkTiiOrXIilolZyb
lK/z9TK2Wz2UxHZNVs5O5dnxV7/5MbPLIOcigii5PwJNI7XNOJn2XCDNWqlNilIP
K2ZHlvnV49ufUUxPFjVPYpZPLDv0NE6bBVVPq9d/0QrM7xk1gD7zghtQLyUx5xMj
ljTS7EqBtXKneitHO/+BaxK0W8diwi20155uqQdToERrqJv5Y0soGa7yUk/J3GpL
TSEYCE81EgffV8XGG+W8JlMfzErD31HRZDamnTDr3L8mbLmAVTywlYzx3qfHiKof
1GfKFZFsgIcF13bw5Ocqum7bipHcl6aMJVrPsTgHvhX/pMZ1uotIzGKErNoLPlPR
PMKFle1t/OfGDvyDJLz2+G1f9O6KWPhVOcftY1a8znxtW15vwBfNZhXfLmNpDMGh
awTVM+SjR9QJiSKsQTNtg5XYWurDsx+e0Mx4cVbG4uZR0KvZKMIJZWICEmYE3nO4
j+zHkg7dVBnBJS3CasDdYL4QIPoxLPrsWQLGTBQsKwauFv8W87INsNagqtZgn8cv
t7Lvw0ndNWmbReMy9GiMu9KRoXEsshYrGRvCNpAmeG3woehcUr8xV9TwvZfjNsT3
kGlVgATFuJQEtGoypNpEww==
`protect END_PROTECTED
