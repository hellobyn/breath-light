`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ryP95d5JORek1LrjjcI2SZE3xV5tNpeyr+RHk6646Tup558Bwu6DgyXHiLXwUXc
3RpiwBmL4OiZ7SVg5MYaPsgJR3nIX0FjiM5hlc/ga6wToPvO8vKt8k/mIDYUrNNr
f2iQ34ov0yvrCP33VRFFBfZ+XcIC8PDyCP8Af1NY0zU8/V7QPdlI88ih3bD7kDPT
B1deYyiZyougAXK+lqh8gZL4uWfIJ5Izjbu6aNDVlhQNJPFPEkpyCD1/XZmQnNv2
a9nSdvyDzcNMH8gaBLD1RQN3G2dnRxPHfsnPeAcSAju+D4pvxDbZ3gZKT9YwZzqt
JGlkeWJkMnbohzMMLuZIvjSUl1IyDXAFb8N7IQXNEa3u3d25W3X9tolqm6K/hDwJ
`protect END_PROTECTED
