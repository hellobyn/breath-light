`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnboJEgPrwaKvOPDh4TXSECVGd12Qwbyyz1W1vqZytpt6bfzcfgbZ/0hwRNbLaZ5
SUhCLOyHjHCNxUBm3ByTvQrvHEyT9AgTe5GraTYGIvNjEep1wAqpQoHY0Fk00P0H
IyWhlI6SQyxOICVXTi2aub8N5+Wqq3X8sSXGcrAUHCrVYFYWvg4I+xCxZDWTJNLu
`protect END_PROTECTED
