`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKc4fXmc4ITmwqVc68zBW0iZJnkkhXSgkmsuvkc8uYwgkOM06TeKIwVBMIOCeN6G
7RBdVyR02Yh+p/VZBEEXpjhPyCXcaN+QB6YEBWsQRcz2q3qkMeKo2Pcj6crkI//X
Nxb88RBMQjRXX5ZjV4ZOP7MpHNzhwVaKWlOCFMxR64xceW5UKGaEHLjtoNFIYysB
xalYTzCtL2LZXgL0J1iE24NHEcT0tfpH4WI9tYxd8Ole+Mmx5IxfhpfsA9zxi5AL
w6zMwDeIgulVpT39WHExfnSpeJC/+BOub3INhCyuvdQONazzNmw+KXZ6/ziPev2S
qkxyt7hQr1YOOfgl/WUfvXPojGqI3Ni41cJw/DnDyra5DwiVTMLprO0nsX6Mvy63
/2zpOFFAgc4+M3tZNIcdVwlSX3RqX1+O1/Ip5kSfcBkuyGBXVCCoULs5YwWfZXGq
ub2aD/I5gIlCROj8zkZxrcqHIjPsAuTFS8ONTZdpHQDdy9S/hoUk3J15M0jGQKT3
xZLvpbxc5OaTtg8SmdCHiKD87IgEU5iSevoXkoipXfK7nj4cia2P7b+5ATnQlMw8
z67RzLd7zYywD8TH6ygN1LTKt2KHdkUPLjtAs/0EKn8ZBIUE0W6pUaAFa31M59cu
WiHf4RFrQ+bR2bD7Bqu7D7p09JhDKk77o9HumCzYJgf8cxfQy6wrHks7cBvv8azn
SaKZhOn2rWR6FdokdfgMuAgpsWjqEqnOiCbfUYMMl6BCpwYGkacaHgkVwiEt2hfM
JOxGOQSFi7fa1R9yBcEQPiCoR0EEbX98pXmGNqQgzJ07ANaPjAbOSgfSwvm38h0Q
o0/9JSa8FNwjhWA7tdo2pYjyjVCh4AwZ/VCu6XLtP+oMxOOTBG05t1R4oUb+G96v
l4CwlCOdT+chmdiqmniUn1OyUObpjxK0TMZfPNcJp/Eh9/yA2fa91Ni5+ovxLABz
rt3sNe+V4rNsw62NM43b6w==
`protect END_PROTECTED
