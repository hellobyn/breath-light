`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tqqijvco12/amZiiaxj4AWX+bZelFXswvXLmsCJKXyc9fhn7/xBlUwnZj8AbuRKx
lq/KiRJ/8gVW+NxfaAh0Yc4ORkOCdIinAhoern/1Hnnno1lqMujqQANGf1JwvP1t
h82HRbu2wfCkSFEWP0ZyHgw2sHmDsO6EiTdrE0JgA/b/jb0pd73MWpdlM9WSVEYc
Le6dCkR768SYnSoJFmR67kj/GBa0gLLeangBTB4HtdR7zVD2npyXzAd9tYisM7hV
tD4MMSFCP1Xk1AYXX/VX5bnCHwWWA7NxgNcr5aTosDTe8y1E+4ChlrkMkrGf3gvd
ez8n+9SEtDKj9eGG2ppiG1NBY/YMfE7rJTfbXczHhiTyzc4rpGqs6HKJp/v4MsVy
wJk/2N3fc6ftflS17QsK52RevNiSrWI0u9upvZHlzcAwfLU/t+3rVbf1CqlmMpJ0
8jhur92MqYX7/prisgeiZzx+yTXYhmzj2tQLKAjagF2qXcPjKlPMCFXADanPZ7PD
oTreGLRfnigflNjUeamHsV6XMGCgy/EC9TmEPbHhQbQ=
`protect END_PROTECTED
