`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXRan/qavutBA9KITcv210c2u5H4GcgQAUw5jhshD4hGacyjCrOg3ZacCgmkeEaO
3RMHIsGR5HLblsA4A94VC7tEnZ7FraekwWk15nmzA8iKJg3jC/DMfxk+7V7jmrMu
Agm8jaOEjpqFUUUl3Ab1m2nZUvFPcuvYwk/Ykvi2c9+T8CITNJTqNHzYI+5pDGQy
m0fArCg6MCh5QjfAGhn3nfZfg0Vzp2ribp95ELnel+gtK+3mYi4FgLXVqD2fqs+i
bRGWjgXM+RAgdc+jKewuj2TjY20j5aNTrKaFC3B3LxRQIAFJ993pCyx9hx+kwxyx
G/Kq7WvwpexlyrTquU3xfloYHwPCA0ZltLbv92clOITxj4AdRTARfbNfZnHPZjL0
3j2MtfYs8Fwu0nIebvHATmlBaYdeN89Ig5bVG7OErwGQNya3sXPOHgGK25yos+sr
fsIfPNKjTpri+zHi1vtpsuOI8IThZQsTXiRY5z2I7we9gW/fZV1I5QbezbhtbEis
nCH3OWzoFInQdsvG3adkoHtORbL++lNjv+PU6fn/9tuuNTCb47maoqggwmblFK7h
CllfhvINtMBITEFqOYFD2RmNDAhGW25ECXZxs3giedb+F6T7gY65WO+f/q3uDQ+e
wHmD/iJrVC1GEbEId7NNo94j9CowmP+Jd2K+esAX01UXzAKKILlPS7wPSlWAw/S0
ISAvgki+eApGkMAoLy15wXuvt8PUKl00RLmW/eLrnT6ansgGtgGEz79U7NEnMiJj
qzHdpnIEnVWB5LLbp+I7v/rm+opmEQn1kxPQLMrcgmzUtKg/PxPPuFLA4qyHOmyF
QBILTkpytvnIbWbRf9ArXtjLSsb6n6C2slr9mebDVyy3w0Jy9r0EiIbLNnxyQH05
G9Pd/L2nGJtbq6yYogWAd+5XK0KpeNLPiBDb5dST4p6yO0poBv4vC9Pt7NyELay8
gJ3ualYczgOc2AHB8cEurXMDNkyYXJslDVaqc/wwm990kR3AGWGVKNq2RIq5T1lZ
IJZyX/xSmmG1WlWFKiioeTgmFJIEdYBWp9Azc4q+PvYXTNEosxv7w9WIbteoQK4E
LIeOrH1V9X9jIPi+avpPhoTeHmAvYDWro0LwbdtZ/uWKzu98ahSbwn/4N+amVve2
N0qQGbBUN6iGCf7BqCpZh+0IkiRQeTvsR7H7L3TOwPzcJji/KqNWQLddX0+z439B
Wl/MAJ6kbY+ZwFT3d9FG8u0XP8vzjv6ypkDm6Lq1DtdCEedVByWKRO291bWz8pep
/iNohsVRrWJQEW4IDnc6bLITw8/n9sGXOENOtmISOxtdf0xCfOVXcIU6pSKopQ2V
Sahi61cVOiI4HpSojvZ1RpAQShpw/bdMZuGYfPO4XKspJjXGW/SO1ZjxSt2rmysR
TqfHNVTUVCCGuJwhXdX6WLo4mpzVWBa2AmbwZ7hvQpxyRWhlwNiuAJdmYVcapo02
0FFc4n2BzJjDJYUlJctv8QCRtwEgyAtKUI9zVbxJ390/ET1nUiTJeC/ApfqI/I7B
IWPcusx+1Elo2AOAEVTt82XJOg2Yyw3Z77qN7MKIcn4/4qgkUozTXz9w9VnEY978
Lin2e1DOA9wr4SLluDC4euTsxFNO+H4wV1qXMWGxTaoiv8CMgXKBKLgQ2I4hCZsV
3FrXjXQi3QlxnMsqkcVh5WaTWSSt7SPbj14OLCBXQp4S5D8g03JKkA+7z33n+U24
Pr5LUE0OBUZ1eZz9RxpklIRyKa+dT3r26VXGTXpxlcuqt/GQQFpKaK1V7K6TJYdj
DQ7IMtggzvDc1Gqxs0n8dKymOd9hAg9cOQNTbFxK3x/y6b+k+ghQgqYyIvQa2T7f
rZZ8dXxqRtjkO68ZDR6EFXRA6Mue1Ls4ZreCIQqI+ut1ZdOS9xmadlI/6wIcW4/y
/ATY02ad3rRib4v/m60wU3gCQQlaoTFYyuC3dChsu/ftMOqtNAykFdoCwQVirNmn
GfH3McD+hW+ssD603STWHjgHKOjK0NO9AZXAUiJEU/Hk+a32J6rOOPNW5NOO+UXw
e1aXZooGT9o/YW/MWXTMU52jWHH7aKyai6GhSbrke8K1AGuoPpAfe7RxA1Ddd6i6
ygTCosPsAf68GfDFIUzB9EUB6FOdfy7dzmk1KquvrjG73Cjp4UFcX6brHwxXkShB
iBqwe71mKWzHm2ZIa6LfTGX+MKKiWxaLTWFJ5IRnox5aUq9VAgy92DojMz8VepNX
iIsWOZe2LPk60a1aOd9Rqv3v0Xt0oFqDbZiKzy/Bizxr1x2JhtGKjaV0Ftknxrfl
x/nfu4qdwz36ENKaQSlP2FqFItq0lUl8LOOIVWVQehOLOGiMte7IKLUeWEpqRVgt
ovLoSFzD6h0csKo7l9O9awweNrvqvSEQttVBUjJF0PLO014CpkJU/lxjwAavdAp9
8ZKsgz60VPOva4zqsmfeaaXMSo7JbpgI57WvLg3npiNSLAApV9rroa6nFzisEh+v
9RjAsq8449WaDNzU+1sC6b2iV7Y+YffiLKfyPl9QQPRbscfn6zOT260f4lmslBVt
bHIYJ3uoDemFWsy5P39EbKGclGQp2BQikbFX310fB2kRUk3Vx53lEUp7JsMlrwzQ
sgDc2gMJWz4C2h9tcAbXg+6jZWhw+PPf+eLW+exKa/e5+VP0JEUrMzFwlt8PK6is
855ktNZIj1S3ViNmlIUbK1CYV4rJtuzeLSnxc1kdza/2Y+w0cP7mIJRsm+gzxYTR
lFrMwoENAnvOB1ZB0DNaO+0jTW4DT45kv17vHozctMaT8SFJ6FtHuxsAL2Id/k1l
Vevjs9RcxhsMdWlgwFuxQXAS/e1jAdYrZdElou+0eW2eDIGm2xQwKYSSiS4IySS6
H6zW67ZqPvxG2lh+KPpl9eBK6y1osd12OZjwfUUwQwnQpoEysfujF5UvyW72hZCk
rreDSDZQV+1veA7nXA88mrVCLhA4BrMztcXPC/PDZNb3uviAn54WbbWu6klr57iC
XD9RR8ao5t/00LKJjjDlS91MFe9c1CJ7CABno0HNyZt4aFFBnpBXqhXSVZo3O7qi
WmISIh6ytgVW4nrXdXtyyAX4uBuLejx1KFKWufYqhs5FHG5eps+I+bogQaQNSQB6
HXB55Mo31Wt4EF0bwTdsLqsVB+cIPhWgUPplR3J65zvJKIZDb8RCKAP1Inwr1F1X
F5Ji3+6Gj4zMN4uhzMcFhihdNDcuUK6p3xgZy3GPWB+D+Ym20RVe8IRas+ZJFiAZ
CkK//YU5v0vIHyduL8YDoIw7Jgv2sXI6unV3CJNd8DoofPUEeSWZ8yWAHNsDIe8c
DKKcaTqBW9y2cBnsExagoPnt1fKT58WkLVIqrXJIKw4xf5kJhENeKO1qV300c2Au
7YPFQVhOxMi+cV37jKnWJEaUf8PtvLmoIgeGH6KIunR+EstCdhXiJWh2lptHPb8V
dO406GDxoidjyCNxf9cZ/P7rTVbZkYaenUVGgiXXs4/s7d/FHSa1t8oNwA83i4Iz
`protect END_PROTECTED
