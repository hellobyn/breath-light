`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gKqTBrdYL0APjFf59o0QdWYpmE6euR9r5RTdtRW5tE5Pui4mNVbsxmvsUs5H3f5
sCFQle8lLwx+U4r3h0pW2Wh93LWYab4bIfyAEdEumXnllvrfD5K0jzzf7gG7nRQP
Egg7h/Rl4jdRJcz0LVlNMsqWyjtLyN0j3peQHQTKW9INzAu50gUeP9v7CKvYz1Wv
wBCbgTzuw3z9hQWmU8rVygJcwpfIIBBKfC4ULC8MKIzComIrnVlhhCQHwVyje7kj
4CwpyykPpWXnNHHNySxS27LUPPIhEnic1bquFcAgelbLifOYH0VdMSUbsEj6kqoX
+XzrIoyIL5tB7pS0GWleQpz1LXeL01CzcwSw0OEkZ5O8Wqsk27JXd+qk5PlyQp1G
ZAx8F0q+QT0m3vP5A8qOZwnJMXN0C1TvB7cqwyJZuia3AbFDs6YdoD3KmEYUPBr8
+w6fzxjHgZY3tXkgKgXqkuD50hHKYRL/XxtUNB+fl96gWHJoHv7XuWIEYvzJNSBy
eZrW0WbwxHhh+O/xHkFgbzPgbel3b43sYP3eO75NDIuUt/j7gLiMAfLy1J5itv9S
14/9rgOxGTb4AePKIbaWF/WFDxAhRLW2sV5migks9mY47oDAUJd8MsjVKw13GHVc
FCoKVi3MxKPD9AZioSIGlvvpRatUTZLdkMLR2xxwYkl/kATpP1z/oQ0q3Bxxhrcl
nSv9s162mYJ/URoeOuYuByxZnaOi/SwOk5ry7NuofUW/kbiErri7aiFiuB+BJeQU
tvEdV34vTvARZrcSOagL3uzlekiSEScXYxVkip9aEbbDls8W2XVUoekLynVKbZMG
4o9j/DfZw3hf5qQ6JfwzQIRG8RJNUUm7J6L+O58enEQV0yWSTD69fj8065/JVj8d
Ckrx5/NlhepZypbszSRbu1NiDsjJYYJ7e4LCQfVb8sLbRQPL9MtkIIxsHmpPoiXt
vet1pEOFMkHsyo3f5qLD0MBgyBqD1bJ4fXCeTjUfaiftvrrjvMKSv2+6FsBgNBV/
ScCPstBM6havPdz5wr2hVL/wP2dB+lRv2PDn9heQuAMKpl+fUnsjPPOZfLL5VPfU
UIExGbtja5gxkOW/2+ataLOunZ+biltyh08kyV67fsfZ3ROkVF4nnvuhitGv/jMS
gs1QTp4KNm2nTBRtCNkD37dvaTi8rGhjOdI/w880T9Et/3VoKfoCb9oOYkcKnqbE
SfGfgOlNQPjRrMR7ALYr46uRWFaQy564IA2h5tADSinjKrYX9/4Vfo/T/ymj3N7u
kMvmy9gJBgvC1zaSo2qvUgkJb+W7++uZrUU7hkh6fDasPG5amrVYTRgpj6OoT6hj
IRtqkX2Idpo7JWEgeyPNvX8mYS82IqW2nziSTKqwTmWx8/oYgC5lXG8wqNaZDrSi
SAaza0YcfbzyjBfkrMRaxjvAvFJMj3E61nSLesk1baMoczfQqOOfVkgOrMR1sbwH
5YdDQMlOCKfwg1EdJGFm4owaQipfvU3ebgwy+ErSFSS4SBEF/nvs9WxLiIi4ax1G
OVkK1/6rQ0PYJLRZBSoeBRaNKUEvGtRc8oqfJCEhIFs6V51W82sOnYGFFU2gnybF
AIZfXaWaNVihmq0TMFKOen1OwXmjPZXmyJ1bN3ksLgXBQC2vqLhwtkGQjhcE2sI3
qQWs3sNd/q14lbcy40+MROToofgjWMeE4UWXnrQczZLxNNjuGsjnT+NA9d1qV90G
7pSmWmGBiOcKg78WJjQ9CIWFvUt8++nAMhV7xSNkis24KJKYAa/9WYapb7pj7t6D
20Q+i/ei3WV2rV6bmB6rwg8G+K34m9K0JftM5ed1t3mK2Mzz9JUME5K99S8N8NFr
yUVYhanD6J4X0i9PNfj+Ts02FJjRl2djpLcL2TAEp/aKWyoQP769z/vG8FxzMsZo
BRPsOpk+p2DdjiaV47qK5qrvDbQFNW8MbI6emgZXVpxxSThOZYx7wCAKPudVeqqq
7LgLuHviTPcgDkUPwfHufbAhoZzP/xHdzOXLerztlVblETk7UtVYKXrwPYhPc/wz
rz9jJA4sYHdXEeWhbwFxTA==
`protect END_PROTECTED
