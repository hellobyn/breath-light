`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mcv+FVpcCNbXpuH3ETCdWPAXZV1Pmff/5e183yRahHxDAQGO1sSB0it1Ma5yQTRo
9L3Ni40lTedLWVTniJjebN79/fS8uq2t0MdElvHbgEFaCU9s/1ZJs+l6CxiUZbR9
4znr07h4Ji7Jg0NKMBCkTB3HK4Z2oyQSNpiUczHZnCGVdYFCXAV/04x7mD6RbAqz
jcfX+ZAdKjToGJmuJRtfeBnbOkgpOH9LN2jJb1qG6izBwliMDyL2cVa4z+8qOC8/
OJEvTLEm+sJC9jyvaizOAJz2ikWein9GasyNPmLQMK/W5hAxj7C6x+aH9cChekDF
S8TrIfWmd/EYgXriv3LtxONqMcH+jvQWIau3X2XhlrwhLiBU3Y5W8jZUV0NzBwK2
eWP8+uIG0cucCH3ah1i7xiv2X2wlWLuK7MUv2do3LyS1nlT6LA3X9kI9/3Xf8Fzk
+dLA88j2oHBpjnW44cY7brEy0/mLtR4Nq3lgFoWPQRfZB9s8vHJt68HoU2gHuoo8
wGCve3Nws3wctMoEZNPNKYwUJPU3kOe0lDhmEKjkgBtMql3qfYrRQfPJ9FfCHmWX
rqI4jh4Zu2ktzjoqzy18Y+RfKwC0Jeq/wud8SAgh2RL7//8fvXtypciQXkh2i0kF
Lo6U7v/qnSFpZUwZwpoWsRYLdvwA/vwfnxKclEeVKWwc+R2GUrn9qwhWrAgZNAoY
nXPNC0OxF7WQyf8k68NQeGA3X0k3MttGCCrTTdet+zDc2EZoDQBbKZ0QgCLxPeNG
V9y7fnYSey4bOuA6YnxX7thenvYz6ztJG47IUJ9IFLpjvA7247NhnRZRDbMrnB9d
OExCWn9qAdU+NS1w0THjTdfLStqEjOXbzreuUKTt7/bIOYPjcyJPx9NT+nByz025
C2qQbq+Xpo5HWctAL3bQ8TVNOAe36P6yfmg7Y84Ua9P6/5c5LP5/pghEtiOpJ3Fw
9WYsy1Gz73elYOeCDN97/XlbqmH8BAsrunSmvIrdFmE1ka8Ull/X788pRFxZRLkb
3WTKC2DBDRvI+hv/lcpYnmsgXhUYN6rEgWuq97yBEcPRIz57sWbh5b3jSh/GACWO
Ux1LA6vJElVf7aFSOWm6+c+UxKpnY2GYaeKEXeltfGPTpxQlZnXUQVp/x5E+rvRF
p2iK+XkJqCnRF5zhX5PDyqwp0DoKOx64t9VmqEWrBqdvmuUA509vQX3x0gKjfqPZ
hHS++YHY+XGTU1rAvZh4YxQsm3HW+FS44ePIC7NMEBcvAYEuV/ZIoRxZebi0ocaA
QoBNxS9EWzCoCHjFqNDNhMYgN/9KXHQin15KF3xIlmYKK9njRlbxByVqDHtCY06v
LfvgnJeh1Ig7+LGrZRYMHCwiDPvtHIJHgLvWOhXzYUhK+PeNjlJeTjv7cxaAPTrT
kXmPfS+XrvTRt+kNp4ZXRzPZL4zG3yWA2nolLIDyeDbYWCbzMerPPLGBXarOcUYr
fKVskYlny12BxyL3iP46ZlZDxj1hERXIjbm50zUwDm42IGw3X/3OKlvQZhJHOfUx
y5Sgs2gWdI78DBJCvMOMWfOqztq0EJ5u9DrNxXAK2TTrcvI0NZYW7eWwy8oqEHCE
3YRKq2V7BQbzOgB0ahWHGBO5osolYxGgQ1vjkACip3RHR6+8ESjs17iysAVUFwlX
tIQmPwouncWKYJeZxmTAwDCXFgaVmkZPo1ucdgP9iuetTD40/jpkN+65u4wvbjVt
Fib3GivzSYcF53tocMeAqvZyVI+BpXheUsqgRas48Jl+qAklbDMiBBIKTpwCWwoy
1PFuGUaXogztXNeyJ9q44DkhFQ9NlKkFg191RkKqgPmbrl2m6oUQWfB7PWzH3p0Y
NJXMP+qOsoEgrWXLLQGgtAfF2AEoHT4iXwr40vx1hOejC7oTU2HBfI+AToJNIOcl
tK0ChNAx14Qq1t0pRu8MVSId/qJi3JB4gIrnVZZcRzlhdg4UledR0raEDdVMKcCn
Q+ynbfnSgkhDpT/xdgGV1UF6mLSFlEKOHptp6Z8Z/ZbTb3wsj6aMuy6/sTwuNWB3
Or6xTFxxH3I+bun3QN6RoApKzyjv/ODRdNQwt+gqz60/XVudHtAKpDYVBiKUJzjF
Ghy/D9mbrcTAZCygOlvqmgqu1WRsO4Wrn4R0PC3uDd1znjFSvcT2Z0lhkkoYkVhO
Ybp5iNbefFpCk3Vwuo3aS0ClXNfui7coJG2Wt2ZcxyiJ4vN2lNMt0XeoTNPXvk9E
uZ3rxDV6FN7w3WBOCa1+csmrHAH2IjHOIBbVWWJGKxdFLEH4qSDUOBEx6byE60Zv
oCTlsB8axKjq74IENovUg00Khf3o+QP+hMSGXxo7b9EZQHqlIBe7PuYbaV21Fdxe
0+kbkFecMf2gNJ9wlBEzYCTYTrQLrLuR8zB5SOWwYpAnGfOVObM3uPFMMW8eMzfw
qblq3yror54RMncyaJ2GrlZLPUT49hY4Er3Jyo9aQV/YibcYoidbk02U8J/nEt5i
/oFjsANcEaAjR95MQ4ZgXN7GtDrxedA7/wR35D2TpugPvKewUcgwjaG4Ek8+nM9w
7s/oQLlvdpfOZNXrhjqroZi7gbqn0DU3kqBX8Te7D7vQF82Te3m9e+B6CxJPCM/Q
gKnOmcQSvb66YK+XMDl9Z4g9LbiKpXovX3/R1aA2P40FJeeOV5/9INMzQgVYZpLR
9d5wYJD5UPs2rmPvuwdQ7Dr96zsP4I93npKsCV8El85gMwGTHEI704++njJtV1Xm
1wzR3X1eH/tzZYhtItfawQESqoYIGHmEDj6fGIvO2h2iz8piLm5PqQP6UIoPLTKt
uF/yll2O9jpCUBnNUIOthdH3l5zlkym0GL41WZAqfDceULlQYbEONOPhCVFXMliY
IsbaLmHIf5wJnboWe9edF2/wo+kKfBKCt5mDWgrYOuuHEU/hrbPs6ZpUvHqVJ4sf
/35u+s8IhZ0IlRJtAIKaKjS5G5csRgjDNDEQRashsnHfBzjVG5+7w0G9pHPdkpal
SKseUC5bOgKhFzRspd9ojM0TiKpz4prbesGsbT/zc/Q=
`protect END_PROTECTED
