`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6lesadJhCXmmDKZiUoRh7/sMXHJkI7Ntw2VgwXDok1TDMg97iwmZ0rWmRGme5GF
i2CV3uQFBI3ZxcIO1Eo6uBBm7QkvDHO5ma9BTLU/+1tI7TYBw6il3Aug43/D0h+7
H6q6OwphxFbLKuKSUwC4StL+LYshY04ZQzm9Jz/E8HJB0SeIqic188qRgWfI8Bmk
K4FQyCYHyqOsndgIMKXiYsOfTi94QP+K5Oby5LhUnubCdQaFU/57eGM3OmShQWtN
hLpN+BHaXyG4jbRdM3GllHWGqqMzATVllfisfZ18VXNhErcLD8zekl5NHvt9cc5p
L0nodKFqYWqg6wsgsdHvQrA7/d2SEIwx5JB/t/T45FA1tApIBKvS1/T3FcC8aPjH
`protect END_PROTECTED
