`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvAT+KMU9PZADAJdU1Q5LwdpA1Ydc6qg5tGHGzhHE6/yqfZIQ1oNC10BlFa7Cr8c
8CEZo5ZjJqRYlfvxSN9jkqn9SFNn7zYus9mv9rXZtX5LJZy3NM+ciBB7DQYn8nVx
hvsaAg2fKEHX1iCNQjiKdt8v1IV/C5gP4Oa3NfhV8sId5nf1ZpcE7Z/EQrQDHhY+
v+6q0cdd7c+Cx3lLGZcikhCb0lBHz2Dv8D6rMJnnOUIvLl52kUTOnzGEp/xEuFcf
5ScERMrn3EKg3J+bEcIzz2jDp3mb16oOLGpkDB3daHwzgIXyDBzVb1ITzWkfSSKJ
p+wxptDLvkxcVl7HvjEoPkjDF3whIIGPioyDWEC2C6kXpjttQ3O0/JvMsdXgiuB7
AsAEzA9Z9Y7fZmzrH3Aj4WjRO2KV+1aMN9dKkBlZeba7Ex4CI9v5sx9ocGDjnSQb
VEfCElWxvAv7Wb34AaBylt1+qC4rgpXE/Irfcqp38vOkAIoXk3OjovdYKvcJn97P
ffNlC+ERV0Qo8qDt5HZ6/kMPJyFLaMggNpcxQFShfeTMy4Q4QLDExee3BL2WII0D
pPUQN8xoBwpFwPMiAz3Dg69z0nng+aNgPTJBSFdjHMuhJSNJiiK2JtOwxjXbk0ok
t1jPVgUnDqXrJURiqWs9JTlM0k4VrMkD3RPGFcEdicWTq48/VTirvZVdeuMXhMhw
+3qMNz/wDH9QT61bXl+mtXUAw0HKXGjMCSg76BaHPwlotVoicVzObjULnvK/uwuG
jLmIzx0Rx1Fv/ZBxtc8pPpAmM/B8cmfiujdanyeUy9KnTPIF+d2vumSPwjBzu9uc
1X9Sk1M3Y/JiiRrsV6qRw+MEb+hTShBp+EwcD27D4g0O0ZahEcM3dXHhDa3CS3nu
uz/4TD0zmBGhIMGw8if+ibUJQRmA3t95JSZBZLkoEj/XWgcJPhuas97AmsNRZdP2
qdXI5ULFYAYpjU8tVphh6c3TvsrBcVJVL1AjzlL5Nx5bOP77x3vSUAeezlSi4jHZ
jJHWxUHPuauMGgJ31wG0voZDWuAN7MNGX9lWU4CgpqWOcoXCPSpj9wwFV5qX/kUD
NBpob6osMSSZfPQbpFifPn9OX29B4eh6hu7Qu64PwJz/h7CZ3eoT1kwmdvpRNbFK
+3T+we/SkKS7MGGg8f2Fy2gQuOzGVaodkuiq0y1CkbSxNUljA948QqGKil06zdB0
oA5/CUilzjhmxFEDJyecofeP0TqvtvqMvgX65s8mbc2OL4pC0DMv/xCMFC4NrjHI
72w+zbkpDiqV7YTyVzZvrAWp574OhJgNAZLum7+FdaW/XYk4kaN54Hb81K/f/M9F
Ga9VcxY72CfyvJk1Us2FMUDfyHH1pxGB1rrEBw8i5MBM8dcapQyicZzffm0LqQgb
6vGhe7Eo6GotnxfUNvlxlqZg492c14cGCHIoR2hqlU8=
`protect END_PROTECTED
