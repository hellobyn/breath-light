`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pc8vO4TFmv7UMOk7h4pM/ToKFYj0TLrTAL7c8ahOi69lb6FeCBHPsA4Ag87Z29vR
dvI9sIMA8fXCPIq4IO/lPQMsNbCer+Y1kzbA6kMxGU45FHg4ZLnk3llHVfd97jL2
4PLhtuzAmy4V3TWElec2BqyeaGrrlE/a4HOPs2dqvBV4X5IK44O8NhhVyZxjQ/zb
3R8qNlJ6UCmq//Jy4NOvtpa5WuKKiVIUrnm/r8QoMJVaKrAWuiE9PHlmTgeTjc51
dOdik9gf2m0/KlDZUtUJSbwEjr0g3Ssydu6e87z8b9yuSEjFlL0vtpWSpOIOh/JR
gaEJiog+ySgKCDkstcwe4ZoxXde6F8oBRgSzAXVmocWj3b1hJHQwbS7xp5aTGEUc
twRhyFV6Jm9rFejLQEWh1GjQLz+sUh8t+k/UQULVxF4DZOJZLx3bPEYaznZsD+Zf
/r4MiSI9LauZy8CoPRgra4EqPbtiMimpEuQLl3NbF6o/rVQU4SylpLCnr1K9akyQ
T6e0e4jiOtYOZs0UoJmTOvEcq41kCsL0RM4L0RgRZccHD110QV6jTiEV9gbuTNYs
46kRCMWD058ZvQRg3nbeMsXAsqGgIkkWUujbze6MbGlarpkDFxx2wv+nbm0FqDU5
siOeDJkv6hkY8jun6bWlmp+AqEE4VVy7j1ShdgzGYEFB3Wc8tNkarMGLB6LecBZp
1imxiAyDc2O94aVZDO1iBbbiDWC7DVcAdFw7jojJT553Ubo4RldM8GU/FRUgXEjI
qzgFVzaD2quvIeforr9AeW8UDJBGXOf76Sfm1wEAu8PIwdp3dz/v/ro/OfECqcQT
RWkU3+SFZbaI2nY1t/THKaBfW+E/fjhFSS9PTaqV4GdBopA3Vt/uM8lIpxWmH10Q
`protect END_PROTECTED
