`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R2rEhmgfn5896IySj6jdXwC2NE6SM2dQtJdRfO3662YUTUvsYEb266s9zE5Ls5ZY
dUNgdDq63u10d7XhOTpHbWbvInPN5EzTOuadkH4cyY/rQXKevHfLfentFGfswyLd
xdbl0ZO353hZAvFEZRAEL/s9sDmVDNrGVilzN4dQgSBegQDQRVNTs8AYph83jMRD
fApVO6/xw7jqcAr1/XlNN3ZEv1EcowOWIJXF+phzWZHBmAycte67jn/E9Y6pT3Zk
6rEknTP2iAaDwpdQDbymtOz2EdHNaOoiqEbGETA9aOFHjHz7hSHt76y4ha58pP1F
6keEIGrKWkFj/HRajMdqctK1e4ZeoWpvvhhJwOPhI/8EZjhiUclzkS0XN9bvafxC
WpM7FjAMgY0H850SI0dCsrfbCE88nMdYCPksAA4mhirnreZjvhYswKbtKqnrYhiE
nusDlSqJha2FfnUeFQ+9NsaEgOA8aqBcQZKiKXyJ6k+YJnA5/+LuchoC9zTeFLfw
wyasBP6XLZEJYWrkpiE+hcPWdyszhvuyr1UZP9hl+emYWqbCuIJeuRTq9S+iSkfL
nlPwd7s44P4vIvqJBjoWEIy1LaJfqKApEiv2GgqmOKGs0zwtweTVznEf2IyzXCRk
+tl4i79TZGwyzXKumu0x8kV75GZafs6DYVKmh+JbWQxYlYOvZjcZMN+5HvGOuy/o
zv0WXhLowllyBbRmRPVfOWMLQiBXiTcet8jrcrTtHy33EkOQe6NLAKDoTvSiVoux
eOG11u74oGMdhcbVTnmnGvV+iT+IRtmJMUaxhZAYyrYPvs/QnH/dFY4n8MTIYDH+
D+ucZkKtPMyDjz4llq0IQo4drNCn+qrkto8j4mYGfqnFMWtZI8n+OelnL9TF40hq
o4hGa5slmZhOek5JSa3uLw+wZzxo/41xrGpiHf779n/TkM8bbQBXnS1zI/kD6ub4
v9raPcUG4+G3FsEo66I3M/sneXFBtu3WUMaXyScsZJGe3fDWACZ7ZOrBFQKLeOJh
2tDoW9Y0mguBpsyaWkvQVmfJRjkP04TStFrnzj/xtAhf9UzMnxTnvSaejNVLSEQs
QDST5Qp8KFdatbUx1iIkEXFjoXmCTG12T3Q5J6PqpgvmP+05HBCK6sK6r8HCD19r
r3Ad0YACv+nBROdugbtyWrvrJiFImnPYXOFG7xBUSHb/fp33pQn6OiNE1phsfx9Y
s9citcAY90DHOJs/pBWVD5+ZlEko+yBWMonOosDoh+sc7+BDPTrQRZi0IngBUobN
MhdsZulfdPoHSbu8ya3LubWH8pem1ULE5l31RqC1ZULYCR1qh058h6oWAZeACKQf
cTy+caNlvvy1At3SEO650IkcIWnQOPfsmIxaoruQ3xsAZmK3vowwwDiHsrhkVkis
C51pPnSEtkMgalgpRMctmaOGF3DzRN5N7A3ZTyNK8xu0YOn/9qc7idzEEchZuPsr
jn6CPz2nmEfoTDVoKF4G7h8wSqFa1fLcJeTcGoE+loWTdkbIWOCvdXNwHebBh1I9
v4ZWYIYj3hfDKVBlfmjJ3bez/wrcMY1aLg7cWoziJxPSJVb56YnWfF6LghyAh0or
LeYwP4DgazJPZQwR0rhRvJfBvKrsQuvfYJ4SC/LQc5ESYfznrfbwiWy30aRLHxhr
0MHKmNIDMskIhRGZXlXVY0t2yR/wfZQgYbCB3Xs42+PIKMwixtoiFcLWp+7tKtzT
jEGwD1srVrio/e28Wtkz7gGdrKE+8zg8zaczNTPm8P+Y8MKMZxPRBy8rMNFEzhsp
RT0cHMGNB6f6EZXtu9wx+bAuTEBB8DaZgII3gJprna416GE5ZavTJD/b5/4KoBTC
qI9f4kOT6phMPilNRXxlHr/ALGON01SzXkKlaGdA+L774yhdgvzpMu1iBmyFwxCk
R42WjoqRxgppDMiB5aF1K1NR6YHQxHL6aR5M8s5e2pm/wnqP2/s0Y78sFF2Uh/xP
IBQvjeQ6WRkTsxtRMtxOb+hVYDpoVcZ9nuqSDmUXHm1M7+qI1SKgvsEdULAkkdzi
w2LU9oWiwoLnI28L3+X/iH3PDQMbQmgosTpjaTP63yW5oZYcIYO7P7+0Tpwg/kXB
+qSCd8jKwZG1gsBWloJMHuCus6w/r6TxnqIpKRVvLUWmbwurMioY3KuVUr1iOb8M
d0Yi9MbKsxVA6KLNs0Xq4KRk1u0PhUBaFwDiS8MxI/tdQGqhPfA6A/ooaOwa3avP
cIYjPj2LWr3gxYQeDLIl/LedrG0AllJnraDkfqgKZxtaDgS3XNuDxg8CTjrLm3eV
rNDOGLuYlkpN0AC4sqJc9gWZ5BIYTJz3hlS2+Hq7yy+q1pWAK++DICAq2U7cbbCb
JHAlIbhDqd6rcODu9t/TIR6PgDa2Wx8NOmbLp/nJ78sQR17xg2tmx8ZA7I61h5ml
T8sEOzRDu3AKeQBol+utsibr/rCEOIxszEWab8KJv26ox0esz9ueJYl/01mW164Z
xNFYSq8NwfPdY4RBzTe8u/At6hHpsfDzKL049G5FF2y1cxQc4wZxcDUJxqGlONS0
mtpegyq7P6KtQ/F11qv1lBWEDoCyxUu7xSITIbLDtRLtPllelSFLLz1JOoKM2v6v
/TypIwJHRGLFU0Pk78RTQP08+PBENCyE054vZFiALvljqTIG1TzQIKiz+TGhSiMz
KgXKBqL9nqWuu3Ydq+qPVQM1uYRzHD7dbz8nK2h0n6sgS92CKb5FOMR5uuGVozjJ
YS38kGpTKcM1AE3W4RPkDBjBTozF/nk2Ba4HujL7ZcYrTqpksx4CWXlGcxcS5CKE
xUWbQVBXz2Se027NQAcutkOE29NncKa7eItA97Fj5ZRThUZLcQwB6K/wnfPKGZua
GpLu/0Gnq5VJH63QgV2FET86VnbvvBuiFZfzOCEIHhE0LJJhE25gBSYtvXscXni2
V4Os20gTw5Ce1NyRj3h5jV1A8c4h7QUnwyVotyXjldBHWC34F8KOElWGkUGOeFDf
vCSwCTi2vKPlUSDGtR0R2FtXc508JD+FuYCzDrO5W+4g0mjV91bVjmaZqX2/TIZN
t2MGvQYCTJd4H5sgtg4CpuJ5/FmGNMifRNFWbYJe/bh3QqaaJM2E75Tmggb/ta7q
KvnrB8NRCfWKhXqv/a+LBf48uSrQ52DhIaSA2LpbmrfUTK3NSx5WNQ6GnZny6Azp
PA3O7QPY4QGraJGkba5j5POovnL0xC3eyoIpbfB42XHYwf1sVzoBiyV6Ep4cTkjS
BAsEcf0mMSwWAwXZs5YAKADCBfk00sdKdK+Yr6NudJnkitx76fUdamH4OzSQSnvJ
f6XVCKmQKg6gTIhoW4f6QvyIkgYXb+Gpz5iSKOaSq7lBXfVbFmfp06LjZn4BvXRn
f847b4x1iawOEtw1qwGu85dPKEt4wA3vnCuBSwJOIdZSWHuogT401hHjevd56Azz
usOiZiaJMErBVI8aSHixpbDEUtCYURQDPbWI2w/1isXknkZi2St5mtghTxF14nDx
qBBIq95Fnye8mVrzGD4Jc7aIdwypp5+1DuSxd54NERfq+YVmhgsP04YIHSISdveC
aWaA9WurTQBLfiqDprM1PSoYRYbJ8a3LeHNynQHH8QuIaXY69o3MVqM0plbimOf7
YlwcmJlBIvrGoUHIlf3KFICcpzmmktBFQyH8OEGCBils0DHwW+Uqd7KVpr8tY6IC
NtA2c5oiVGv/CVJHlbVokqLjuXQd/8L+vIMkjsywvOwoSRGvDxiz2zF2HWUoeujD
vpJjfbv+qpbzlgasX6OsLthA5kbCJ5k8HijSvv6EtQV6XKSJxNnTUM9lksqaw7RB
RvcahUls+KifLugG3EWgewOOA+KRCXQeuHfdSkeku8VEK0E7Q43w8t60QuuBqaFd
ZUpDn8KsxHkoyf2SPDj51OcYu0+9KK1r830Iq4k4xYmcjZqklJP+4cL12D0CTSeY
ajMZg1M90p+qGZqLIsXClasIBGLaspuWzwo1rCq7xquE9v78Qohvf96OdglPDHuD
BQ+tFudgMjuj29kTWbo5gES0h1iAb1N9S34l/4t/BXBsPRPDyq+utMW/jr/lFlwl
cDgH/14UNkzGuFcuIpmz6N3mOO17opbeg4flyCpuPamrTMNm2n3Su0ImVA9xJJge
avRoQHsGA9Zo4IkVI6QAD/ehB/gXEaaRBXYtOxbf/EzS9/YbPm0SujHV4hq6kDXp
9Z/ukkJb8g956XmI31sr9M19oILlegjDmzz5Trxk4u8ZZaVglYW5IoyioLlUfXWr
s++SsLj3sIj5MHu3YFLbRhxannoGdguTXdFhrFmH8rg+AWVBRGI0miTGjusmg68x
LtTgBXwXgvyEg9ptBPidftuJi4eoq9+97MAO/cgBF6fR1Crm63eO3xDbG8RrAWxg
LlVzNrgQrER9NA9cCXbQZ9Dj4JJqo+eOWdmyhkfSS0/VpHCSnA+TWi82eSlvfw6Y
oXUENYUFpus34irlfMamKCnC/6MPf3kdsSKNbe0DzPq1s5TyTbinDHmYN3I0rRlr
L0qFbhdn1nSOJUMQgffLtxySdkHeVDdo2pRx6AMcSYsMltspurWXwzMFgAE7IhpX
pgd53Goy1lzUERNQGombqImUfj0Q7hWSPy/l4l+5/RcyP/5ourzQB/WXgotHhtRq
QfawPNXLqyE78KsMwI9yHPT95+n+dLPQVqzST1OwBeIgaSSRcOGSBbQNksNYTwc+
6du7JR9jj3GuiHzplTy3pvwR7CnHmOkx/aTykkmujAv7F1zg4zP6zy9vPCQPQQDa
q2ACBARggqWDSxPNmUYQQ44mKrh2AIPNVaD+optdv5yqWEApN9SGSmsygTNfHesQ
GtKYUPrzA012HNapA5V6wwyBotTKTbmNfi1rxK60qTmUWX41PJi+y+4dG9Jwxjfa
2kBW3g18SXMMxxGpiKsS0sySCPErWRcWxHHZ3fYry3pmmldbkLsZVbFxmcZjwVYI
VzrHKiba+0WnMEoversg1jvYzd+MBVSt41zABtj7IuumRRtr7k0nzlMBtJi6w0rY
3SiFgXdIF4jd2VsVC7d60HLnTsLZylUXz03JeDyLrleqDGy/MvsNoaAMiTZ5r6vw
QjawHy5OqJjIBgAOoERUph4buhEoqxozXFYI0gKxkYe1DgsDFPrEoVNhe+QhPLil
VxQIjsSGH5XXKPik1PaYWNQF8BR8o8BuRRlkcjWqQ4ctuFWaN7byuHXW2ffl3AaG
WTeHPGqQRnHMXToUigRw/Hqvy/MT8IkHSlbJZagy+OshmkX7uXSPfuxygwJdorjM
OeAV1tX61BsuuVklxcf0vimLClHwjNcqTF6m+wsicEBxx99EpeS+MpaAlPtuiffM
r9yQmLdiwCYUHRLdacKBCGiyAkRpaQ89jSwqTFxOgirxxbimisL0Jtkotw3eTgeh
ylVmLn1Y6Z4fdRqcRVQcsbG18dOWTsnKUeHBFe91eAMp7/elPQWAeQq3a2iL0yuU
/DzQ/+EqoUKD80vn5ovC26YG1znpQKsbZdU1d3PtFydHoX1mkvGKUlBdd5sPSfic
dxT11Y1ut9ycFRObbksE+BtN7x1dPC6pjdaXN+ZA/QhNLDo6XcSyKwCoNmpSDCaD
UgtxjNm/PZjGQzzk3UFyuV7amkYsFjMvMPtEbmhAR9dSTbHtUIcHLIfR/qm7DlML
gBCaQdbE2mGvaYZhBEA8GprdJOZ8a/eIYygpxVEwK5XdrZ5v43Iv8A1wZQrQguUq
DNQcPL4XakkaRUeNiwq/UqPTAncciMnXe0pY4LLhP8+pDcD2JrcjpVoRBwXSTNuZ
CpGgjj4CYXlCvUqD8XNr2WIWqnO/K7aFvZWaGN1Ts0lHLtHb9B9qPIf3WRTtzTpZ
i6IghEGBxCEy1uzd+eAr/QXsnVDlLedRY3ulFq5VIUvlUvCkYlo6E3kt6w07xwE3
SGKLAmx+kTXcVYqi2+uwbp7/GnNLw5ZRpeVAk072fUkyNEuTAOyVGFe+EjfVVN9V
pKIZqAFOU65otgVJfcSqfeGQYo+Cha8WdLG1lA4x1EHUnCSKqgfzvILxNTAfpm5q
/QVIsy4fZTUVGR4amtnzeCMHA91bhsFzyWQM+kI78OY6S5gKCN599WgBXzAHodDM
eIrTtNvprQ5oVYSJb88pULx068Z6gGE7Kr0iiUUMiCKZinVR9l1Y6/NEQzYzbbR0
Z/jwo8eISH1/9y/07Gy0u7qhunx/V0QqoGuqEZHXe5Su8tw3FNp/3s8+AG6x+97T
iicYsjc4Ozda53II+O2NuJHMWrT8KosS6HAofLt/w3VyMbFkWcAdYkKrdViLIoaY
+DOeuaKjzO+FfHAv+z3FZCwH1Ra2+Gw/zNwW8G2EfpFeCVu9ZJyhCh7xbv0hDwbP
NzQ039uKUMTp2GGfk5iTeaQZJTLMLrYlN6Gz3UEghH1eLU9L9z0LQoybN/CNrr3V
RQedDVE/19Sd7hGL3Fm7sgcEY+ua8003icNodG8G+EVAYs2YocwMyII1UCDqnOTX
AaUJh8CBl571LZelPHs6coHk3upzS6pUaPAb1vR3xJpRlK2RfNK7E0Pwo01uVrrV
gqRonvc2q/nVNRwQbipu/a3szLJp3uwEhGGDcWYiaRwxFFMQNTbJmYY3IcqJotHZ
ZzPKwoY97587nfcRDNmNO3jtezl2m34BQHaizlHR8coLgzzYaYt3SmfVUs6N5KPE
rH9w32Giezl0XB7VxgZAKCx0A+yKCsRoLZIp+C93Sg6G9zvwlC/HDztFIlvj5tmf
ddTBPvdxIW5RvJ5bTU0nhKD3FFP+bClE//VGvo+yFjcHIUi/XoVXbv/ARMlzzMGX
hs/Yt/4TVrXBJeIEJvHk515cYbSqCtHsyB3hAzUpR/xwr57UG96XhbKczDUOFCxn
jD54ew92rPMaFv08ixho3MBJ+ngifU6LtxcF3qJeiqx7DhWQolRWuPD0xTZLc/6/
zAa9JuCp2ftGz+I5j2A/Xi5EEGMDwPDa+dr1k9LPel3jYXLe1hkj5iJP7VpshmMN
DupSD20n2WXhySjm5XkW5LPSJQidUiGN6LFyFQF5a9IWtjzQf2KhbyC17Ryeo00J
qx5GHrERmaPrMh/iGshy4029Ji3919wdzghR/8EgzkmQSPcIDMAmKCQYg3Jp5J8w
L7Vgi0IvPtoX1asv0jPGjmoXyA18/QUNbXxw2+KdiJnjTOJrB6Ve2MS5fSMwyyEz
wcfQAdv2tCwOLqfLxy1Fgzccptgn3lgRMOs9vR+50j9zf5mbP54tIYskVRulnr7e
K8LGlr/9t0wNLvl5OO47gBvrW1FqPAR2srA77mmwiD26uo93U/XhgBazohN/v/D8
Hsk1fx/pj59qUNEo8vln1xHrpdFpVxZvTlttj323fEno7GnirT7qHZZI4auaD917
xS+yIpoz9XGUsKS2neM1/6ZRRPEw+5sG4BJ3Js48S3oybpJWKlrjFUYIi5UMjv7z
mgtHRQzfEWCxtARSIPF8CcRA9CB+vtAmCabOd54BYl5UpbDJibA9AnR9zbwNG/SU
3zVAF79BkNBhXaTaoqg8ut93cOc+8rFAdpQaDq1QDS5GcAuWdacnXpzI2H4nCbou
UHWpxqiN+mjs7bO6dmqUvuxzi213VBzvYH3o7Fk/np27yrvYLjuUXYIZRqXaagld
zn/fXACmRtqWATravcE/od6KNJjwMUZbYS0ub5f1OOTEZy8hODR8lpVaiOuRTXQa
F4jf3RulJkcA4LHbafDOherjCj4nIpHtj/lu66tq8wgRfLbV4fYtedB6WyDtFjQc
7SPOZiy2ojJ+RmNPyNOKSOlSKHecyliKzVVO9rVC55cr7pnjsI73SZMWVBpPqF04
KbpM5Ju1CRwJJ1vZBIDqGzKUhHXpshEoulB0nSqMKy6JiptOsHb5Flaq0puP2VIb
hWEhTDyexcHthvabkCMtLu8Q5a28UXStnRLggymvR372gwScNnHmPbSrj7bQVf44
YElydgxvjVoSwpGS1IsuuHVoVBPMEqKYl+q6whVKiP5IUNALEIpcSttzqnRidGh1
5HQxj2YHQWmju0lifUb+E5ufnX5sSbqbHG5NI+qtP0y6CxJmG7FpLGdTFJhjclT8
VJbzPSc6/VCQih3mge+jCH/4fhLYnq5mSpatje+QkgVdWddIq7Z5IyQUfEPT1zao
XCeiaW+elvWZf9U1IX6x9/lSUiF312g6W6sUjnUAAb3G1J7fGOH+Am5eNdhXr9I7
pRrA6zz8oJfm5towbxEEc9mDU0SKbNgtcaYLW2ymQvm+DAKR1+//oYF938X3KjUQ
CYxYee1ye/mjjDpAkGLJ97MwQVgJJLBii7EmcXnAAS26dcZI4uccb7Zuzx3uLePi
h6aBz2CMJdcCLvacceZ2RtkRRtDX7l8Vw2sAYeaWGvgoDitwivxIe+lx3Oagm5Bl
7EEPvkGX0xEEzrSZlppK60ihGlHXanyh/i0XmAE/dcM+rqKCAnVXwCSFWumfLusF
k1gErcAfXsXJWZyzldPFsybbpDmHgADmA8vqCYGYVIJ63uuoe5r2OeSiFJsqcUNK
zH29lxdsov5MuTrZGH0lCXJkSs3G20q/DjYBSz8OfWIguZuJvsm9KQrsdEcTsmei
8jh+NoHA26zNd7xgEBLRdVNliDQOl8CNBtIxZ/ytF/bEZisEBWxXLQ0nwjBTh33p
Au0v3iYKeA3K0I8UYoX1lwQ0NAs/vc2OmnBvfrcfRw7W1n1Ebo0BNEvdTahF00re
Byt/WUqbXBWgIAy64AQiKBdDY4HFRaRtwlgijoQd0iJBsONkb80pZKHWVI8GYzsP
g+2JBr/k17Wy84swmDPBhRDqLFMBMAbA2ExZHqt8pOC9UcYGYfl4Sl0STK6Pq5cz
nNXce9EVMQfBkVimXTc82uN78QrTyYeeIlBaKMVHR80gQrvNV7NMsR5qFcDBRS/g
zaTegpuhmRRDoAYERg4gk2P5EdIF3vTbXx30rBu7s9vpmk0qzPecTZMKBss+KJO1
2NraInNAXY4sW4m3Jk7B5uocVQu+bcLHDol/gzLgtYd/bTwspicaG2MaTTJ910nY
WP+cIxm3eyXRC/L5PGGz6Ob8kFHAzKNHX2Andj1WkM9+uRP1AWpPyEXBwBjExoQ7
FC7LZGs+HgVA50H02uIT6AqhmEGE2M8a7wDnp5W9rrSgPMYM62HRchxjyPJ10Pij
mMolyQ0O9mJUo/lskkvWTVG/oF3pLEcgckbSKH9laHwRRdgdOlSAyWOj+OSTr92w
dMqBbnvpBOP/F0FUFnWgUW6wqWX9Ql8cEeQxeV4/y35yZfYyJ9fy9XTx78YEvLZD
AQ+DMquZNxaCLtRBYP1iWwZMReuFocNApuQ90oOou00CTw/vgjxFr0FH5AEgFviK
S9gl9gQDUcReVLiR0azsXa8Baq2O+6zLcTWLjkr9vg3OYkQqSw+obwC3d06gbp4b
xSp5sr2CQfaA1iBG9yCosRuZguEuvLfao+YkXqVSDshLNpCyDl7RCgwDIhCWAZpg
mhn32IN5PlDFj+E+HuAI14ivILPnin+6TODu63REjmwAs/Vql8d7MpYsxnUmwIdx
9CGX8fv5/VLqUVq6ELqk9jy883ymX6CBYKny2s+fvHkKFpvj68XPddonEINhJ2M4
`protect END_PROTECTED
