`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cU6OCSteYCtc45AmAVpQ+B0C1CcyBccqZGCu/vsVTfiPtthvCg384TELxGyhNaCC
vpqqURiuoylz3kQ5tqCEPQjBbgZuq/TgSb5sI/h1e9eMZz28l4DAIs4EWePAu+1h
tfoOUtvcBeGVNPJY073KOgCXYIV3uGBMgkVWsF1FHcFwA5CsHjqzRp9yGMDjHeGz
F706RmC3Mm4JeEfW4/tST9GUET9flsRHNnEjcwXsmjfg477Tu9aR8zWDie2eL/Om
JLpNL4Qxq4WjRfeMwUO8hw8I6Lsw3HxNpjxpWBYpNTtiQNjGwN/AgpjARZ79JiTv
u6VqcKmzHbJcNNcLlCLvaQHLXarrpPrpNQu5nm5gaEX5jQwztE2tlv1Tj6UUjodr
sj0jhNpMyFsxY5oDdKC5q3sCFoFnpsrH/tbq9/+uAKVyw9kTQkz6eVpcJ89bgkHV
usniALc+M2R4Vx/CDL0nUN13/16+hIkzCtmSx675cWQ=
`protect END_PROTECTED
