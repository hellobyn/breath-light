`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABF0Y17fwRJ96KJaxOWk1QVyKf/ETlc+JSkQpMWPpOFJGbfpcS4fi3dE34uZQACb
02VaFQk0j7th+vDj9MhKDq1iEdO/qCO/F6o+nXBKVcnLhoyY6BkAYOBrhddSyLGV
JGdjyhE3szlHghS3mi5Ofdf6Wi3PD8NPXswcZjNlYinORGQGVTtz5RhmLs+w3rWQ
y3XR1gK5xH5J8uKCFM5jbYLbXbabhCo+nmn7KIodM1v1OTCc11AkOo/JmhW7/PCb
mLUYtJCLDNF9RG23pb6SycgYnXzsyxIAgVJA02saL7DOt46aYIlQOzoLMTOIRvur
PB9J9wfPijsQU7iALqBm+73SsWnUl/UPN+xqHLmAXQLh1ahJlJbhM72IesXj4c09
Np13Y7gsfT6yeoy1I43BzJ7IqaTZb+qcXucYfmPVH6xgyuSOU6oifdmnHFbUFEMR
ff6adAMoPMYD3YAM22U/6HEeqgD4gw47AyorFzi8Obo0nMTT0NzdHkDi7NTe/Imz
YqWf0uKxoIcuUr8CxEU9V8e0hnyv40jazP55ziNRZVq0KERjQDzUGapd7wX1lxVm
BAZQtERBSbX0W3lVA2JRhndH7O5siSqpX9tV5kT/UvNj0ozUMvt35BOOjQxjSdfG
4oAg9qDT52XoiQpy7zvME8reasKPYQZATTnpzllMpSeaIgTN8jT2UUS9StXZUe7M
B3vVJ4hxFfGitev505orXz1U0nyIU3BlXW/4YmeOWuYJkG5jMUgMGIKBnO+jeMtl
cr91XrMdZN7pjffwtsq80FODv8terLdXJoW9Fs6Eg3tyz7bIvjDrHg8aRQEv1E81
2czpt8nXGols6GRYW/AFXqHBhOzls2JhPv941pjgCQoo9eNDYSvze4EArZidA3x9
7teuesphU8nJ15U82QxXkdErDJIWEQ8qVSQA6AKMPqyFIN2tdzEEqKPSNDm1YAdu
wK4+2fnLVz5Ioiifa2fGHb+Pl6ss1luUpaiYkzrzzaHncOXZBVpihxGA9UMyNMxv
xcxPfCnQg1PVVGOWQ2wd4n1N3B2F2Gc7m6zbOgCOELaksWouF+kQOPZc5cxdFS1G
MHzBKrzEHu4+Je5FHARf5LYO6k/X3gdpYzpU9jRwv+iB7D3BnB7bIOjfmts+pQeL
J7Ki9APb9LKGBea9ha0HnOXSAyNfXsi246UC4bWfzqvaDk2NBmAKTvCq8m005HHT
WgEX79tRFQhPYBfvmuToHdrPbgTRD+bAaQN4ZWWN4zDpFdL79BpIGTQfT4xIrWad
QlcLjzLVqQPbRERF8IOZROcSVqoyCW7yJUN+ARSXIm+ryyfDDuR7TwoidEi7NALb
+ZOCMA2VgvPdce7TlVotz1Czq9QORbdEGTnj9CaB3zMaEri23j9hYNwYnMBuDa7G
H3EzRm/LCSXXxtMkl+zRb/HsoyTTeE1oWNpGscpKl4oP+JOxHY9rIWCl2GTQiviN
Di0oiXEsN9yi8UD6ljxP1W2xnObMT5HRp2bgtaoGtm9mtTlinfxg0h2b5t47d7Gd
wIGbtvClPfjuOmWVwbMI5GliigF2ZtYy4Alvqj6nxmPvt7T7hiI7P1TB2ToRAxVW
T1gw/bSVB6Ljn29GmISSAXCMYsrkPR7kCFtm48FZLs+y9cmrrTzyDkGZdN9To35w
HM08nUNElgPU3xwz4DTcC0jlGuMyEUySA7fNyWUAVAhNzctmULBzkh21tYj+UkUi
N9Ycf3cfnE7patru6g8bZiTxyUkTU0EsyjUtIaQdlOlVWk3Fjp/GhCeV4DWo4Ikw
3fnPreXXHfij2jjv5vOUPV3xfdMFPrwqQ16ARFTaNILVfA1hpgQyUlV0NM/N+8hh
aCQfflHKPim+voH3ngc5oh8AGzUp84kaQgPkuq+uvOXGsC/hAplXYSkuvUKRFGE/
kxTZWWSQpDSkTLQA9cOHqrH+xVe9jFOH+kaBSCeaxPM5fWFjLJOqFDQAEfD6+VCi
JmbBB3YJFlldrrLXDeOu8BTKWaExiB4SZG5pk6B/UIHI1aT1EsRuSdHtivxt+YRb
pjKYIzPlif+c9Npc2jW7u4FX0R2dJTrxXdPtGAXZXoZ09iWqpXBK94w7VGA55Rdi
j5dQqfqXYXnPziIgja+QnSHP+e0ueMIUESKtxtfTZjltlUUcFKxUHpwKHuXvBiR9
NpaO2utuR2yEeHti2mEZdSJuRR0nFc7wtmlfpU0vcEg1owMwB9JjkZR+BwmJgGoo
bLNmASxGXdfFYeRlQJdGFP+bClH5W5ierLYLSw+8KO0quMsLktt9krBNnSacx6OU
+1CJOeF1eme6u1NB/rBkvYuirg8Ni7TxLSYKJ+qaN/5Ls2DnbZ52Xv+pX/7SsYop
qf7p1fWu6xiG4xKsh2ZJEjW6Bny3zijd3JklRILkiILvMp9YfZraZ59ID8SQLrO1
112969riWmToLDxWdQTYfRGXh8qyNGhgL2qEbEIfM1WBltavJMas8KEsjSV8AT6A
2pVb6myBLV7FmkgbQRuK+bk+LcAnZdmaiejTLCHSn4ZiRsw6ELL5iZa0bwIRTDi7
yH1ZAUZH+kE7+EKDu+kZWPTbZyvPT0qLycQHh6LJjueZKb6rCtdsD1NYWtr2oLvK
dtDfSBJpq2tJB8Twt2aHF3QV7MZZzvvsYNU7BYtSO0kxscqS6jORo1Ir9+pSMTBx
aNb8xV+i2rqOEP4h8t9if9N8UXnc0id3Ej0iGSU5IorLPb5IC1k/M0OKHN6vVTnj
/TrmAXm7NzCTePsIPIaOtYbhE3I6dakdAMhhBS+uMvcGf/qR4/L0PZXlJY5UEtmy
1nxd+BTID/lczyKQfgDzDH2D1tefebjyST4Ouyj6CuhF4v94aii77brBB39sk5Nx
E/mgUIrvI5Zkrdp65SoFHm4UbKwdIi+oj4LD5p/BI15ZXdmScVXfHrEFNIou/8Ef
Sa2aYdt3/EUC5Xsd0sAaCZWDKIUX+U3VPKlMSKLRTI9QdKxuAyj93Zk/QpDcwQGM
AGx9ewFje3prjc75P5PYXTY1pgtaKZMAI5cdw+XkNnTNeMR6P2OpBuB5Fk1zmeXT
55rV64gCLHoGOCzTojDSWOhOd2cc3VLkC9+mD/nBtN7z1eM4eifGbhWe7hpKD2fg
3ny6G+WOusUrai5IrU+NPvIKFYEo1dYDnoERN74u9rodAERtDCkTafEdF1m5QRfK
inDYbucVy1AJoTt+htQBMcYbDYyRS46pT8VLnTEw4Q/BIatImYtgtgd8wbsf3nBS
cTPHBzSeOB0TPHR4GcMSC2TP9vrXAxcu5Pgll2aoAG/Y/i7oajPl4nKRvbMwJAMp
tspXSxFAUWsr8slMQvERrhCzd+4OgWDvuSEdbZzar3luPtf2YRWQnyEFad8rsvcl
5HNm5c1sqnjW+eJPfF/Tm2P0H57h2PxTBNpPGVieHY1HyCWSGTmLji6mWHAMgCyd
ddTkTfcziT8r4HndGHOJWc96K4fI5Ih6R0+/vbM+0VdEAD/7MqYZb1voxRFZaobF
P+Dotxk2BygxAVcdsl6SwMsCh5D+9YQ40kv5ob7YfcRpCySVIBqCfKBi4eZPIBly
68xW+hStaBBwOGSKCXkShAlWe3hfqPhHKoPFQKlPiuyIToCD5h8THBPaZMAfesYT
w90e206hmtETHJVjIzwAlBb3LERtp+slHypVFRJkxW6HhP5hxqH35lVM4UXNxMHe
K1rg0lxGa1GWsXsk3niZkWuytNcOip7okFmFPZJyFUfu7n3CLoGAFAf3TsBxVTTO
bVR2kRYRoWxStre61+N2dLI8rh0fr601XTvGTgdMe/4wRHDPdwF4n5YYCDwoi4G9
Sy0fFDvJiDG2gWWMWM9uOmc5EvN02G/+snAwcQAUjsZ0DSynYR6cwo5wwg3L3xNN
Xtx2ch//VYKMkgxQAoCKAf3MaTyBVK80fDJXhIunffZTOimDOasXQXts3HHT0n2V
o5aUi+LjlaeeBdapVYRmZpPQSR2oOT5bNvdgCYvJse2naoMeaYPCemtyuaOl9vj1
tCFk8XfaLDOGf8liIGf46+6IPfSOmLNh41Bbnep/h78h6xD/rTSYI84x0jMPyGr/
9eCA0wGXG31tO2awKpQUIDpY62jOG+vt/AMm+16zech1kDgJwbYU8Sv85lhrJ56h
ONMa80WkyEh8OoZONyXLRBdYCaI2Bk3xEX2IDMg22rGPJSl7gpGUihkg1TNmtHyc
kKVV19vV7wC0+Xh/f4VrIJcyYVgx9mFPIGBeiY9s1e/4hJuNNUDIYDVIpf9W0vQ5
LtHY9Q1sgd253qQbHE52xVnUvgOkH2VByMezEVnqUu0kf+70mUxfXwSVtC2egCIY
/FwJjENasKxbya3fV4s8S3bI0KFWTfmkwXWAakGXIhL6TVQ35rbpTQWH6fk50avb
4iHGDDaPMqn8qCyQxgqsxOg2/627w0t+m6szsT2zWyLX8zLdylAvVSI5rcA0Bvoj
FRv1OlMNwrj2EkhJxnqbcYFmF5dt1CQIoOmLYEcmXr9W4GnMonTbT3b0yg2FJdVw
aRxaCS3YsFrLtxrLugwu8j9hoLM425oyfr8zXvpTPDPUsFOFuehVZ6fNUljcspaA
ezKVdhIfUhtCemFaC3JBSlSlKEQ2aooCKQ8sn9ROJMSvt1GVPnEh07NYPdO+Be9k
kW8lmldEPRbKg0lqtdz0UEQqsfJXY6pA3fDc/OZX6KT2jITHEa+hp4Yad3LVvZMs
iYeS3go4T/b7s3buOs1T72FUX4KiQo3ZvsMWX0jqUtjrUkvLimJM2YOZirWhEBwp
kwGNFzNpHnbXHRBfRMAHd9Vcm/1zZ4fUFC5McwT7GXT/vus3FDkGoEpzvXq5a9+B
GOWwTctRafa5XVlHxmP/C5+KnRa01ktF0jHQNWHhWdzSqyEpjevFjaySFwj8gY4A
A2UH82iNVtiQlcMneSV0ZSVpZAYF8vE4C0GNAd7yThK1wPuBBB3kWbQpjaYhMXUv
Jbv0/dSDjjocUGXLGSU09bExz3bH6gb3a22ZO5kA7Q/NbM4/Uow0CKkfw9R85yqT
CVI60m5jIVk9QltqDp6dW3VDR57Y7+kwvu90zkhHPPe6RCPDxl9IHg9Yu3h/Rp2x
qQjO5s0TFl9a7nPuXBgSUMGgsqMm1rAemznLaF130T5pZEIFjwbJBVslKaapqoKH
WB3Q71mmdzMKc+2qM/H5BtFBN9TqG/revBy9lx1wXtIlSMfwpuAFu6ldtMeow9BE
z+ue+i2qaV08puFQp5oc7gtXF6fBpZCO6uJyoQoOc8lCw25DHo4kTMHSz7EoPlJl
XZxDgy2F979laoAEUhIukeZzgaoRuaOxi1Xw3KLD8Pxyzml8RnTmDPTEzU7LESz/
fNsFVXZXvF5pK258XA7gGCHCamVSeDJ8CdvuXvRDv7yPDkJfnSAlAaoCEe1PfV30
RI7TlEVRzSS+1xEdUNX6Bh8RR2sMg8vjxA2KP72skG7oo9+h9SiHqc1fc78SS3Km
LCLKJpTJvp9RZX3ICyWz9Vc1bgx7XHMkfIg8opc3rs4DES3PHZ3QpBGSwyTSLkkX
tFqb7pmiHQsSfZCkWOdu5XQ1EqYjqNwD6DWd3smwQAyg08P0hLnqs3p2A/RXUot1
BXFkpOhJlStk96BvoKtBp/uX/O5ms/VNvBnM1K4ZyNgzWcqbInG0yHNaylFu33qH
dw6aHeuaJrKnL/coDQzyq3/60c6ojFOXrYQs0mIA1lcBBSEqu2ADibFsEryLk6QW
CqrWNpz32JhEaXReLdHGnNWBtJ4/2jI1sd20Y0ye5rZDLUcP/m7gBqxQnqtkewQl
kgw3eOstK54tyKMKliuWjOEHuwuIQ09+vHRZNQwCro/uqSjlL3R3bejBy6HGylkD
tazJPBtXX+BB0W2ljfVFD+Qa7JJYNoZf+flJAXW07+f74wefS+442Ux1on7GkheR
Av9JZD7RctVQywo5uCFt6j0MyOvApiTc+JM67EBN8uMf4l0ZbBuXVEgvcFh3k8HP
3YpcqQrAyJdxiE5izZA0Gqil054x0GPvEtkEqz3VKN90UNiRt0jLyZwi2LmkqOsc
iHHN3Slh6KzhPZfVx+u2R0yGOAGOUh4ui9PNG1Zz+iEOAnPj9O/0NiKxgxlGO5pV
cqTHxRXWm4mOMv0cG78FOiXMcudPuxPzXjUi8yBZ8HuI+ZTCH17qJnDpfvaJummD
poTHsS9uTfgDFQuWCGPzwY3uGexguwOCyoByTtN89acvn3d8XqwWFF4gWPtiYIXM
V0iOC9QvUjM0gpelRGN3Dqv512CtoZrQvhfI0LnznA/SSQsU86b/hP6KEHXgznXQ
64dlltp0ZaMrjohDhi+/HuZb08qJTnbrT0fqRuYW8Z4Ka3vVTPcTuQBaeE9owknq
PxkKBn6FnvlSMLGQxMBBQzoJtRKTzJQp5XClon8bk1F9bFMrVjxv/zcEJoiRPuIR
r4fkHjhUuxyxGt6hgeJ8f3ksd+ESvj9slVPoIeoRCP1Vx9pX644x9qxhjd6wx3kw
G9tRvB76L6zn+aH0BngvW49sCiy8BFYEJPDh7D9XLhBxTCbgH6H/P1+HoXyqH78b
Mvk8akdpNBpmI6HCXega6J8hUms0Mtwi+Q7iw5aQODjJnXENVIh1+7VQb4Kmxsb3
l2kPh6BKuvMd2LHF8XSkm2Cz8a8Cz5TxGYokCpSyztWdUWlOfn8wzA9FbwWV8OB5
JcXhN7g/neCUyqWMihDGPVN1pbY9T3lncgJQhQ2fr6IxPQk4HjRNqd8bC68ZOZkr
8VMc0+qPhoI4LXPOx8AbL+VM2LfPjGSPVpqKh+lyZEyEEphqKvgd4dOyCOyqCfn6
bDusoGhTeK9npkddig9UHH0DnJwadKARsk8jLp6O9cGzpcFfzqfwrLOi0PupWRWE
PBcZCL7T6CBQHgDrYybL6eFrV+jyyYLUp8bRhA6N/xilFlLV+mYzBA7tQFlFWS9k
j9t84dwyVfUmEz/KAHEQqB4CYCrgNFNQM83C/ZBvYUDZAIMeJ5Qzl8xFMmNcvwjh
GNk+cT43F3/h6zgx9YkNijo5HftESJGkIWPoEJ0ulBtTmZ6Kl7kl+bRZ6biBDW/M
9XOd1RTXCL+LhHXjOm48efLfqUj+1D5KI8ZNMsXo/p63X28klQfGX6IMwat1kYZw
668kv2ooOiIT/E0ldYtXi0fpzU845gQe/6b302mE0RSJ5sA0S8hkMmYuX/d9OrRb
wiozYaXJa497Y5CvXmRU04xjL9wIQKpjpuAFglAUotmEqehNEKL15NLY7k4B3Gry
rjmjak0vAK4nZ/Vop7ZTLzyZivetHP+60SahCRYL12eqmz7UFgL+jSiGMV5eSg3k
atraIrUiYNYgECq5rLrDlPzIcsJ2MaoOfelIeRYSFhbDLcbDZr6J7Ug4kthQmc/K
iBKrHvKPbFYRfghDadiIsrl/iayS3YTxsbQ3ohpKYPzJ1A+pyx5LyDofonsiVYxZ
VBpPdDWz/+Qqd92O+LcQFlzWkp4iasVYfoVfCySZdInbWD1J4Z3TgMLRhXKDIKXZ
wk1UuQvdcNUTfQtl13ykVM+inBWX7D14yUU3IcVxtf7sdKWsu7vFr1JJerhRsV0w
+oZrbZ3c9soNjeaKV8d8nP3EcdNseVfV/B5ZpkWpVd2Lf9sLstb6BJx8JT6mht2b
qLmW9TM10FOlCbADbcLyaaG+zIMu54AoL99gQsGmxFpwCjtamxFpNXZ4UOfhVXtV
l3rjKmI+DxVWHP9ne1bLz3oJybfHTDY/prtOx0IqgxeWxBHmHHnK4onQaMAhnkks
KrWsTYQ+xTD81pApuOxIzydF0wGTnnLBajfsfWoVS2UQ1c/Uca4Yc8KRLt4eQdz/
79MNenwaeUw+6x0MAzq+TyIYIiurR4NAF8vgaLpNUTxrqh1QvLYSUI0E/mltnFO3
c0TlQYwoN/dlAg3HYjd5chS5L+EDegUxT4atlrkozTsHhH69eWNrsEJhCCL8jgT6
NGUCzfw13l7k6xUrtheOnxflH8XAuzkXPBnchi3vJyV/+6W1axqXplOth8XClfdV
+WU8fDPS807yC7HKzeKAVd5avvDaZolH6q8uLmG1FuBiUiqIK7nh1NLijQVaOOwi
HMQ7n1ZA8QSfVcz7o49O+VfVyiJFXIhdlg7aCIlHqCleMDur034NbSgR7b9eTrSn
X/5G0yiPTYkLqs8gXi3hMDuIO3nIr/pv04IMrGOBwZlVPBuHe/SV8sv+Nh/lEryt
ZtdQv8TFZIfACxZFJ0/LYyZcjzKbONO0Z3Ew9pH5oYDELH+at61hy60WeG8+HDjt
9loVq/zVTx7vo2L45aa7zRBXKw/T7b7UzC/FxgxOlT8K02HSB/xb7cWRIbZFpwuJ
axSOwYfGPyGPImFYSWcJPARJyz061Pp4RQernxUIKD4c6+ddOqHtJX2t8z29vIKT
LphtSKNIyNlfrn3HpDGqb6p7H4FQ58tXssfdZixrUWPtRDAZb4mI6/kP3xk7wv2h
tL+4mAJrDqPkUzO0HBReT6NZGAZSvSg77mZwkC/SN/RnJMuQWTff+8ndnoqwB7+W
ktxmW3JhuqSr/jQc8fhR2Q4UMNIM+Ap1UCYKT0ncRSk5ATPmkH3/rGjUE9HrxYhb
HoLwN3kYh01wSS8Q1pz/cmOTZuGujBn9/f6Xwj/AvF51FDAUREGJk0PNMZks7etK
lw8w0hW2UHxfZxMGUXRemEBsp2udOoEin+rK6vtCVdnE9N5Wp03mJ7OCE2lDwLYE
LSPkz5QlUtIz77S2jGr9j+dDTgAo/O7e2tuw7y8UsVsdJGr7ZN08ulwiZBFP8AHd
pfB251+X91K+XFG9VMJohQYyPBj+y6kDjXtIYJ/Z3vBia7ABdrnSD5/puIoghw5R
WzPADWGsKnz5oFCL94uAOJ39egSZoeL8FAEGnTr+u7ftgpMnvABKV+JIcVW8TYLO
A1mITqZO/yIXINfwYHkfXS1HvM2X+JM2xiyYTbNglAqldwgVosI4n/sRVzProh+F
AV+zn1z52aDtVz9l19lzC8j90ojifNviUIBiG2dctTW27SArYHTsr7DESFdrAtGv
QjYCU4CH66TKic8p4LGBXRbSITFRzkD5AgUofQ8+L/2O6UGuo870iEFKHXJ1cmC1
VCOrgulWcwSBFwpfZe1+z8H92e+cOc7NFjQmR1ApledWb4pOku9UoTY8zmFKDlTV
JKoBMZRVzy3ld7MDgPIW5gqXf2R0WeCy5HBPSUo8FZdaOkD/Q9w42q8pTcNT1w0E
GemDecY/VLSikZgJ3pB9GefMfNaRbBiPRKhVd9G56VMC8FRaLox57W9PYcHHuPOt
fUNZigI1WtVUUl3YhCRryv3opa2PnyqfKGcoQ2oFt1uqrOqn5PYwJuGdbsv+eJE+
z/yESJSs1PmlFXEc+Nk0Qd9iI61mPwVZmr5viCNxmN9vCr2LpDvw8X7+5+n8sDS/
OGT/vRHPE2X7DaCv3Sbs7IS18lX50rbmfFUAmOHD6j6GPDToRGZURw2SNJwWLpDt
FF5LOmCnTEo72uqPe1bbWs20M4OdIXAv/7MMTbb4V2QBCjJErOlqZL3oCGPb6Xzr
rW8mT7lTFL/AZTvxl6mkcX3rQcnBC9EfnlEsRZvbevvbwCszrKZuQ7jgtOfmjJI3
IxbijHcqAjU5qERSZNzPA/vveqd8kQJXiK3kCat+VyFIX90JYv+FdQjkVVRM1EnR
7rpQv9BjfYTeA8kZoCH825WKEJPe0LDhnI3kTBLfc7nNqgubJ5LljUL424ruJFOW
MLAbr5vzNyRHK32HMaJhldrTkDuIGN/IbEd85H/1PifJrYzPNsu8I1CvIwsMBdDK
jVJ04rAkP+kBqBj7ArlGaPdzS24VgMTL+rlEeeC8zWbv04GK9ozzBCYPQW/8xEyu
8nX/ykgNyzYKG0dHstfjjVfjOwTlgjrAw2Ix9hi2jo+Z1FKTc7ufDklC4fBFmXiJ
WFRBWGpcBRoNfBaEt2+s0cxe83Cf70CB1VGspEgw/tBPTukU73tXqrcq7n5NrzyP
pZtjV5WsHa7yPNjgCjT+JMQ/zkKWqyeDa7LRbA6mikjBkzv5PYKV0HoST4Sv0UrQ
TmLhVoMW77Vq9Xbf1CBp2la9WVPA4OPwGvDpMiDOkLfwdbX1nGnrySMFUNP3OiGa
/kk4M7Uhby8lmUJ7CT7+kiwHgowryKUOPP0naaQl4Q7KrsbKV3CAww4l9hjJiEIh
4LLFlNQsGmtWP6tB7SgPcrAo0wPyX+3IPHcHzlHWxM7ALEFAPn+HwzGFnZ/v2iQv
HnRL9Ay7E22MiVE18V8g3o/EDUdWBH5AJwjKLdWPIr7sOx/HaDgmgMLneSx4yTWv
UXMpr1R9GQog4x0SnBFFnhU+k3i6onl8herrcEst+yWv5XysZZZsNseH3LWuRBWZ
jMeLtc4vSAI/hdj9/pP2uhseY/3f2jjEoWtK0ObWC2H5T/6slpptCQCfsswpp/FV
ZImdov/gkp1mx+DyVo4uaNQpEH7SJ6k8lsh+2ByHwZdeSK5jJm08U+2vY4I+mf95
y8no+DahKfwDo12ycNdvmWi8VrOHw1mkpXpsZAaZuWXuU8Oam/vdpm1+PnytWq1i
2MAkJiguxU77GsWPgR0OIjkln7qYpWJ72CrZ/eD3MMU3MP4HQiXk0Ih71n5mGN/l
TKWJnNGBVsVbswzmqGi6LQQyhtg5AY9OAJB+2yG/bKzCheXVc0be5WJYYpFyKXoz
2Sqr1B7G8Obq4QVrFShSGWrrt/JYtsbo5NrhMFt/P7qRvIMyMyEaQI0D3SGcM9G3
cecXGvRKFUx5v3yyKUOGG6uwoPGWQ40UgPxrtCC3nkk9lPpdDYHcFdZtQhzbhBGU
Du2BfLAikpjHMFqN8DNcBRJUWN2yvmXnlxbp93rxlRpCT+Gc16SY1dU7U8sWmRIL
B/zfefqdSwZFkVVh48XxdVTqOUqkAd69Nhms1tqB+PtvKo5mtWvBp2teScoMhhgI
8di7AU0lyZeH4dfzsJ4GqYbYRONhsdzkikbE8oq0fRuR5xHxxz1hzxByS7qIKIO1
RRSNk+bB85zggtWWh14+mHyOdHN0Ra3sQEGgeQLJ4YgMqYsAfCeE4pLatLNAmEkM
mEYjD7eeNMfZVqJo1hinJehHx1VFlin3G3BQ1YIU8KdTIZ+sk9TmTAmPo6PThE64
Bpz50TPl6w5GIJNF05KlJgbik0y6XOJWfZIICzlwosgDOIGPbpTo7llTShkijRwA
JcD1HhbopJ3Fwz9lfI1mV5/DDPPksSewP5+6YyXc+hqh6g8oXN7XLO1+CihdgYNE
TNNdnld1TR1/ADWVDPwOYMv4YqNSjFasJ4MiTATEH3c9jy42gd/TewICRJRPRtai
MKUF93ljivsii0Rj6D2DCmIIWF2XAzXXpf0dfUw54wkIArFZYdHwR1kZVEGIrx4O
PHHr2AtDKTYdCuQmKJ8NmZYwIk69wXYJErPh1uSfWh8DWkLiYgRmWNHHmEc6coTk
EQmJNCUWLj+mmzu91ME3aa7VRO9zuV339R98wmo90pbfE2kSa4i2J6Sf2f4bgYNa
2hUjZv79WskEH+3+u4+PvroRAh17tlMOuN1ropijtBOud0DZNyL2pAxlJqCRWjrT
t5goVxXsD0eOhQSJRH5uOj8+ZGY7WkaPHWC3a7uZ02Sc77CxBRM+BR3gBVTFbgM8
cISixw3gGRWnkOpB1tKhjp3KECLaVdIQJbrFtkoPeHq1mpb6CIkMQ412Yoh+7lsP
3i21iq8eypVd0pq/fPX+nL63LL92Q2NI8r5fNoHgvyjtXhA5Cl7ckBNscTVGvI37
FQ/OAjOVEBYg0hOXULv2JqY3qFgvGaoQtU1SMc8mZDxerBM85ZzDiZL8qmci+d7j
EqDGvkrCgpzvli19eHYUoRW05F05Saqt/8Ro3orgXAKHcf3v99hnW9zLYPx7UZVZ
w/SausM8mVOOx05/Eyb/GIiOEI3n3EkfqiIHSGupKesS1PlSpn96rr477tfTIg8N
pw6PSg9xU0cpr16mAP0m1RoWeYWlyWRxWAkI/FBofGzfw+jYCHuxJnn4yJPr7v8m
YQd/7W6cpiHniNfjKLJyJZbY11pjdZ8kccKrJpNkuswgyBFhwtf/e6btxwnolLHM
D3uwoIAvkgfvXBdf6JKd2AVN6/+zl9TODvzCkLec0hxQyyZ+BCWTdm3KueVTBPZl
B2byJ4Pp7pPp0DMbLbyexwXF/qPmUCNgin+GC59M3AVuArtGG6DHHsv/VGVC7SAM
3BrQDZVMFevdF4MLSX1e9l7Umrq0sr4I3KZoB2jHfg+vxgX9uNVyjcN+ZM6L0sdy
YJSHkfzV1oH2hyknpn8Xdg+gp0o/YEbRRt0gRRqxPQXa4yeTknj75WlMbYRWRtjE
kP3IHXgD+uTfXHGlSuPhKD7MMwXUdpsjKhKjQYXjyxQjqYREhtpZoZF0MQTPGurA
KQ9bmClQDOSctrRRAU7Dp62BIAshXPndVJYbOITPUgttatcKE686qG30D6Ku0uwc
kTRLlg6+PZVY++rodVv2DgCaoy3CxzAePcsq0ZZX2sTfqZl1g8ms4lBXbmemG2k2
2AkR65ewQ7c8F7IutRPThetKLHbtdXIQDUKLIP5qp//LrttmO8cFiwf1HL9JygMc
DKq8K/RShSwTX94BF7CuX+8JuWNDKTQxCwfxm6VLL8XpRpOYQDIHFvBIP5K45FkT
xmSBOmKsQmlvHE7R2tv3T0temiUV9DDm+6xJ3J8n1PfOISKVLz5gdBTrewfzeR5S
U6++/xWZAY1DtyfrSH21uwOqz+GHOld0LwxLPPHVB9Nkuqa5Gwiiu2v7gfppemaB
JpfTCYXuDnNp+ZZ3rIBLB3cuieHXItgcoZPNGGhKMEpTNp1q0jpUkFGslgVQE7/C
/9S2Sd5FqLLXWW2GfN58LD+Wp6zIB65+E05jYskjbguw/s127s2tfppBF88rrpK0
PpHB8Mi0eXEDoxzzO+CJD3n4AFkEsHu62Jo85XK46/E8bt6Au3M3hzpjyOIV7ewm
aTbOJnwEFELwpBokQEsmdEPXKKv5TQalnJWTvoxpe+wn91FdKnzztGSNubeyKXvn
ZWrpbOd/dpS5VzH7KTrl3GHiy9Fjct9v+SXFQV9dLHslHo5BA5c6LRSPi/n8hMT6
9oQdFMaQ10cvVdv2N1/AtZKeMEWNA8y7ggSiTod8mxlKHWNQLJ4QK5f8t2vUu4HJ
dBcWnpO8HSLC/M6U88irLuPRprbVGWrDhvCnL0b2hVpbU8Gks7EQcJXNZrXM7puJ
ZHN6ON4Wnf84gYlgSW22hGOv7SCRjsCAC86pwWvH5uANxaWyS/X9Zzhoe60brNvA
33Lr/N4+NFm19PGDSR4JL8R9TYANBq4WGYJMjWaYNQuDf9W9WV3GMmkIN0GTw3CN
Ej5kaGiVuMjnsxxuNzOzWH0wW+E5tBCTv0yZHkezso71Ym3LJ3EY+z5XTwf4wDk9
FV1Art0Ux2Ukngf7pMMuutc549xLQnaB4v5GwhMLtjEFXmyS2JuZ8Bv5cJu8v8Z1
zek2eKFBXkZNfqRG6g48RTqiuYJ0tQraSEjSMrKb9iORPFvKcKepwJa6RgRiY45k
EutmQVtbzSLfyXicbozNKwIo9zTMjmubJxcDr/X9hSgnXzSco2YjSK16jZY/iFby
2sT7qLtXa/G7Xg6qrcmWNulrhoB2C31hidB9CJf6Ww1PJuNqBLI5Us7axUpFpvfN
wXUQXS7jxcgODILcbV3QZsSd2UZrOwDclZ1flCsOUf3IFktdn1DGPhBdiLRYcBoa
GMJm+Xf9eCk/LyvvvFrTgnrPA4KmwYgejouHZHKyP7pQmXpKFE8uDnw5mdZwpRiv
NNyrdpICDzMeb6cZKnbyxSPQhz6bjedK1JnV9+gKH4av9+VdI4W88XtK1LM/RnSw
MbQyYAU1uBrdCD0kSFycG5uEzo9ndMC+S1szIDi8JEIaFgEjYjZG2pEjegRU3rb5
aylNGZevUBUlH729Y+zxngM/0VMsFbMpzWquuHWyR0WU9FTAzbPMntjB07D9rDs5
ABuqS7Pqfe+A9I/pUZC8kcX4RDfiIdBq9pRWDMkDiY+t6n0bEEaw7FZQKLUwTzIU
vprZKIC8+UgFUdW2K7N9Pzg3LNQUuE24AoxCkJRa+PoAY4FjTY9rfH0EGe0ggR+A
rPlD4tD49LHr+RI3ztWE8Yp6nVSJvBGp9Rpa1mQzSRPCNSc6jfFi2PnfI/rRT5ZH
0ntTW4RLozXMaUMd7AQvGGPjOxzbRYJ3zEhTIt25k485TyMC4B7SD8Z02CR9tsEG
VGqfrH/LN8Pm3Bi2zfUeUndEG6Oao6cbBCZJ5fXDtksGMXRwmHCB3xu2s+WzPmsN
zCJQG41cXf4iCqOTLP6/Yk70YGyUGcfvbN0NAICTM3XrV4lOGDILk+sleVNQH0Vl
SjD6964IHWgN/cRdgR2jTLCm1CMUBn/vDs8alRxZeMJgb4UNlH2aDb8kNFF14iZ3
Vo5jphJyCSugUxDU3fFCLAXnAT9lJ2Rp0YiaM+E/B5eYSV4w1frhPK4NcDdDgWph
i3blmA7eCCMoIU1TFqWEdbaeVBn+voXawXear9fCKRoSqUwjHBbcqd5WU0i83YrA
889QJaktgPbT4GOJh7Q3O9GYqww5wulhAAoniMeQlAyckBLMu/8H+lXco3TkYFne
GkrW0h/uF2gvNSf3wrPx9c49DRNXG2fBpW86FASNHG5Zmo3XIdQltxZybhPyjd7L
L53cbOBsP7azmfKiReojijRIgVnZGHyaUWrOazcTMuoL4DsLFrypKloq2a88y1mJ
98frcX4QEOmagj/YO6/H39AYiObbB8ckESEVQ4eTBi3u2ZTc80TI9SCIh66AoWfD
n7R5v70j3wtA1s5DsIABs0ZcT4towGutqumM4NVkBr2m3t68jUthZl3JZUHOsNxf
N41rWS6SwWeC/BLBD3S4spLSYd5G/dGzghLRxcGqMTVUpzZRVbAtxA8Mx55ETKIy
3rnF+gC8il4Ah1EAz+FT0NuvDW1s5sX1N/47ywUM0DqiGPxuAUiOVuyfyWQSfLrP
nIimPd2Y0lXiHo3Lxxa0/4+1u1ve2SlpvmczIiDoNGkA1wBuUjryozhvNthFNdre
r9AYMfl/229TNDm6/33K4SH5ZIO/uGaSB+ElqskD6fR4zp38LxQ0IB9aApp1coEI
o9xdIVCZR92bwob74qk5XJOp+d0jixLEAZHtyLuNUKrGwvd09Lsb2iwDpAie7ThC
taskz/QIhsQK9JtbAybfykPai+7KrmcQS83vBP+xxVxbjtiJDxL6SX0vxhPJ5kl3
eIP+9UsbVxgxmy41Dpck59MZmKtgsvD9y3uorGk34VsomIuxc2NzkTBors/0HoZo
/hlPwwWORchzX9sh82SyTaJtADdNWdq1f6OTpUgogjdLZ0+wPuaFDu0hI40NjcWU
qogw1e/k2dBslJpHYK21oL4k4kpXnSzo5FkskmQVOtgHgHo30BCOViNO0N8DXWSU
lVdPOW0Q0uWzNhrYbfscK2lUQsNJ/4xw6iGSO9kUjx/JlVo9Z1PNpVuLyoV/fqMO
LblYf3eDuNxMzNCJf2HWAYfJ1gjvtq4ojwvXYhn0oPJeFPKCyBGEBazSh9OQRqEy
VniGdziKpaePhjTK3pkTGUC+Zaq0hOd5Koapcb1Tl/k2nkBkAZ9+A8EDfaDZi8LY
by1uefd4tCwyTmJdO0GraY3Mg3gNKLK8Lzgesr7JfC0eaioMFZlMAjAj0jaIP0JL
mn+U/DQXXRMBcGfC2XR+IvbsvgAJdr8BlQOOcnJQfwC2+2RoQk1vVPAZv3O+Jo4N
l8Ba6kiI5vXqEUdherpjzlcN7Y5mtluYP0eTCEjDvH383W5BCRZFUOwD9sD5iEtr
Y0GYr1VMXwXEG8wE7+QRrfIkvfaZSPcqbh8AF772tBlDGtdwoaxGjNTVwuJEDL84
x9TY5VBk3p2Bm/BHPi8mnx5GbBSSn5aM+52Qy2Z71VpvCFpwNp2GmIDfYDKnn1Sh
r4ncU61iiEAxg+ETJVYAEhiPlrPi9/KLMA4GcOvKl+n7tUOFDrVxQgjmzLBoIHd+
Sb2EWlCmW92BWgMkDOXKN3K3yO2m+fpU1Ody78xMjuKKA2QfF+N2Okp6c6ndjJFA
U1wn1HEOSUljeE3Vr/FKJLauM5t1PaTo5MvF7WTXByjoZUD3OA+pOGRK9S8LxTnu
/YrtwLPfpVnmIahW39Ep5ZW6hGRc6WRJTPADB2UN5JgPM165xHqsCg936MW/W+LS
Dk4bjnhim3A0Q8SelCjVK2bNXU3KZJ87+DgN5XoE+mv0pNboo/ojE7INoiLo/Mw3
mGuqHhZK4J9iu8qu+c+ZnfD1nbawZng8BSZZczrruWIx6MQ3idUtANyJRYwsKMGY
Nq9RbHseDjJyyAw8qWXrZk+9T9Z4iSzpmtkIdSYD4Wk2l7N1SX2dUhPs7Hlvbs56
X2kUh3l1WigCWOz/aHJ+p9Bsj3zepo8MT8kk4Wg0LJ40wHLUmPQbO72H/Uf2XLHK
dquGdVYo0mLgRyBO1NayEBYggI8OEQ5ZcngtS6+GqT71I5YTuRpWbaG9OfV9h6q4
mFRsA56tj67ZEEt2WhlDI5FfVsV3XX6LiMagqBUwm4MuH3c3FZ0TqaDF+0ngntgi
4t5gLDaSNg094UsTGsc+dpfC6+gQvh2j6Jcb48byVnAAiQNZIWpggCAiuWh9gkNd
5hVyXmNWKjWsns/XFDjtsOL4ixymTSiwIsnli9J/qlAMnpuSvkoo+2KhfUpBfXPM
kfuo+1nWfzkt4R/c1MyVpcR5CbsaP9wURR3u+L23m/roYQSOjzvhFMajmtiQX1Xm
NMNMI1dlLYbTHs3YK28XLqci6ftcw6+D/ggow95/ocZw94pOgG0jKzgilc7z6YDr
0/nG0U9Yf+Uu/x81eug+xBTKyfUtUre1ZiV+c/gtmYXjW3Cdb136kmAsYoef/4Yo
9cPp02KzRBf8sgCrhmIt8CRckuAjoWkq7n3R4z6DQ4kecmGCSRdc23RVpLsSN5uS
QrIrJrTIakedGmEudwl8spJj3v2GbfI6fh7guP0Xc1El3lONQLIZIWYd+sAw9nLE
zIJSMTRPFCRtC0e2BJcvgZnc7//V3Ji24nXwmR7ZMDwzNSzoPC75VbOe/bD6q0zg
TscT1xc4fBciEC2ddu5WRnStb94Zv1gERr8Q9einAl81CeHA0w+kTp9hZlTfedDT
PviD4pQBJ8MBOBMRWLGvsGNRS5tquQUFZTmx5fGrAyerzvIiUmzt55i0jtfe+ZgX
9kgm32tz8PbsWhenDd0dQS3JNuJKTIdB/qNSArV6/QekWL6R5NOuuIGlb/1b6Q4w
4+5j6urnOHJBlDoHtcTmW8rGtH0Lv8dkP6IeUhbmGtTLiCbO8i2epMQBgGgWMMXT
+dsJqVUPPTk6JrQC72F8f7FnQnS1V6YPNRtTM0fktQyXSFw0AZzDfkrGsk7U2UPd
wSv4mRlT615ebrE9SAO/dZaa6TMUNAUNAlC6h5dSaolzzRUG6gaQZEvj+BQa7S9m
mOWAuSRkrOlq2e5g16OeoqN2ITdvhTtXZAmQ6r+l9xsSEgjZa+ER87AL3jkyEg//
Tv8vRc5mBKBB3PhGWzikhN+rEnyZIa15GZS+LH9fCBWZPsyzOq/YdPl6t34eK4s5
bnR1XGCOwoZP98wfXgOjD2ono9UiKi19e1q7fHRBY4SqxhZzx0ZOix9QU5oCk+oi
WoabhjEXaiZyufhmqgf469De6zIiilr55ZCA93OdNLUNCvQLkCjyWj1cIEildI+j
c17LhHhg5B5gfT6eafmFhAqH3VOF1sXOZGVkrm+bJMmTaEs7TCMp40hiBfeWbAKu
Dccyg0rFiLs1yHIa01BGZ7PooG/80hFr7fFbA4ptDezOsCMoVBYz8ukpWJtnHOll
OFOeWQvaI2zfR0bByIJjQDS1Q/DvYPs9ANevx2AZLujDYvIIUpOPjghUOhkH9ITF
F4irEvpE3M3GdzymCZk1b2A1jjrv/Wv+kLIQrEqaztJQlAtaw1UWpTMi6kPQmjdl
PLexPX05S7Dm80vh1veQmgE0bOCEhj9OqGWDjHGc+h46Aj5AL4ZfRK9+kQoXMvC7
s0wC8BU5mif9fLQCc7yslPtJXuALE4tU8oHZFO6jaDKxvFqp4EzrvdUXZS6KVtjB
Um2i6S8fpTtP/VOqyyCc3UYdFKkK9aREGA7iVs8JQvlmzGqPHe5G0hcLNS1HgLRs
I+w7fCNt6QCaZ2I0bFot5CHxe4I43J5+7ipOs9bSN2d1+LuMGyHDRVsua/Cj5xpI
s1KBcZ3wkXtv1MFNhNRAG3hRSzghqOFo9dg681Dd0e45LbuZ6EzAy+Z5GHPZXIxS
twTr796ZGWvAS3FpmwTGglMuRotmBow+xeTJPHwtbs4JSZjG/IpqX5rZT8oitOsl
/GZKT4Jf7/mzmwMnaRtkq+1Gven0YXmYTmLj2hr+Kr46qUFp24bXgE3ir0/1FK7W
Wj/ywlLlRFJdRjkjLHfc61GHE2tN/AMhu8kYBIW9AiYxPbrK81E6iHJG0LSDlZNj
F1pT16f0DeDhenA9IL4A0cV9xcNSKOR7FXx6TnmAo4TkPmvVTZDPvUClpIZCiENX
8h3ZL68n1BpibNaXGyzUTVQloBscMu96OxWdFrlui4HBLdVr17kSydrp8df7fWqV
Sx/5kA5j4AyFN6LvC07y/Y5PiP0fOF+6dwkmEEPGDL0+I2ZwOGhsJC32bYv7LLES
IpQSKExapCvIb0P54bVF5KVwKP3kusbpnnJOEppSn4PTLdNh0iYJAvN1CE0zHkSR
haTw4j1VYA6p2ZSu5q/u9Ek1u1W1aKR37szZsnVQ/92rC9rp4RZ1cActVn9uZVVE
l1ty0xU0Re43C7gOmrwiejbr3ntCrz8JVdkz+L9PC95vHT/w5Acdw6QZqwHjJqUa
v4zO+IAXUYi5aXoLI/AwCEVFLnJjsf5TGxIYdPGmJlVWLsG4mziFznoFqmkhn0/8
Efcchsn2r09YXvjiQWI8GvghMnMLZufLJiG+ySJyKtoP2DRdVq60QfYtwxcFh60G
iNSYIPgeuGMnDZCIgmJFt9k2CauTrSXoxAILBUzZHyzMUhqwM1zpBWc+guaROUEu
cPpRuxSqfmaie1MXyC2gEVEpfs/6rc+3h0bwTKOzj1QWNS29Fb3OkcBuJfBIQKNq
KhuycSR7b4dHx910r2nmIT9M6K/gia76gFeyoNGO9ZUqKi2usoSFFPW4KcWW/9M7
5YsVxJZ1x0OiZ//W6tjBVFZ0IiyWp9lyGvmsnWvfY0PlvrdOhJ1LPPYhTIKe6Xch
vNRtI0osIqDummLhEumHajvaGK2cAIWrXq0HeR+05nulNytI9YoSPp4pubXNuUeF
VKX0MmCNS4G49epsOzxeBZ+g9h3Wg7KM3HmrLgssVnqA5l8+cgIiJlWMuFcqw/fr
lYxCsFz5mK+BaGLb5Z+573j0Nr+1Z6YEqmKUcfVEjkBUf7H3XSYhfdYAyVvtETsU
JGrvWe9GInag1JU2/epCQhEXzjipUWOJSHgZc12VknogUPbv9QsGrup8V8RI+cRa
Ku3euVWPnc1FGRpci4czWeyXjtoccp8oEeTe6pKeG38PdPv5DfAyYZAz2LQnRZ8r
VzpvSFW2KQ1Z356Eg16hlrSL+FG9AOC15FaUqq/hv5RdUxFxpYswE5O9Tat5dWjS
13pO4nbA3qy2gvsJuAOll9ZYExCWIXGlj7sR2ZRgFlGURXya4sfQcra7R1pUMirK
LSO+dSkjlObkt65hPyEtJLcxG659Oqo9I2DY2QUT3fVlgNxv7nmaTJULUq8FGonQ
U5g3SMvk7NG9fx/wf+xgK2wHtagtE/8kdwh73URvj1BGpQpCj7mUm/CYP0dBij+t
O+JBfMxpH7IHNUocYhAe08SkNBM4uSjWyDKNHkPwZRR5jt24X/rSl7iftq1JwgsF
fKph08ybMBA1kFlnTdlrw7I/CHgvydZpcxgaJCjkigXpw5g7z+3rhGtahf+zNmF7
vPVob2bKtwwc2HN50duaVCjVslmSkhsiEF7OX0xpC4ZRObRVEAogPajWuhY3lzna
IDZIyG0NlpGAQ1ApUf+UqzYY1vTxDjg9ULUZ6udFDbr0gv6yZmbmoLB9nVuFu4PV
TSgHnuyZY0qx6uTjAcY6mgrTKzgtV/iaZVcMtQ8HOx38sTs6pMUidLCpvosQ6mK/
uncmaKAPTdeFju2BrnlYm4GzquQ56NkdgtHaHJ5+IrNgI3fFQaWhd0IXKR05UAk1
c9BH8ARwkHAfJhhfjyHQ1P4ZpEOQdhQV6O9WwMb5cF/aA3Qdyo7/z482N0hObEOX
fIl0MTXrR2D9F5/syLGSrWxpfJ6Wk/rWanEBfd6Hg7q0u3BXf6kC0lbtrIaGbWj1
ub3Z3Tj+m4dDYipqw9mWlFeL1g3tyesUxXEx7zeVLOfrdOnMiQshhKFFq7guIOeJ
gJpenpuy6JcxwYO9zTubqGaPCbOshYvQvjshdzmqu/NXaEuWbZOGwvdemS1kVpfe
ybS6RewQO/s1XBSUIsxxf6285eg6TmHp8JlkB5ToL3UB/xW9mwpXJPQMeaDMRspr
uAFCBGLUEKl59/EFQOulktAW1fYdeWEJOl1BiF+XYjzU9Pg2U/1LqA5aFWQQ6cbO
Wxsi8+o8+x9FmZY7wLxteDNgnMYliKduglAbQj/Kz8gcbKz9QM87OWJDspYYfhge
3HRuJgwzfFez/h6bg17G4cgIEn+IDMY1NTZjrCsqOir9k/Jc+Vyry0bGkb0WfMFs
qJrEwhNKYc0DE2+NVSePCF2IW6nfn1dOJLxgqRNVByziqUf5IdXtg236bsiXUSyn
59WgW//xZKkzpS9BRrAykIvQxwBg2Je3RSwiWXZwQnTXDKkREZxDYvHtYiYId40j
19X3A1X642/JwnYcutorK37KvdUghpY0XQwsLxhrq91BJ3+CyVS2lKojrc0enGXb
fVvWw5Pwzx3NZROlNcTP30/ANZBd9ho7Yy3L8uSgGLwYhbgYQCs0qjPkwveuSIiM
lRZ2aGH/EIJBRSb7lLBeAomCNsNCDp3aW/3oQkY+LOUVb2j+584HxyHC3vGDzvSp
PkooTJIgawqKv39nZkn0mgoLKjOGVtLsQy1Hj/SXJHB1ev/kABVh1AjdK+1VG9Iu
LefVLDD5CtB0l88ujwE3u28blCumNJAreD1p8prK3Es=
`protect END_PROTECTED
