`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17d/I6zebFMszHp1dB60LrjbbyuvBn3aYdzSVhruQ23n2t/QBccVMnlj6EdxJ1Y/
Z92nmQI3ZDIIjPCokZYN+wufyWX/41WAb671ImZtK2KUgSI1MZog7f5kTpzSHncu
QqS8FyVDJlWYM2UbZdoMctJ/JZrsRnIbcc6EgGGx9lXQgBgJ29mHXXPNrL+xNc+G
MTdQGjF3eQE2lnmPMrs0P5TSmjdiZXvGwR0CwKSaeI61BKVpwzVvlui/vDS4Z/u0
87aTfkYBpyXB1qv4OhhV519uX3V97rr1yt51licCDpwHwRVDXZNstgpzrW0LuyBd
NaGfOjxgGC7f8HDf353Brp9KfBSJ8jW0H/QT7Xf8vF2AqW+RY5VyUrHO7+plhRsL
0E+ZajnNf7W6F1YNkfwjDfmfE3eU+73CAT69n/GhVBHEnYSICDpnRARtgWDNqEhO
mwaeZA78UlGa3fo7aEji36yIAqcuP9f1Cswen/U+Le/iWS8g8aUYlCGGL93B9yZ1
v7js6tbdAX6jjlO/gTgMNlLf7pqQiW4vPjTrKi2D3ql7azt2Opq6pFg4QRkNnNai
SGpzwhb5Ab6HWVrFsCJ/1EH3W4N3qouD8RiAHSY8qneXoqdmjzzIPKc0Ctmy9/e9
b3EStc6ikIt3xWHvAVY4TE19dskoU2k64VL3NOlPsoIzPlm4eLf/QU6gU/WYAaPz
oGJ3UreRqtEhkNdqGkQzGlsUDX2pGtOqXSqi9Zxqdd91GFyeqX/LekkA7OrS6vL+
DNwvrbEXTaU31TAhx+t7znzu2sQNMF37EQVOgopawmKoPpIoJcmXc2QhovBR8EuY
3OWUNB2X7yfDrdtTfVEqvrkCFUZ42uCLNtZr9LLwnZo9xCNq2AnrY2p1ehWVqC25
S4DtzBRibkOfTXyfJxkAXCg6VdC4/+1Hz9Af/Eb7sIwygiNC76wrVPySj4egTZ8A
L/xT6ingskbNo1nDeOXL2CDDmiZEPKHxwINNL55nfuNB/1vJ2kgAPwd7PeW0cs7L
+pClDvvPt/vQq4lMxgcjQTgKrLAz/bS+rsZQtRVnp1VhVPRVQedWKVbMjOmLT3vj
oGiHTi0J1s7DMWn8sCh69PYdkh5fT0EJqIrdC3ku/8K3jLpt0S5+o1fRkmx5NRzN
/qzqhC5dl1xL+ZB/FZvJ8fUCg/GUM5Ne7f3xa5q//hRGs4D40zqQ++Rt7oF1rybD
OWdrVNsn/dn/HKVQ2IQo5gddQHyMZWtDfyg6wneXoqCO7tKLHOFowOZSzZGkTiiC
BCJH1fQfA1fOLqXku812LGaKUPXe8Ash6Ruj/dlOnGvkL4oR06P/RtS0gke7fbvk
EFZNt4oCT6evADzbTs1DQw==
`protect END_PROTECTED
