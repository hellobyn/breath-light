`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkLmORa6xluXFUqbgXqJadJFDmiXj1Y1d8vpY0JYNoTMoheZoNmXQq3fa+qtOt23
LIuvaJxWXP4EbtqF273LqpH+fEjQz0yItnckmNdU3/JrvsB7C9zrTztsCpHldHz3
DZwZO0kcyaBhRi9KSZLPr6hgd53TqlQSM5ppIIfv614I5gM24drfdawBnwrlVIYK
l0f/WFcdTyYD9OrX3X0OjKm0BxwuaTIoFH8lewzSC2r/1AEmnXlivaf32MHMMfVm
WOSLLuGOpcpHq83rDUpZSCtcQQCorqRt+7a3hRmkNI+7w+MPbJ76E1Zs5kvsE5vk
3BwqeYqTKNEDqEGt/nr8J9ZBbsnZBk06VVFcrUbd0RSg9zV6+13YIFKzb6y2CXLP
9RCG7NG5oHZHjSxicyH+iSezaGsOnuSA+FVPoEkr9aycQ/SGRssTkTCXSRhyi+Dd
uCNfLi3RdLuKtUqDQ8Gzag==
`protect END_PROTECTED
