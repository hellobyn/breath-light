`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbyMss2V8OsLW0KVAzLQK4Z/XtA4rMOfMFJKvF4tIun0FCX4ZiqcUqaDFjKtj0+f
5H++IcbthC1vTwbMMCPyAVD44tdNHU8yzO+4RVQV+PmN+MaMugubzPViTlngIi2/
AXVrqL4WSPWYvDCLtC+SSNNtdpnSek8E8Chmj/aurQMF4YClfidGD37xe1ZxQc/D
bdIkfYCN2VDe4fXHmCiAcpnByIFOJDxiceAzmutpNydba0zeGr3gYxtOd07kvd88
OqQiMHiHz5aCI5LdvNSuiUv1BLu/eNlwnHdMFwRICIpoUM6cQYuldT62kbBiwsYi
Zmz+j0LRUjeCBqO8TenAa0U8/aslk+aMo4EUeY8Oe7NsQxwirwgSA0rgN91vLM7m
w6sibn5dlaJlDctdKv1dXR9xqnpjMBDXLFCv5A8gZE+fKg+cpTbguFoHj/5eBh1k
jNM9pPQNuLOcork3oa5k/VlltY0V8AHi9nyd0S3yqHRhOuACM+GzNsaBYE48Czut
52RUGVdE4GHgkQdXlm7UgDIMlNxYsluqKBOQe7Cn6owKQvAYgJNbjKWdXKASTk6j
039XIe7FxFYGMaCHsAuVEU3gZ9DRNjZbqWFVQSpBV9oYaOxTHRYI1F+9abOKrjO3
f+ExMdym/SZ9v9YFnUximOzaCx6r1ZhP6hKklthjAAtmdTIBsSltOqdE5PWZlieB
JNBobZRq6HrZKmEXD+wT5WRFNEHNxnLEWgrN7f0pYQxkaa718SIfLA2jvWzmz/i8
IuXIefp0ddOeyPH+0chyjvSPfucGzLLD/npRnFDmlsraW8Y/ZDDIYWp66DXsnGgx
kReoPb2emiuY1uNgaXLfLsOpP3UtaClxhBSo4Hz0C3lQEHGJiBfQmjGaigiEyeob
D0FaPssgrJeHogi4Qc7z2LaZsc+jqyF93W+LrKEu/oy1Vm5zlFf+wUIdx0ak3slB
PQjlVeTPEzWtQGT8MQdg5Xd5S6ljlLtlmktDHlTmmE6gjn8JQ/aF5oXXSfjp7fnm
7mfYka6qb0Pgh+7vpORZn7E+MHZjHMR1VyKUdPRV1JRP8ArPeOB3BcP2g1hTwAKb
Xd0IS+nlJdFvuGrbZ/r7nDAkSNtAbtFN8Y82We0ft9rZsH2ryEsqPexM2m3MGxKR
HrN/QvMIWJT4aLqcBAPtMAU4UMvsE39JxiC3dur/3Mj0aJC5FDFvLsbjgn89vnNV
0mrS99PSKh08uXqKFYFzXVhqu9S5wMAi7xtjouOon1I4tkyAQdrPBSzwSEe4/22a
1Un9bAVntUw1ztt4oU9CtGJaSk3c4oLcJxDVnc7inCLITHYzcvDe+4RZPh6+jC4j
4OsgtKrlXYmSrwFjYHFDSOVfPaWKuvNsCYIzeBlhZWaXvKoJ0j1vu2RC9RuUqz8y
5uJ7N7AVMd1hUr6v0tJhE9+T9goOyUspt1peTWTpinaSVZ1jgIK03bSInqlHLF90
sYgHuKVQYJrdHqGJY5HfqG5kDe92RMW29J9HUz0r1GvpUcSbyDO7LFpSxY1zK8x5
32+kTXffkrOWf0EQGot40pTByWCacTPdf2zEqMhX7a9j5xpuLZwvRNQkVWe5V1jn
H0Qna9hqrGQpIDRXGbeJ/ZBK09sbkupkqS+RPj4D9pRPSR7VAfZ7Qxj7JY0e7rG/
F/9bqgwpX7EwHLEyVZAHkHrsBlsjU8QlT0bZm+D0F92RNLewDJl/EhC3yKPTEUKl
3zgYcmvqf+HhtjQevzW+RA06tT/iauilRH6SpiJKODcV07XsHWEJA3lhvkNDO7XR
kmdbTf9gSna7si5g3ZJ8BdHkqWQ8S8rswqIfoBwZWxGCnRd18oJCcn67lLk0ctWw
08iFuT4slYu1EzkLweO3W/1wzqiNw5afRBpU537ALgRaC8twKeZaSwxj0zsdRD7T
pBVZLMd8ne42IjxaQQrXyTvq8wrIKZXL7upWQeCv2ot6pOHE+TdlY3gSnlAawqMx
kd1SDiUrbD4Qiv2ieFlgnkXu4I7edG2HNio2VVjSmjHF6thqvgrBLohz5gdX3gX8
4+tjBxR5oOhVTqWhq1YfDAlpGSt58qobUujQ5MSkRiP1tpCy+PzUolm5aIPzg5ew
vHsB7+LpCN0BFJSrL6J3Ezp/lm/+QA70zd7nrnpfYb+nYYDLnpfjZy8ryOWHnYLK
KB1v5flDknXFd2RzV/oyeyZBQY+pWpYAo53UhrEcY3QueBjys5vBnRqhOpkYBuky
69yzutBHwjyBeUwuAcKtckRxPqj487at5GajqoKwKM0O9lsjW0+EYht6Q4TYNcis
X5tALo2SJRG8LaNskV9+k8sZBsf0hSn9GEyJEMAUpxknCtuysK2qxaPWDbdkI6Ne
QMYBSWRFfGnR8YnDr1yibXZ4IIQUOhefJ13IgflPJCF77YxlyjQinIgwR9AUAMBX
nmz+df0MPGQ8gZPsWd8jnWOPCjBRI+Cp8umBgGGpYYOYv3oxtFbeZIJK2QCJoFTN
X1dyYY0W+yOhFotTGa9zJHGUlDJJhsFVudk35nvZTMVoOurhi+ozq2XBqLCmUDRT
OpXu15Zcr+FP/ILCMHyWSpo7LgEpiMsXkFIGLcUPT4U90diSxgF0CpQ+0OjYocJ4
O0u/p03C6rqHpcKpy+HD0ifoDCbntmZnLrMOtHibI4icKGRFmZYrMhOq2wBcy1uL
ZtYZ5WAiMC5zftA7jfvZxGP6AL9+EXCPpwh8gkAftuJ/HnI9QuwXXxLNGavq+2XN
SiV0N7kedYke5Ww002k1kDmk8nSoc5nj7jyaGeAGIb6lwEulaHYoVNu2AFu2pwRv
iZwqAE2Pcmj3Kgvp2GdTbyM1ywr6vBnLvzniKfZKaXAB/NyRQMJSCasMKJXne68F
jWWwB7NuQ6npchz0qZeTC8kCntUlpKnVevEB1lph3UfFibvgWU21hcAgBLEocmrP
ZyAC58boL6vDGz4RzbBQAMInV3PYuQdSX0w5QlY1PaAggwwr499ao0MG40rFVge3
DXCMeFxyo2X5UcoD9ymNG2rlnS+t9srwaBg38os6LltJMZ1DiV43fW/0SuCHNzkM
qtCUypHoc2N8n6Y9sbpwGz+08Rl5qZbUcVGO8LfaWRuibjy6YJv8m1os6R/EJLdE
HNQSkcwFxtdnIW4hs8QXA6hzLDLHoMF0ydzXYQlGdM6b7AbRGmcKacu6uNB6YbcM
XGaiLgVMZlfaraY66nPWTpBf/fRaSeM92FuHE0xVSromeouHBqY3lhUbz4hV8aLV
d/iem8pA9jly9SVIPy8bI2ori3c2zO7beH/7KWoJ6REXOndsQNd+KCfEBuMMVoN+
BMXJPGZ3WvBXRWUkXLIKysqY2rrysUzMVhYrwkxZhNeQuO6/LZ3C0vydTT/701mW
dQfRcnfCpdupRXQS9SrhGtBR5Ia419boQUNxPBJV2kK7pP9YoySgP5sZl3wFaKL6
EDTLIfg7Jn29iDifRkD7ScHQUqhhzSfbywd81m9399Hwzm+DQdXbWg1Xcdrxtecq
Qiej4aTtZz/epfUvv+qaB6HK0/B0SqBof0aDd8z8Vbu3RCVgv+EtEXiT+9Oc54KT
yhnAB/Ysyz5D7+xMxAUGCdp+sx6Jotz0KkIYHFS4XKt3gdcTdw+Mms3YImd2sQ9K
0OaQyT9z9OL/CCPJS1R0SWWnAm3D3x10OcMk6xYn9hlfP7jrEcgi7T7ngrPtBojP
sAz8ttbABSYAMUI+jt3EDNqXbwp9gTwVkM8GN4Zmeiq/2TEk8+mr/1wIbq36AVDd
lLKwnmk4kUlsnNPxJ0B4EUs+ORdaBfUDKKtDHq3xUerKJfW4ZFN0mdM6xmzFmls3
QoR3z9T/HX1mcaH8KDY6h+QBp9LXQH7xgHsgGCHATKpa3HuaoLDTOYWeB/Q9pUN5
bRYfZgIhtCNdBt5WUyTZ0BiF9OWWafjZekpiI0eWp0Lhw/D37T8OsO5swX7klFJV
ToKKTIWukmp+g8lQo74FcHePk+GmSwyRrQ4Jjx0OaWw5CBseacM+10iH3RbFIPW/
cMP2ADQOh4dmn1RJs+d2pqsRC4cL6B9W0AJoAjwRvCRbeIAbCaHJUXOg8Sd0ekW8
o7QZmYYc9hw+d42bm81Ub6Haj+imTqK/ZoRRvSgmsdip64twZR7FynQeEYk15NGZ
PVtw7f/bwNNMbWlqGAaRYrLj0wVqaSG3EsBShrSrUAqHiUOqP/XcWfTW8rczeQt1
gq93m0/1Ynp8YRSWtcBR5IgJ79mKMbbzVgeCFLHmyJHWI4EZvSFQyLO3ETxzDdr9
w84H/Lv+5EyUj1A4I+TD+fpiHRY6GiNvlTVYiKY5jM085qD2FQ8c57Chg5sh1698
MMzgEnAKAOEwj16F4CdGj1umUlpd5srGHak9e+Wjr2HtYYNuOd8TRW2uHxtAZiQP
Vt7Tdr8br8LE2m7gNzWV8g0QgFsDqjvQ7vtlUjBrU5Vhi51f0AXPUHpKgJoYgIJv
aYTceu6PndeyQ0aAc7bdalBRYbNqL1eVTo7O5dJgd8mtJKArReVJmfuV969CCxeA
NFFeNWrP8WerbdoyZGl5LeDEFpSgKs5Z7QLGRFDrGyEw+B83r3Lw+iSNWxrZxhsM
/Zpcekw1oXgBhIbokhUUBu4XQVUqRh2YID2Mq/k/knIYlyVE5oJkKTpOSbUh9HSb
jSPbnVZgBBRbda+QSB+XLg/7GO7jehDdHBsSOidrV6ZI35KCniaW3gys6ph1nGoU
UHZ8kApdoxzaPasXybhbQ5iGEpSiW58PXHmSpSV3CEfN4Qs2TaHDYglqx5PSAfMw
2esZlDc+N15KM4LCZQ0GS62qy7S7Zvtj6YxqXlDd98y4MM5FtSAqfcefB/mP2vHY
J9d4f1KEQ+Q2T+dq5nOwBtRVEu57hyKmj41PP0HEfNpU+4NU66OL/aB3AmkgefI5
zkIrmDWS1UYXPhW7QZjwx6ZFhg2MTnQ1sMfK1JwRa1g5gZjzd1zwW7Rugb4+/vUD
VwyTye2YEjZVg5KGhP6qLTCLEen56ZWNVKTrk2VckwU/+sGZX0hDEd+NPVW8+Kws
6exqELks0lZ0K5sl9dOfexyveRKfA2EsIRcOoVjzWOhpJQ+hr6AbmQOWEoh4rhDI
viA9sTMniSxBJI6H/2axrpmLe5OFzFQiZ+VWCBfs294TRwzJUIFkmSUeAXQIfQcD
j5qfSK/BbHv82Z6pPr7PmDIs/effaSO4x3/mDFotRRroNa+rO6J5HC+IGEgfb67l
jSOfmCB1eG69CIty6Dr0FaLFvv03lY84kEHYIoFMBk2lPQ4DGPPvuyZBMLdWJ6iJ
/QL2CBGbAmOWScLnmqP8gNrwA1phYSTEc8O/dtGiETPDUjMt0hzUIytp7slKCkF/
+pw1l1gncZnmYvBXWEAYUKttXP+Rje4PEVatuy4lEw1+XweIxBeRn0RdFgtxqH6y
qwkZQPRLG9oC7dWkEyl5PfLl7yRGQBX7kwRYBadsEGy/+v1UneYEaybsB1EF8y6P
iBwoC4GXFZiTLYbd5nSTYc7XwgOTafeV1htI9R99IXqqEPzz/jevY8SpmrgEACho
lM+opvGzEu/ToxCjOgleSMzsYc7TOf6NRM+f/+szMFKweXYeoh3UIhEPjG/GcWIj
f6sLacUR+lkN6L39MfTjgJRPAh6lQC1XgLCEYjVsw5E7Li47J8LDaHoa2ZnltAsy
hCVU9Z46h72xAcbSDcO+AbznG4qaj6NmMVqfvD3BAYah21sA5xA8oy1Ph1oJ4CEo
OPoSo8/K2PCtcKB9TSmFCfrTXxfy3Ndd3X1U29En/sFMgASZyUInxxP0095f5Wbo
XwUsMIPvtUf6ABsdMKPmSw7BJsFeGsQsSuXcfo3B4u2QSEdee0b+whNF/cG5IChf
npFWDwVe0ZIIGwIVHDVa33nFmhxCgLGMEN6z637bqJYiANdFqYa68HkLwGD3g3XS
jurImAOA3z+Hpx6+sEAy/7Y8IPrY6rlwxai3NGjrkLCw3tjRw+tae3UPbjJZRG+7
wlLlfbLmj1cNmRfADPkyU8MtQVoxK7Yt5vh8MAGIA/ra8Rfjc2S6t7hzvlq9rl0m
Mb64lsTyd5Lt+e+M+o3f1JtGIY0pH8TpjPF9zE24UH61is5sC69W5MauCpCo92Ph
A4faDZPRuMEvEqwKgYMhEaDLwP4sc+ndcoLHE2IxkbfYoutCjfqTOu3HgQDjoGVY
0FzGEpzS71TqSOSnchUNsyWUyz9hD/cCNAxjPi1osns4KkQ2f4ti9Vqhjg39K5mQ
PWaq+ep4FQU1Vl0pGp0qQ3hFeUKTJ0jIX/ye08NV7RiLx0vU35gq0JKf32DeOd9U
EO74QG1F5sV9wGFBJQBnW56IzPh6Oq6JQAFLabULkL1q9mzUTFAC1NRB8ewBknTu
5fG92dLuufp5uxgru/cw8T5Ui8YrLkiURHLaKUoRXi7GJhnqAHkVnQrlZFHZUVnT
pZWRdYR/T69lDaedl2mr/eBSs2NMhEm9XiBare3j6jro2dwagWHmbe2GMBMIU7LX
KZdRQwdjqgosjFw2dooNTFhabo8EvATtkDPWwCscBcY5EhGbRIvprTse3PgWn7mO
pEVWzJEoYnV7gQzOwEdadXRNd+Eoj/SSDI3FkWeCaxfJWOehmrefXr/1NqAKmC8U
GbT74WszbGro+c4Wpf9YcMy6Sd3wgol4qwS1+7ygI9QGS9a3c5EomN4KnEPQaQwV
OkE+bUDy6ft0S1KltS2b0KpxcGH34OBrvNcd1WlOxtFym6Go4ystiYK1HbQpSbxV
WUTSonF5yQMdBPSjBYYVrjXnOq2MCU645nnorSp3I3njtDgIu2DCutzbxWjKypss
ppLj5owJs6t5qD545u/oo+SVq/dsH1GQCh5GYkic6aqPJcmk4gezvJyLR1MUXLRN
eNPW48gdCYHWbqk3Os/MVmxAnB1B+KkKcBkEKF3p4CVNgdV1pegnB1RoEAh4SRKS
raE4Qo0wazHJPEZ4hIqKIPcb0Sp4z7y65eSbqfoGj9/YcKqENC5ORSFxiZWL+6px
ALVO+OELnQowG2s3MZkzYJO6i+tPKuia9o/JOLox9ISpclc/4Bs7NguOgOqeooAf
lcJ7GDCrvBjSnJ0+RQrIF1RqUalSsulVwWxTgRDKDtiNJhQsOXBJAVtQxm6BEd0T
6oUHenj/oh45SQLurcrlIMO/UrWX24B7EDKJ68ls276mWBrguabh5YgWIyvKiECd
ZyUl4BGNtmvgOFc09N6rukzVtKxnN40Nw0CdTCv7Puc9XMynvesPZh8rTWrgd1id
RtT2F+50zyzIr0RzvdjCOoF4QkGF9YpbgNkFCMURoKxXLviy8pbntZw7/usPsLZL
N8ycy/9Ur5rG+QnpRRhgjFPML/1PTdDUyj93/pMbKkJB7ujWxbtXgTVuQJ/AU7x4
YCcTWx/6o4QCaH71OXd/Fj6TDDS6nd0CCw0BYDr3hXTQRuWoxAm79kLC6zuiC5ii
vGhZpNIpmARe785R/bM/W4CeXgqnkpOrapwj3Oj1yf6wGVM38yO9Zska+ZTG5PPf
wvm/i+cOqoL81RRoYe2mAf7WtcfhqsZs0VXPZ/n1jRTxT0kwlvPNARlQmRQ3Ll2K
fsL9qsMiiZhIdvM8pNrJ86Adxfdds4Sh9Up9Ot6ntgTg+VXJwPUjDGioZHumUubc
VIURZNu429+jXgWw1P5gvPcBNpIUNCm0TOnwSWCS6CypUixr4gU0kgpPD+Bba5xr
ffkmG3/yxZWgYJvGQTEeIFwqgAXKgdwPzPDcpAUB9UJaflsCrnbx4Cc2fXr3Cry1
dE+uXkHhrmXyXbmz4ICD3fuvpyZ+B3oGoJLSYzUVN+txnYM4PBojezzlG283k2xj
XwM47JiDYO30GJKn7jCkOQxJZCohex8AYvuHMLBZs/5LO057/PB4TvQX9UAunqBE
ayIZj8ACwsbPzLYA6Rm3r4PFasvjMiBzzzIpO6skCu77bmj7LlvV/AfTctSrOg69
aCHbeYnl7ipc1bQu8Z8rN8U2rDg7nnwi726aD5lmlce00k3DXIvOvf6PsDaxUgAa
u+/GW1c8riKXPVFvH8F7lUK4ljkTmr1mWY8uX/U3PN4JrCE1LyGeyoi5VxDu6qOe
iKMQ653T9V6i+fSbGSb+RMHVXeDTLsXhp5L3PuPH5ssczZwPGUiSAp0+ciT6bzzb
eCeQNYH5/g7rpZw8TlAKyHQrnDcd31uMzEt7T9sFrPapIbGRN9R1DSl60tWbeGQb
gtCpFN/WRosSnikZmCfLhc2Th5kURm+KARzNl0limb89SCs/9YlKCdlbRgxkOdwR
d/A4+4eTYEjChogrGf8GtYajVzrzoIgT8Rc00VhzKvGjxpGC/Ujqq/baDtwdX3Mw
3JZ/koSwOAZPwoGicGXwyS2gvdd4NZigMA5iUzNqJDrbPHn0rO6IXGImEWbQvspO
EhKce2qa6eWTmawMoItVi0gmYvY1bSNQ5OnF2GXWpDjGvxGe22FB3xYtmpHfFqRv
aVQ5NuJxQkO5Vc9WfOacueYSS9VMZJ5Sipc0zI6BkLAIvb9kiN/kQ9Vq9qmgTjDh
n5ZEjcZIAi7GZAbjbKVg6w==
`protect END_PROTECTED
