`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nDNPCpA74BcXdYJciTKO0tl8whDXBZolTNBGnN56b1hBPt196nwFLVX2CR0R2RsS
pVZv1Uvf2MUSN1MyqVZe13CAVg4KQNNb4ktzdFXrs4YxkZ406BE2nByLTzNIRquh
O7ypt5jRmP0rXBr3gTYFABKAjczUXt+ehvjD1Hck6e092L26axalXyjTBRIN7jf9
3YrOrYBpbyghKxQWyjNSLn5kJ33HDO8cwR7YdWw94Jy4GsEUmxqaHY8Tj2l3OTJb
luAb85T+6iMOCtlkvTmrlg6vtAz62f+gka1+8Wb902UuxTyf9Ko7IpSZKvJdP07p
jMcHQ5GyVqWtL5xDiEcDdHIUSly/5ZbJryxxzoV4FZofQn8InBykfuslf7ctAsOS
uGs5OO6MNMmAlcGmVZXUQA==
`protect END_PROTECTED
