`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7awlwqOJIeIPWBij0JXqn/68Yj2yk2nMOpKixuaAVrYhW5NK5rQM9d2GPudSpCUd
Ba72Uzqewm0m95MwabWOsPtnLIBJAc/aMDMQOWsY+cD72UYzxN/45bzUm9WqyM7W
uvELVah3CJBxlydVi9pPnH0k3YNmNUdUigtwBKbYYVKDA/6gG2ju5ABlbILKpHKG
D7oz/0+fQQy1N+dmjYnImpuedDr7RnAU89ttInVTen8tVXFruskNseNfLvQwkE8H
bhBPCTYfDm1jCAxNMh5+Mk6g9aKbXiIHqWDLbZFai1n/f7k4xEk5jLrpZJgV6hM5
H+oShTjskH/jteLhOE8zEQZQs5vdQC7woxxLHmcmURW53iLa+Hrm+0fpr4yJginB
RsZXWomiTQxO1pups64lu0jbzwxNX7fVrkz/AA9+FDf/IyUoqiXRZb5EtN+glAVa
bkk4RdeBMGS+w1TCA2HAp4ehRrR5ML3tvtLQGLW+hj5RdrHYQmOslKbnkcdpVCeF
m3MHiNDn1rTK7lvdkGExH8WMsS7z+K3khsd80kJR1bRaNMTtPBlaDW7DPvFzMavl
IaZFaUxtVnHKK3lkSLO/inB1fQzp2S0k5/2VTaEXhDr1Pwtw1TolR9OCWXnk+ySt
tSzAmSPDEu4LkUTmQSlNf0enV3ZAPcSrEY/gFaDHNueTI7ZMsIT1vqjoUb6rFOMt
w9o5yM12xnspFOTuHp7RfyQxIgBqQwXF2RCJf1i8bSYwYljfTXyYbsRsigoO2kv4
/uOeQMlMZkZcoWwzsCdiCOXbxUB4bTtjCGjV/VXUz3+vQneb/D3zZy7XqjBgC3X3
XwsCYpOF1/tly1QaXEiUJVhMaIf8TPhPno+chpagM98hmNTx3pe+YuTEwaG+BP4/
NFamgsw8BraYI7n7yo+eAndSV4cw9K3fnEXKmV/CD5puTOfJHWOBfkZFc9xHvAQz
q3SotY+8fPENeip5Zpz23lliSt1eaK8BvVMbvDAcmebqE0nXrfEqXNwH++2DSC6y
vMz/VKqQQ+lrnkXRaHXZG/DhiJ33iBe3jFbrofA0q/fJ88zCJ3RhT6ARP1SJ97t4
jq5pD5ocecV++k5u7NjWBY5Ns+rccL8EzrDwy2+M/DTRpEtmH95Xsdofqlg/WTRn
/g+tL74yAsNt69O2fIDZxJdGYh8QCGmAAQzW4KiBEkixxOeErNK9GRY90svrssFS
l65N9/a+cLdIHlwgKfo6AvBNrNm/D2BpaGTqrHr64/NluwG6VQyPuDNoy1Z2RHyK
36A6yAT9ftGTysNuDfmfenFpIJtZ7Cld3N4DrTXJhARJvKy1S4Fb33YRhigSGbia
1eJC7/WcApbKxEEhtah4sedis8CFFJrZG6z+Fw8yEeoFZ4VlxtlXU+1FDO22Figp
GpMPBtkvO1fG/SNDqx1RZ9kd8HeAAqSzbSRRYG5bDE61YR0KJY2+xYDUnIIg3N0+
/CkztV8Q7Ah0tJZ09YS8wrN2QQcp2R6x3VCuEvVix7WK79jdGZwK/bbCf6pZBpWR
r1dFAeeZW3ZPYwat2aF3OuvvVKxV+keSAcZqIxcsWJmZWdbyHetfSnZrZlApqqYQ
jI2F0dwXEvN6I5/iTQXVJRQMvNEI+PO9ZqQBUDb3TzqDmxc9OzYFIeJoNQjTCSDG
`protect END_PROTECTED
