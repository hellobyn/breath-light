`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3iK6ZXGYZvjNqNgUMSdaHEr9jhaRu5np7I1Sy8wRu6VXvL8dlO0sjXu9TMd1vbn
ptQGYEFRJofUGD3+4FgUXmpoAOEqNuLcJeXZmr9YjDmlCTJ8OyaQ5uVLmYLRFmXv
6mg0O9xlJiEDvZPlrsNenbaG+3fEimEvFiTvOPxUiUWud1dqPBle+VlVj/IOxTWl
kmspcUaitTG2g8G/1zrDE5/5noBwgATR4xuGg6er7bWMSj6Rb7+fsAr0j6kJAP10
X15+Pb/iKQRN6JoRtIRFGt/MPu7eYX/ZkVFU512pV78GylbYbqNv9Kdba7lXBadl
bYG62p78+J0o8rIPUX2MweW6D2lS6ewL3xO33olWuM/+wUSpcXAbRo2rKwoU2lIo
UHMBdhj0uB7wWz+ruAU5I9sjJbH8LVi9NLA6zQTn5W8Dwnk1/aBqyCjk59fnMfga
7fLNi+uVhDWx4a6CtZPLCChUV7aFoN4nF+8/Mege0r+9c7L2cEsktpiYjNcg0yMG
4/uZhRAk85lDivC5hVexft/HQDTHYoDQ9Lpl/H5FFHQGiO0knxIlxaulLTJFO4BM
k6TTMPIvJVCm96GJrWxhtQv/hhBGWuaSvWlXAyZl1tc17czzYkdArUP0HUjSAhLh
FthTYyD5JMudAogxsBHnMvXDIKbYhOs/+zhqQtziPlb/Dvpz72qt9NmUCgDo1tjW
uqQKKkMrPoTPWEE3aRhosB6pUfAgsqGaGGPiqoCJL51tss3/1aURTnx1ehNibOxA
WKMTHKIwy5XiaNKg+IuvBpOGOeea7jPIIk7tcoVCOHIX5oUknM3kxmh6Yd9WDwKA
Gtc9OmaMlu+8n5AEYgZyUYVEIwlHRvm+osq2GvXtRXux4zjk3JHiQ3JhEtX5Vz3U
/UW05pCp2IuLntn6bxQ1GoKuY6f3OEDvSrAsvsH4lFN2uTRTWlY8sKphzy2+YUiE
O+uruLP/rkF3D3QsxN/DKZWT+2so8nx0A4bpkzWO76A4BzlAhoEQq3I8yc63c1YO
zuk0qcBeYdMTenJd+t3Ie+cDuaOZB9uJxu03cZxeLsjEzCyeADU7Kn1Sm0caahTJ
JkjAmnWgdMgwBDmJuAXal3pk+FBEuKwjLF7f6HdY48QDhcQixyykFznBQySJHbSp
uEpj41QIM3N2mODoVt9NW+pFb+rnPfJ5Q8FEJQZq+DC8dB91R7rV0TPqiWD9kP6y
4Ezycc1H7jaKyVKdQxCQE7iUvxQy9jhCnlb+X57BZDMNt2BjZbL93vkBwAcRriJA
FwF+Iy0auWwqem8TPuA5N7AlXzdelgHnQDw7DRudFeBj4AxjQqykismVLRVyR+js
Cr/qb2xpjHvnbd2lVv6iWxv/2K3qR+Ion6Vjv41kKYb6SXoUDcd//l9ApgyCWUkY
Y+Wodyc3vGZyTDelyfDCVYzdkdI6jLnPvNVh089hNxRt4NmXVh9N50hpg4nWdnC5
lK8aZRgJxGSh/ztOYags2ftuQOZBGCeB64spwHBha1/5nygQWhH//X4qa3xeaxI3
TsYw3HKHm03NUO+1p1gkS/f/XSlxIqUMQpq9gN4V3Dgsmeurm3vX7ja7vxopSq9G
D6XK5oFKlpYZ9S4SONGE+eKUwQgUtKZFaKQLZzOh5czfJ1Wf6v6Oh46AlRWtBKks
dm3iGgYYmGmmYZC5F54fooqfX95hfmzrWDq3N0DSS36R90BjS72VciV4DaD2Tc2Y
bEXldo7JCz/vS5RVK0vf8Gh+MZRNobTdlY5tmb0sxwJws0QPC9GF9p0iZKG4Uf8P
bmcGHPZtbcKkPAo+Fd0/D5Wx5HMa7rEN4PlcQb5WmiNzilC18k0HoDr5qzh7wr+s
MSf+j+f8RqApJkGI0n46Wpnc9U+6R7d8kp7W63v3YIOlOJUPLFDRtiLyjocFjhZS
Yewhr0FawJbsDib2orBcUx6I0Tz43F6mHHOQ3tIhVEmyX7T1K7cnK6k8IUU1D0Gw
gQIvSBU5Xn9zdCM4Bs+Mg80hHnevuGOVq6vpGC07ZmJA8W5EkUUmJYhdQXR7h3r3
tYn7UPmhuQ8IYKCVOFOaGULE/3CX8EXAoa3YSGb2/9mof6LkWjrexUB4EjnZ3Swn
kSqz11/Ul7h048r/6lTVTSGA+2hVrtwMws6ztzf9Drgxu3XGlL3hYodkJIfB2Ply
dziDK79YspEilxns9icRvBmk/2TGLuVdoH2JsWY4FSqunTVA9EEGmKg/PKUm3LTt
GIqSIrcwactQTvoOPYc9m1xNBPpQBsQ6AQfTuHIWqbcqQSDZZ+3XBAMX73eNp4B+
MWwvx42JiRzi/JLEjnfI0SqxJQwIliQZAXurw+f/4nc+/FnznhQMepYvb8aWq6wE
krDPTrV90kO/549GJPjtdJD0ktOMUNUE+W1TeHmSHYOb0REKlnrx/piN4sk1kH0P
5Wr5uK1DEOEyJdTLqvKlnA+73iTtj2G4tDgoOL+nbSu3ykZBdcFF+3SbZNuVhLsJ
cLkqRFE/jxhpGDsX7OFJ1u3QLSwtPYHlCHJ9bxnCJz2tYmmu3vfOrMVjfCkX0OxX
QjsAXwQggSPzvohD4SC1uziRG/li/8HWD5P63g6sDLxdkrNTegF+0R5TsRrqj/hq
aCMnjQTjHudpnoYsvSRJkpr5I9GsugscIrqNgonpCpV3G6gO8iAELlRRTxkiD2BH
cIyEX1948VANsA52oy9Z4YA3NVPTqIKl7HV+Q+BLF0d6WJzL0zCa6R6pG74XB4bi
MylYsq5rk3uvUtw/0isRoYFQ1fJl/l1CXEeKZ7WrjUQp46Kn2Gi58OxewsVIpFea
2hXdJpPeKHhcgBPmPlqA1D/8XeAQ2YSpspxOxjNa17YcSJjTRYOBIrJN2bpqdzUj
tA0lG6ziaPraQDvOP6b3PwDUD4tk+/XzGxomgp5Jv3ChZxyDISUTYPLROFm0ntcn
tCxJVzonqzsHZ+CtV2ZlCJFlxdEX2fDesTduFNysfsp333JUgU83Btg8Ls+1rQSs
400/Qnyz72AYg366u/d+68x4us7B6h0oJFTVS24dLyJRsu0JTl162mHAFqkas1pr
xyeAIuOL8oFGAaZhvvYDlSn2cGIZOPyvS3nn4xt9mJFMaP+wuQ3WMz6S+FN5mPBo
HjQDl8jkKYPN7VGQ+9+i4Iphp/mbpBVQl2f0K50vr15meeLjYq40eZ5t5H4i79S3
iNGkIMoj1EgmqNa2P/VUE81GFNgqJJnL7lwr6pZZZjAnHxGKFZ/uh9bCjIW+ZB6J
o7ZsY4naWiBW6o2XCvCpsT6ZiRUHwxTkpxSIedEmgAlmRylBTCJMV6lV17uiTOi2
tc5lUkMuj+Fef4FAI38e8GdxoMzkcmr6qVHmDXCOCTL+mzl7TdYOXemEqb4Y85T9
oDPYt8C6Dgj5gmAIoMZXDOOfVIK4zaSxqtoxIC4WCo4OCxJqKJSxjc4gqmSNjRpc
qHITTz8BpCo1n0MpSuiF0lQsgKfNJ483mgnYMzhSiCdu4Q78rG8X+SvMBUMNvs59
HN2vXP4lZyxplaicB8qmSA+vMzETdEXU1egUo7GJvMwbZ8AoRC3V3ebdIcj7RueO
Llw0Z1XD+RpjQRlkTfHaDXJsLbbOModC3t9ZbnvNFH7m3LmoJw4AN/cwDvUMHpm4
QfarHEr7P6M19XDg5GRydU2Z3ib6MUc2Wvta843tsrtP+b/fq2uCkhBDLIhc3dv/
VAXd4DvrSygIlCcR3MzDrXxo4ucA5A1wr4iM0XKQIj2yT1ZuHPzFZH4Kj2GI7DM8
cgH089i0/hdP60vqEqsIsulQ+B+O2L6a3wBRLlvrVcfPQoSEA0qeIL6KlqFGOSHy
xu7tbme0CrxwfOIdEH6WZxCJkOBHrU7PZhbeJA03aah14GsHoSF4FBQGlfb4IXAG
hZoMDmpR8dKhjvYRdAewaXMXtuGrsy/gQMdUub/7lg0eB0OYjblLiAC/yJSNNVR2
F2589OmXzU/X4F0K8HzA/YZb8ZkJ9a7HFrzc6uQwtogl9HjJuGUDvtRhmAFIqzbt
7SNILgF7F8OlfTomdjoZVzf6Cv/BJNrkfI1odORJ8XTyRAEHoMaeKBt3FBymnk9a
z5S0vsT1oczlI1oXSkZJLLJiSOXm61ds45EbR1lth6xryef1CO9LQKd/OvLR3ASU
L1sMyDeBZh0ec9muNSseIo7IzvDgozZaU4AoXOyN/8knipfg7Mrjbqt/lO4RL2jE
PIoSLi0XHc31s/z02C6hS1IZDVjP5z0cRAZYBG9iiQmBeqT/lI+MqdxyfbFSf4Os
chpdftM6eaIA0Pa93waFWmUzsByJtsF2aoxNaj5IJ8/6DcsvMyw6UOyHv54Dwsh8
5NaHO3EiB4s/AzshzkX+L9A6CD6D1i+xb6Zhjohr94MqlL7g4ToTJ/YTF/uFkHSe
X7AJjKc0od8UmuOIddRqoUadu59Q4RX9ng+IPuW2yfM0YF/GCwMgjBtoFws0faAL
jm2JsihCE7xIltXBvmiE+aoMeMn2JYMQ04hfUs/5MyLsFLpcw8EHF5jE0bwyeVm5
N6lx4HDygS63ICXV0a9ezZ6KdRUxzL7RnBNudMGYxWZMdbc1Z4ovprTftrroTYVB
PeahgLfznezDf864LRlv4A==
`protect END_PROTECTED
