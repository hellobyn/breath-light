`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edULAVCDn+wjMxRdpL1JjlXgzcAWRRl9jFPRSHmnEeu3+bp7MxsYQmaF/C6knN29
Emq4OYcR0VqzuslE8KwKy79GN6ZtIk+Rex9B2z22OXM6psb1EHjpxpG4fSPPJPsV
42g9tIP33nI4slSLIqUUne1u7MiQbJIyvUfap8AIlH+c3+MIeXlcJNb6Vj9zXuDr
QnzJdnAxq0u34F6XBRK+6nlDZGd9I+qg3tJguuw1iVcHmgjAah0FGA+LV2ukb6uS
UarQaiyoFQKNVSXpPc6ZpwjN0qGDMeWPbbrVGYhg2JD9QI7CbDBQabVNBvu9NP9/
4MszmCdbQIGMD4OYAr13yiBo+CZJ1xF52I0Z2hGHiHXDCm9pgnV9fdIV6+gg51UL
e9n/RTdd+RUP9Er08L9irDWmgnoKGjhL7YQPyTzGU23zpPE4NP8lGDzm08DO22ov
ykSOQA9N5lM0jHpajJqYeS+m/IaOVjUFWFlV74NaOm8rAX/mMm1QcNFl3HKWjqBz
gSsRDHqBon9pdxsejgmk3TnaOcsO51PLYXPRBEK6coRk8JhsvwAbUGqf5Npnw6Ml
W02xgta6OaYBS41GsnuTL9S2lb4KMoFhZaXwdvypOKvNhWNRUELojDc7DdgWTrL5
jTUcHwF1lhdDUtCO66BtxXHLT6AlvovZCXPrxp6UtAv4uKJ5I8NR3qALzjiTIT7W
/XK9D3UMsUBwyp1I8SDuo68mqVU616QACj2oYpI3XmhdCABvs6k7j8ovRSPPxgwk
jBzI9MOiUa5j2uvC2i2PSdhP9D6/OF7Dxg0eztFiQ6HSeumuSHavj5kkjXFxh8+U
bXA0TX9ub9GxmBSFDhIdOQEjaUJaa5nz7liwNH0ghLrcf6+rLZN+e0SUR2F9RQN4
EGMrvwAlkkWVKshlTFrxSxwxNguGfbAmlbPCWXR8L1tqRd+P2Gpel8KcxksnloET
vLq0CAApyNFFxRCUZOGNQc/xulKBj8nPz+2fIlID1etCkwz08ppfSYDD4bcGOKsK
FpE4xJ45LFIAEd0c03A9Upm3s/h5Rrjt+N8rBMqbh5Dr7JM69Q3nNxMr75Sg6+5r
s+QHH1PeXWw0/wjaZlgWRTRtI09yeW5nM1BZw+PdrB2UYrfryH/RWA2WYMZZi/2L
azAi6KFdvv/xBIp7bBm0rXWytUshcy4KsM8eYY/2HvSKVBF212IFBop393xTwRFk
xDNhvevSGEkxMGbOlNKGfaUgz7eIABDiaIzvIxroItvyPdC9uD/pm5S9vUPP6d2a
pGxV+haAarDbnF9ILjoGaLoVnvKDumQtII3bgcCXKsJmAMUag3nsNj/ymT9/9/7i
g8F5i7FQFm9zNYk7YCAkHTov23OTd30oOLqOYA9Wy7SjcU+82Sle9Y5OSDku21gi
EzCMoCKfAKaiF8iBWR6dXKszLUo4GI3OT1kjMZYVhOdTpSJ8SFXGrxQTLad1aqtM
ePoOF55NarUMSnBgsPuTLEgGKtr8x6pJLt780eSsa4tq4y8A/jIwDJWZG7xJduvz
EydVYPCsOEUQ60KkHbHpMl1JIt94Wv02gjhKHjCIXSxhUIvm8MYOiX3NWFAjTY6S
fjJhP7O1cppVqBX79oc8HjAird0vFvUb1RTZv6iHk3bPm1HRFHIbm2dqyowqwcoj
odHlnifzRvuXUeEeECXDduJx59vWMXuei0s9o6CePqeVVCQFLCWND/7QAYdL1BkQ
O0LOZyEqrpWM7OMXVqlncFzZ/IiqNji0W2CpYh/+UfqC0bWl4Msieuh9jU/VAsHd
XNXp7Excpt4mJ0peZQYGiby58Ih3Q7OECFqb6ktuTFjoMfhlCWhk/yiA/y3rsA/u
dxXY29cRzBLqBrOB95zegzC0lJHDTWKaPlDHIUQHAHNx57IPRWaFl9uDhY367bCj
TqQE5e0NNQowbls6P2PPJpQWiHafLroNDi7Cp/PQpCWuBESy3vluSoNph+hVYZOr
H5KTN/7yrum9la5y9j43nHTfQENss5RZ0JQowues6YaOdVv9M7HOAVxuRWSZqvCn
bMi7upnkI7V9X5Zdcc9kYsncCzQWhM6JcICFxfW/t1ehb1CXnABLvKis+bTR9tVO
Ru7bqUzULsEOgHpDFj3/vZkwEkVQYig9uOaa1S3LkPWIl8qgwrrrk99QC9BJS3lz
/JZB4X2Ufpax+2cjaUVAm9RDOXBLoK91XhAfr7OW2K6DrmTV73ctqydp7njtWgRt
KXV70qx9+8ZLJyNheW8W6FmLsBU1++fXFF5yijb1SX3vt2Yp5tvHbVXLcfs1hWxl
3qRVqvEa976hdmSRV67S5JFj6JXEbR2gTyJnTq2qweX3PLfmFZd60eHDu6mfIQhF
VUjQkA/RaVx32zhzMafWHeU2B/uQMzwaE8lwrsNtB/3LYf78R5s/RORO96BplZUw
D1/JxEI6rJ57fAP4CCV/4owKwhdppMLyGfFLR5lvQORWHU/Ypq20prljXV3qdjBf
JehjgmEYaZS8sGTjgbehtIXWDl4K6QHbA7Mrx6u26YjSq7U5YhnBgSdptmRr0m3N
jaMLDQcVXAwXbthWk+dVbHMZRAug7mMsCQcrm2VCkE4ERh17SpvQYiaW7rBx9fxe
wQCwvv+moBomGqWLjoA3KWqVEXnaIeYH7It+OHn/SvAS0FhT7ugWYymqDAi/2gtk
XzgC5znrh4TcSri3scGgDWIHWZArZy0c460md+LjKaaCPGG9dFz0UEt1gvz6DvHr
KvgIodHMsr85tIUWZuaViCn0UAZ0aPWaKBv2CrwSdUamM2Z2TNEEelqruCl5NUdP
1Aofpmm29aNeFX8GQTwA4ozzC3V4cKqWXdrpMKHqGzWRf9sBgmiCv2s+42ycrxBE
j+zR4MEVHu7Xx3KxeRVQd07lXtM8davmkvRvBPdy9CvWY9psXre+ftWeJnE+NdxU
y0Uo4H6N4+7tMbn0kIeSx6oYO5arMjZcyrJJrGK9tTX9Tc158jzjzFEvvkq2XPG9
HNvjuM7V8wRrxo4prr721jIrE8RJrka9VmQq1y/vJRL3Y/OJvSU4CaI7NTWVHC5b
zSRYjE10EjVv9DI4t980CGWX8hTiYadRoEQHTKzO0HCGOD7aXjRP7zaYFqGyCTwO
A0Y3JeQMywWVkghHFLSN0vNseI+juWho3Fus8lubUz8jQ45p0DhfKp5ytenSWrMh
OY+fYEZNRdvSFQ6JFc/e1Untm8EcsgUXL6sur8vAH37vhA0GqkpGKaqNo5ZNlKOX
GgwPCeRGbanKC3+HWUEtfHYyIYPqRONBTwevHxW3XhRkvMwBFXyAltfM2H551/zG
5tXnle4CKKtFZRkg/aeFlzIAYkLFpn4d0QC9hNlqTewqg/8j8PzRUc6KwW16Ylr1
cJwj+/V4MyYoo/YXdVGjUPRcLtqAOBjVnHln5/5VYbA14k6Ioh91j9gjqJjgc+y2
B2HNK9/Slyq4oqz1/PVKSPHlV+cqZNZXKUOpwfjHXSSGl0HFEXI/mQuMM9L0uGzt
X9GPhFXcNzrDv+yCa6QBuA27K/ZjOY61v0rOVsp+5ID83n7atdNpi78KemcZz1H1
Px9G+tFJCMRIHvztArs6LKD65GPidCYhI5fupfJAVfmmFEG9ZGRWLrjyDJwnP+zT
XenyaG2i7ED7FESmjqQ5FbdQ6lmi0rncwa7rYAb6zoKrEhEpPZSdvCq9hBMRSENZ
qkRgbL5zk/X9cS0uzeVfJuOS0A6qX+rvsBLgxLxoGDCiBLLxqPKgC6NCYeyFD+8h
V0pSaXjqumn5mSaOR13S/+nMSLPN6p+BtR+v/UK6ZzjJrIZgwZnlN9n3bX+iEjB6
0Cs2Eye8YoYZQuGr2b4PTHNuLnAVU3G4lyyaoA5pRcaI0puufwcr0ywQf3CfelL6
hD2tyYRBsosoZC6VM8gkPgxDbLSX0JZDv1hPElMGVgrYLJrPaJmQBpGCwY456zVa
Koe0TkydtEqrx8d4VeTs5BilIP4jQejkoyVBF/aAFFJedogFD9W+B8hqmJwFufQ0
4VteMX5BQiD5+qecIXUY9IFTt7i++B/KbcH2j+qDGljmqKSfQ1nv/hyRQ7NKnbOE
lcO/V/shFCWM4MpCIsWuVMazGf9VZZZadC3bEVIE+IhArV4+EK+YNEyTgAQCUXAF
7dIa7bvuoI7UM0RgKaWVxj8s7A04OtY7QdkBBfHa74eWQ6vuavl19YGV/F8C40eq
ekKWVT6E0J6kwUrn4ptEVTAP3RkfMf/bdgyryPHvpAmCxVqFdtTy3MifAKePVo/7
`protect END_PROTECTED
