`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNskZ9XdveQFideE6jPQaUyLZz0UDnO/iSgZB9i9S5KVDL+XuX2LWz14DPJV6oxT
nN90dT6t08mtHwgGM8nHYpavLBfDOMW80887oS53H1G67lffuw6npZCqrzy1BCsY
GAbrolZQDR1gWFyCJVKrz0mguBEEq9TnQKAHxYBe4tryvipYgMcaH2kwVGp3KJU8
BR1KwYftBj3klohzoSFgmvvx0IYW6lbgqvz/gACmnmxvMCAbrheNsKX9JBtHADPv
AM9ZvVwJHv3f6cnmZ4J5qB5RVZDg7II/JpB1WRj2LOmkCTYez//jGzQovSxR879s
aI9uo20Yfo/c/FG6v0l5QIugcb2ELw5W3DoywgYRPdLbMxUwQGpz7ierS3IdkmR8
fgqMHObjewov5IiX/HfVJqLETgmbxcMJQ2CA0ro58xJYa8kSAPXwndmH4/eRYySM
V3d0F/wqdnzdGDIi7C4P8iWB7o8X2+4OIDTvliaR4RbkTjIL7gYTIZCZDvgOAX9O
5Ipc12La9Vd48m7WJirT6X7DnuKhyGf8ekRkRMjrWQxL9Ea9gDbSmi2lcuQIWe9M
uH/M9p5uOXvhCik4bzWVUGxHhaxUC7hF4RNOJ/76u0DFeCT1jsfF3d+YGTx9rd1p
YEExYtBcqNqy2r6Psg26zPd+MebwbBqBhNa9BLD6Z5dgLILDQrdY17OzsuEFVoIZ
2ZBfHmC3TFBnQIXBSZfQQEEcjLWUVQa8DF+Uuq1/n4SiXiwYXOTkA7mBKiuPaCxn
9JYxT6lIgelMUmnbkQR64XacYo9cWYT4SvYlvZ1Y0glSiSXAbBJRxM48GqiTW1oB
jnS6BYiH0tV43Xl3MQ5yWXB8ZeekCu7xigenCkiT7YII/zYM4uTIduZjP0m40raM
fw8C+f2jTkwUwOpC3GyHcvO4BXxljF0+T5OekIeobnH38vn/SFlLIaw+IJFNnjlG
rSPm4quLViXZSW42b2wv/s9CdECd+osqCnTILfTYVKTSZODEkubLN3EyuVG0kr8X
wdVNY6QPwNX+2cb5O9fA17TobsjMhwUosjzIgzzV1yEa7tdwy+401p0KqZ+vl6UP
9yA83BUvpQlsefnlQpB0bMScC0t8BD1qjjVJkh9VMPoCnD6YSw0w1QjdYJW/yALg
y/juJEyjHOwMJUELvznJ/m3KQRyzzJEudTkEFq55nnGOUNbwdgUTmmwzOpWTDs0E
tnYTSVjTgFuI31HG8R0tw9g9X7iEWCHsMwElewvbw7nLmH9Ir07BBaidLcEeqac2
PwjFAxiFosta3pGPJLE8l1bXEJsEDjXtGJV5z0WgUr0/za7i2VLoc7vwPZGXf9jj
Ke23kZvnFnUIzc25zaUXiTRq9BQRlmI0ZQw73oKG8zHBYX1xylI7kiIYUxJOyGL0
G1Uup6wbUJPD89Q1njcQOFQfsEnjbR7TKVqzJwH4d9uVj1ApT8O+ryOvlfVKbceG
BxQe7Yn76hNSuJno/gQv2lhUi6j7xZWp9g9+qQy55ySw32IPu5z8pIMudQ0RZhWq
PeOMsM+38HJJvS9VdfBDIA6e+pqY6cUxSRGJB420xvKj8R/YO3r/KNBsmtv61kJp
RYIrnTUL240i+hPK0A8v+/BGZ2+rjNGAewrN7XrIkWdbJ2B8e7EjoiTaEwfGqUcr
wAYu8yBPVFbyEj3On5HxXL1L0mokYRcbv8d1D6saJV7fuGwVom/A0k8A1vOQZXwO
ZbssnZCRG3mXt6QLHJPwvt7Loy26UjHP23EJ9WJ+VPI0MbZLF1+j+Zx6RFF3LNsF
1Kwrj8jbMtV8PxseQcEfp8aC5ixjCawh/DAAK1ekYeLsD0yvWzejxKcZc7DgFPZM
tO3IX3eYe+sbCGpIZ0P/RS6TitWP+3QGjEepBSJtWniuKwHNgqokMMTHVv31NPTn
XFyjl+JLykcaVDOA/LkXERWFCBl+5bkFykJPtF7e6ptfLWCxoII26X+RLQgU/iIQ
Bg3eaGwJtuk6A7FrwfxfWBFme/bXRjOrK6/5NPQsVLJP84za6BP8JNVH7Prthcj6
ciPEhJ0tgy0bPQZBkzAbXX7p6IQt8fgvQ6ez9GupkeNXHBrBmfll3q+8ns/mq1g9
vv2oMCWl7gb7pR8pg1hkQkC7R9Ff2f1t0238kAdQhWbxS6PflLTqrBzc+t2oKPfr
napUq5WGGhOUvPepz8uPzB94i0eNs0G3EfWOPy0U/pk1dXeKUnl20vYYf4O9s+kG
/KgCth+D2P5RYrNnqKMf/3UMGd0stJcTgQp6Q+tX/UZSlcLjvqpg75kfIi9LBz9C
I9s/lq7FFSnBEf/NS8Jf9w==
`protect END_PROTECTED
