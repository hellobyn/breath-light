`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wC+P6NEjts6BH/F30Keywub1LkqU5iFK3IomNuWoGrDglkPNgwjEp5sIBjM1hXd
IZGLth+LnG2k9HGwjnCoXlik/63ZjPk59nfcOSQJ1vXMg3Ql1YDIXhe3Xzln9LJy
lm/yLHGm5SnKa3YGFnWegw3/npj/PwLigZyaUGcZObX5mjRI4u/Yf8nx/pdeG2D0
kFVNdYVJyLhFM3moerTDt32/gF51qJ0Yvhnr1GaDddm9+cmwX7AAVctC/ZiDueS/
DWPyevLGgLBXixIuhkKJc41xppJqQW4zz1qBEvuQdO26+ouhKS74ZMtzJCkPxMnB
ukI+6KyJ4XrP9LAJPxQlY7GSCk9gijsb7d4FCCN5Al5sV2OdhjHdudxxkp1ewd71
4Zzoq+grGYUqWwrMCfmfSiPMf4ZCeJBp42EEkkE6oI0zSMeI8fGr5kvdXGWWgx5B
LKGJOQASP3HrmQaNV6NCfQJtoz4JtcHWQul6ldnSqv6LsbigDPO1f2Jkz2kl5IPD
YYEVmeR7oMzdpokwUxLbrhDgXsiY9DrfTJ5I1uCCMv/7AGHeSzRdH3wbnCmb+6+M
SAAPG0xB9BrlTVtpUKj/ocyBs9fZqDJ08vUn4WM01sntQ2vTTScipg9hZNVDHhFS
TH+e1TSNluyK+LdU0MdsrXy9wJAaHtgGrmi63RfRA+oyL6xuz9IkLNyOiWvexCq8
FiBlyhiPZSsTIwH0v8617mn7aooeVHglTPviaVH3TvzmGoK92QYKvuku2VjSgB66
hHPUUAf9eLqAflvZDwhoXVGa8WNS22i5brFLzKqe/CcISR9MoM6HYEkszdVUjYu/
XPc1lK0gLcVr4/N2V+BO9JHWbh8dIF4+2mutlyv6hXMkfI34Z4BZWsRKYzCvaBfG
JR79s6d3ywZxJsbmuOPKtBBS10L4N4xNQpp/yv5KJ4WNz0MIQ5nIbvSYS25w+PDS
Dmju9q9Oy/l92xli2qagfyv4lf0NpqaCkaFJauOHEK26xxsAi1BIau+SBHK0x9Ct
E/ddZvQHNOJ8nKLSbh4o3YkVmQrPVd3wPc7YMQ4+xHboR4vAfYnuBa04e4Iy91wO
Iw7VdDhsdZSj00a8/p92sBIK5VwCPtG55OYEOzvsrNKGYKgD9genjh54u8Em4fUs
Rh3QFbHip0qNkKbdhRiNhg==
`protect END_PROTECTED
