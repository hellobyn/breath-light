`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rKm2uUMNYQIJ4nMrnKLa/v5an3YSBl0o59AQIvHyNgZqx5dRtPEvBRpui4WFDbY
hKC5rS9OFdEZTBNjsMtvoHHzEyOCYWnpe0dLy6mW4y0hOggSfqzZywZMfbZiKSw8
PeWT92DxIl2E6/pJfIF19VMGcUm3b64p5YkU73FJHqf5Dpc608q8BcOCQ1ruOa7j
bx/hoFP5kpUHB2AhBBOLY/YPftSY5AXZ1uNAwlQ6kstrmEKDOWtF2suGyFZ4/5cN
9fdkqmDaK6LelDy1F4JUGXZ1oAbL2hnPnhzhLPhKxi1lLN89ds1sl0zrFHmkHeQi
087pxwYyuOYZadeAfCl+zXoTxaVzuFGTNKvb174xFiO266fCe+cY8N7G/rsmMNWH
Khn1tVV/FBoGpyKqbtbSpwQ1aqQpZ2mnWnFahyIc4BeQgiiE2iUVxZZt8xGz9yI4
y3bIooStln7iq/ryCfUImNn0Pk6rOyXaG7CxlUiz8UOTMUBRbiztId1sZVf7x55U
vGfUk/3/GwXK6hBq8SV3w5jdKlVxQ2UXCIPOO3hFVmqie9Kajiw7BlZ3AiQjG2OL
SQmpL5pIkvHLMCV1EyBtMWiztqUDGsNENCdxxhdSixy0+W2zAXwNQq3jELuKX+Zq
92/OFhQ3Mqo/MXpB+em6e5nCpO40c3MVD1VwyBUi2l/toP5L1srLD6M4IrHGZqHz
TFMUOM6S3vJbhQ4sc5xHdTUD9gMjC1nwZL2Jr49eZWUxjDw8MFTEFsKDhxt6kbne
43I6HC5/tvSVRbuQKw4Sg6z6D89JD/oWokYE7/6Ehn/KVtHW/hSOdt7t8ep9bDFA
ncQMFRpWltegKU40lbkhDx0A9ag9k0r+AzwLUucGJJwt/i7v7JPlcyQHVA1gyFnN
HHn91x+scgqYs/04Jg3CwYDqgF/s+KaEVo6aOuN7b5Zf8YtD+PgqC+juktut7a+Q
ViOdXNwzxskivwy1VhLUOAYXzYHiXSND7XKDwgB+a5MZQHqLiqQRU70vI0Y1nKgz
qHTqpC48cn15cjzLx+NYvX6y5Q3tD93wNStZ3VXqfMT0hX/n/ve3LkIIkUW/BTLH
mSksZr3/LOQLjF3CwsnQH+ov9VC6INoN7fznmugvhM/gJbxWWdsetmLspDz+4WQt
lhfYQW6qoepyq0dVV7JAiSXsHYka2TNbp1BW/tWTxmCkvrrM7Uy6WoVbREokzF7D
7qIYqz7tZaTWvD+mAD3XZIP+/Ckcx7zLqJc2ck1IGnX1gQ9B62/ywWmPTKFWI1u6
34+nO4D7ud8GTylBCkKj8fSGHwyeUB5/DdeqTWhDbjpk1DiHOckRfLaJvXOT1z//
WsPK2C3IFl09Sp4LDKhludOvGllDpCWEHMg5kt23xKezEWkIHEYuUgwuHRQouk1F
cl81UyU7GCvL/49XfHNB88ytbk1TdEI/kADVLJ75engiRxCjrYcvxmTkbXA41PkK
aJ4Z4M8piJfBDS05xMosMw2kQWfG5Q9YATQOXqXp6sgU7QVaRlE2K6cZjr0BYDO1
pzBNTjoRZl0Sz2FczCJqAJaqAol4Z4IomNV4KSew39fG/V7Oc50kFTSY0fvdewRC
1B1rh1R8W1vpJeZg8Y7nnawfWHwcN1SXr+2Vfhbo0Fj6Cs1H3iqsVEO/c3VFrlIM
GWJrDBrptSaLt3baA9dGLJGfLTk//TbB+l2JwvxNwIHAIm+bFmqcotsHvylAQDcV
zBYKX7u5bVPiV6p9zTQMNHDrXC8bXREHq6zSBUkjU9Rm32XA7bbgtNVnkK3lyHIt
aou7XaT9WC1jMFe2ABb86S25RxFQ1DHME5h1ko+i/niwqMYHqj1gspSXpNY2FCzT
QEYKCBKKaFpnR4wRXlFzS1Vap2/fIq/heKgnzAUZ0WJjRhtYG+3Ak4DDJCDIIdFs
Y1DQZrgrqTxMubOeLd8bWBxDz+2heRv47xmh2e3/Y8Gjnb5MsOs0SKz6keONxLWD
meaOFh3nPBkTMq2P/oPgJgOgh9h3cXj1CmiPKjQiVfGpmRyrN3X2ErtRefwvCpQG
Bc2s3B8bJXkC2qmPHL3C7ZHhfY7i19CjOjlwt9nJ8UGh493U9LB9AeFMJEtc4fmn
c06gvhIViB7H9MwidUfOgGfzEQTW6bHShu2QV99lK3gZlfFPOJLCIxZBYpteAqaK
knERAh25PT44uqewkKug05WafIgUlGxbVPW5fsiXbEQ66CC2gq1XUDhxfHF0yWzf
0A1H6EW+8LAkQ8d+/a1DkWobUcgkfsBmYIVhKSkmwyRk0MZztcN+5XKIEQabHrMD
IBsZdOdNewy9yBNQkh8SWXU9NxxSJgX0gn6JC0KSj/xgVUZn5yA5krNaVfxvfiai
UoKTH0E8cuRqWzUuYqig6T62cVXsKhp31TvkFKS2C60m53AlR5BZjNmpl2rrJUYV
C6BsxKOCqRcy68HQQMsuUXIJJpAKZ5zBm+ueVyOKVjv/Wkyv1avmqbYJFUuWpDuR
6UH9Rh8MyCf7nssU4Qj2wAsL6f0TZodYxG8Kkko4UCfKqqw/kmfp/LaDGmp6zLe8
bJBIahZP4AkwIY8XWwFWVe8IOuGszGpuLN/L/ijhBEtZ+LgfvanUgGk10LkmYm/G
1LYoc+qkCftphoMhFUhmjZEgsORVQvua4uDFLWblFVlwx9+4H3O3QtWOH36woOSa
oM3oLcxK27+BAcyEiWWozueFdbszzeD9arSW/X3Zj4kjUIx8FNl3w+4YvNkXsi7C
RVXvUuIF8m2sziBQuVN3GNhvQnkqCd9eap5d6jtGlD+1wk5gwlMo/rTNNlxzICtI
vK58TxkPnO5+UsvQOGOV0sXgB1xBAFVKyEJc+0YdguVjEvUXd+arbTmw6LjIVIRM
xsHXSGdTTXM+HDQQdHOCdUEBH+G1m7ZRLGemyI2o8mxG6Lqi4RUEAigliSmOUDFp
n0I6cUVpGucczi2MvUy5jKnT4yeY9CJnxfGVF4Bhztkyb+60GfP7kXkjwXa8h3nc
Oeq4PQRxV3A0w2p8j59ePlsc/RKydLC/w1MlnYFLvM3wKbWro3jNhjsglMnu1je+
1fLghORRgcHsaRYaIGDkxdB7exEOlRlaV+ztEXJLVQSoXGojelX3fjUQ7sg3uGfS
Cnb8MSEtNpO+qhzEimdocKHwfi6nP61NV4vOj7WtpPpHtv875q41qPGVdLlHVgho
7AwHYN7dRI0tK1cm5L8AwC3eVkAE4hUslR6sdOo3dB4VR2rifnVDWJCe6cfFchX+
qgTXhiwqGFeOClMTI/FfOeEJMjsvLGFiWXK6Ee3HKcDT3ladjjndBGaiVXXWB3tx
YQNQMmdSxPwRp+2E5m4l/o6DiUUj6oWX4e/GEy2LedNaRqvI0O9IGBHXXzCnN6ZT
+Ttt8OhtxWGR7bXNHE6gtez01PdH2uJAz3Q6DMwaa2/xMatXHptxFWtJY6k8r5/1
Vpv2ViycY/WFO9QFKUsQiA/A+WjwH/k35q0rmFxNveT4Ajdz6KktjXVpjqoWb+EK
ZzpyF/skUtSoZvzMC1CaQ9+Xd8E3KMjOWTZnmtodXvqWdbeguXbcG62lXWEUo4R1
NpHq2rqHO1vBmRIwRN3b2owm7b4WfZSnch0WSZTzKcT1cGNv2CzY+j+xXUd1+BAb
Pv4xXXYu9qtcg/WPb/1Nkz182Vd/2nqIGuZm10ggON/iSjVNa+z5SO2ZS2y0jNkh
MfYP34QzQEjNyVX7g8UGFBPLVhvYyVrK0blLKI5T4JMHfK+47cxX5Q9ydOrszF4j
7PWUk55UjtIFWfo8qrTm+Bl6ywXmJd+DdGmJV17zIu7apYslJ7TRv5TzjWd+jjIC
LoNkWqhlw+6gYvb40Fz4p0RXKeHOAA6gu9umWcdCoeAJZ3sHhrktm8qMyaGTRm+J
SOxkjHwIfm3HgCynywXqFokYYsgXwH3guRLiJdqd05mc/GUimUtXkh5+o9DmJZbi
jA7aWOjlA6w1kVWYt8BwNaCw2EhLuYm+wFHkwV6tiOAgkWgAFkV3k4RqN39z+z/l
keXxYw7XQEYc0PFBP+VetaVH9TZW0ttwfN0ESJrJ64sJMPd6cNCZU4y6SXoCJ5jx
9HDPxTEU0E0Gv3n5df9TmYbUFRcE8VETlb9a3Wemvd6uil9mcghEXZJtmUG3wz3Z
PNt7IcffgHSn0Pvcl68fUYPO9PYfJXklIWw4V7vxuryXUH6M0WB1TQhwb8CSZGj1
dOXudTHB2Kj52Y4qFgrODALNqjQHT2R60chb5Yf3/1K2XTQPPLinANCibkZRxCFV
3BqsWLxRnK1zpM0VrhWM30pSAxhkUhBEOkmS3KEc19BW72nfft664B0/4uEzfBH8
mMFPNQ3osB17ydZFhjgE62kAp4ObKiFW2FYpui38A1YV5u/aTrhc1HGBxKZvoq9o
X9foSBSvQf+9derDVbZKPfh3xpxGtOEp+82ZF2Cuk2r7eeXWKpVpZnZVOqc4KDgu
bOVY/c9tHzknQAcCY0BhMeC7G0baYgLvjrsYfjjEjOPZBq24uDc5lVsTZCeSY8Jx
kiXhaQ1Gi/yOYxcJhrr55+5kTgBHDXgyf74TVIUXZaQ6j4LoU0Y1JqLnwiS/+jaq
vv6Vj4J/SOvto82b2poPEQBMls2oey8363JxbxNc0x7NmotHP+tfPmeOPJn/XAiD
J9Eo4SQLnCvqC/lobv+iuJu//L1h2B6dt4SwoesbjIv01lMB3qw9k0Ty2wpzXdZv
mstnpmQvu1lRZtItmU0+bl3l2lajxVJOvM30nVj2V7jKLdV93NyBoUFwwM6hIRW4
FBYq2TbsywloNG+wvB7y0l0azRtW2GG+TyUKKYve9FYEdHqE8z5opqBcuBlACslP
YdO19yuH/TPC2adpE5u/QEFf82/v9oCKzCHpGivMrpON+/uwFQ6hF886w97BUvMD
bg5JYEemCwJV4gXmq6iH+q+T//b45KyWcxXxPoSje9/ISNSxvq4nrPO8/YRxEG00
bbXERTPLfC2M/pycSg2PW7AH7izYJgcLhJ+B6xBvFmEHBTSs2coOGmWO4MYZQpnU
9x1s/l/oaL1C9Fod/xwB346L5WXUAOw63SKFFPRB9o2HWGFsrzkNwrudBax9948q
stmQ9kQiWeccp3XgV5HF1MqhBBWfthWciquy0aDFcGb1X3hRgtl+8ocnojI4u5cx
RtLBXzUyrs/ACkl51GI0ichzaH8wX7Uo/P3k5RUXzUdriu65FcTNWxpxzBWwXn3K
LbJ7k1WHIqF0Ecu0D2gQo2gPvvJO2PKGC1pQo8XzsnajT3ijeicKccSMWVmGhN1q
QwN9UYHqs/dlrfNL5ki8JLPWZWKs0FsY0qa2B7darqI1k2RvDiHxlw5uKNz7e1WJ
C2Xh84Bp5YPxU5NgmVmKF5KgzoTvxMtYOYzKJ0g9t1GIonfjLcuovf4iUzxucz7E
Rq27Q2EuqiIMBkzRiMhl37rPXzuUrYz+l5QZW8Oi4VyVamBwPd5zgNDTiyzYkPy9
pnbBB2UUy2qsR3Xi6Beh39n/MWGcrj+EZapTS/J922mzEr/JaLY441qVyvu8E7Nh
+2NMyeECrxUeBUjyVVYybqQqTir5GveFVs/siQsHG4/rQS7FckIw1xU2CG3OyuT7
SwM24WZDX7IP0hp/3dmgRvVY9rfuVktaru/VaePwms50Zh6owtpVZReYoy4SiBdx
WUZNQVdciC8sIVG/uE7wKpq0Qfn5PRz3xG3bmkqpGCamiE4iXRbaZrhWzMZ63E33
llexYR5yXjXxEsusKTwm9aLLl2TcwD4oCuyRHtIX4v/CbsgXMebyMVNzizqJpn3A
rPapXmXEPOcXZbuCZtRXU67wXpzdlduFvchz3tm8lWd6Ih4kR4ZUufeQWhC3Dc0L
tQ6HH5x9LBOG3d6Sk6BTSmLrh7Y4PklXdpLTJQwcpAVEoyzaApzxN1148E8F2Sth
o5vt6FDbRtAVzJWnLMEnV2g+9iI4lOwywLv2eKyGCtjdOk9GGGeu3N52huiX71h8
JEuCARsaaeEUH6H5nEfc3VmcqGyk23QBugyHG/H/20TOcZKkZjgbtsSN3vf7AzLG
d803mskrZoPhs8bgBHpnEkY2GL7jRR9Qw/Dusy79gz5G+i7jFcsEFSxDo5Vh/2xx
zT0HE0dE4A4rO7DMYY32z7Pu/O1gwPWCkJBIcFoLednZmd6nKCwWB7R/7iwErsXl
JSNB1MWQt/lgNA8fFjhXA1U+TmYbi5d3Q43ylZ9FwmdtrvF1kAxXXlOeJvz74FZg
ljyU0D2x6il4rCkHLQLfm74tO/KZFkV0W+0gklQrCPR7Xr2zU3C7ryjAMo/DGBpB
`protect END_PROTECTED
