`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNqhmueQSXdoFMHTSczjex+MWsHD8INyJbjwORdq5W93zaTgzYHMx5Rta7zGjHTi
HfbFK9aHFBI5yw+a3TdfxU1p6v/FTmbJOBTutDGCzpJ8BIru9SgWeWnrilNoXUf4
w+g9Hd7OuXPIizTjP3V2gafNEkGcCBTJcV3nGdL6kzWncmJQ1FLcf3PlirFrmrgW
nQ3tGTFQjOeIK23fBGQsp38GeL9HU2kOwRSf9+kN7t9KZYDkm7U2vS9Bg36jiZaP
jgg8PJNcgr0S84BGGtkcsUFlUxTnz9umeubst1xQZIrflW462TrAnbrc+M6FzcNl
sjDhA09ztkNDYnVDWSDQKl93gNWhdZ/7e9fFHQNUPgaj4BL66YK4cX7aQPFz5ZIn
rCMUrSs7gGYkNHu/Y0cnh1vw94GvLtH9vBLeKi3jBqZxA5EPqeOVq49g+4m3Na67
5eN3lDPtVudApM4/ZaWEX7quLCn9GcKlN9CmkRx4TNZGtqH9wBRVlbxWuR+hMTu5
CSFxGmGFwFwSM69H/6bQR5UscMkW9XKT4XVLSXi9C7TekKBTBcEPOtnWl4km7YEB
pGcj5QadBkMDqnuW9zI8ZCgYWdOCgWVCG9NNYQ1zO9kIGb+rFH8SXtYgyFClMq0c
roh0ZEvhw9CC6ApS3pZEqKuNCdVmqsC1hvjqXQrGzGB3N0JBncSSpYOeniwCQNfj
yNreC4Q9LbKekjCLSZFTaYCwoEKPzJtefhSkOdfRnXhDyZzakE74dw9DjoPEUvgV
DGXE1APmHQ6iBB3eQLAr0LCIZIRDezVo7XoeU0EB8Bshs7KL2Xk6xZiAu6dQnWB1
M1pyQj8exDPY7icD9n9Sxs73Ps8LGEovGEVDzm4+97BlJzwi0nPsrlNJgqDpI4x/
S8FW6wPVjavC79MrSyPcFAdX2M2ICyId3mC2odTR6Q3q2egM+cG1NN+i06CQ4ahi
4Vpg0N4nY1g/YTJFoncyrbz8mF+19ejHWVRywDfXVo/AQpZi2D8S/t2+k5KsNwAt
guehepqn8GtByUxolGrwPCFLQqrTaSOnThlmRJL4OJ3AjtSoFXGe6rshh+DzSyPM
NvDDVg5RP97BXT0kE2wuvuyGV4FqnfTNWVJVlJyYhU6fO7dHfKcIchlYqThaWdip
Ldnj5R0gK7/5vG/35YkMsWQ24H8TKq4Zxn/fKhRar50ngPqmQenn0QuTXVRa744F
4aZ13HzDNxv/+Yb6XWJzO1ZjPKXb4NZ4WKocc6pwdAwlAFf7VKeika69L1L5N/HW
W6/+Tf71r06v6tnra50nSnNkbOgpQbqpDg4T2CKCWWJ4TvFxY/UtOuvxi0nhzZyt
T4uOM+1ce/T6jAGKfXI65g73husPU5/gLDnhWazj3rrVew3M6NX0emF9YFE9lrQw
PeERaczhXvtW5a/HpB8ed9VPBIp4FCDUSLAlqHGtbai5iFtO9XoW14pKeW2saPI3
unbfRRRMljNehRxCzhJluxQpaLUAkFXh+Dna++iOVCf64GY0Ds39bBGf4roh/X2K
wVL+mtYbkJeS7+P+uo4ImOHnU9+Cu88AsOwwO3smZUID9ev85PgRpGvGaXt+FNnk
fjIStd+Ca8awGHbx57VrFYpKTpmgcVKpY9lpG5qAw4n+VlaxabCAwy2HUKbDUTud
9Y+Ek0Yx2p65ciN7i6g55nhotWgrkbsjIxu8oKToUoj4zHExew9zrVAVN1xkglcL
nP9kf9q6l3fP0IC0sHCNWSe2T+XSjLimgDUF+1buM48Qe8DE16Quu4V+n12ffmjT
M+2pbCfCUDcN2InVc9VpMCLpmKLh+BqmXaCsL2zW5Ztm9HuPcI42XgC6P52mD28f
8s+96DtYBfGTR6ANMFzZ9fo731B0R5ZrRVCQpAA8oaHSN0KgPlW4FJCqM+CBHlxR
vO/4DEnzMkjxRoC5WDW/6zoPnNj0YRz9GhAPN6i9+jnllbbY+WVhqWeevESXm1kr
y+I7a30ker/8+nz2o2mfSOw7EYteuQsJVJFOWLGvfvswyopsvn9VSmVtiAAIE0P2
tcd7CgVKY4mBnHaCuWpI/pPoA3dFXOEBNogX4GTtRyqO9TsAmrKZPc4zJ/wbSHbx
mHL16A3e9jj2Z3A3PlA4UGf6l45zuFttYvyBigdolCEwOzSyQ2C048ccGn6/Xkwr
X3LLrebZogz63muYosF5ImDr81ZiW4kERGZBvJk/qMyKgXxOcEqX7C9FyYd+iVYg
0Dd2ixk9JUoPiFh0mU0CMQwUP0RUbspVGCateEVsD1eWhfHDdslxD+mG3ZsJ1YUW
WRTgV8JZnd1aVMMkUs3jGrt5S6Td4p1RarNbbo6keIDDHr4wZ52zN1V2dH9L+PhJ
IdRWwI/hwTu816SPAwFGQJ/VkDK0QrW0M0Hzv+r+flWGumymI3OWfBwNPMmoZPln
sB9WVAbzgx4Bj4feFzy9LcFMIrrezodeaS4vrPwwjofGwB5PVytme5KuzgkRG48Z
pRrFhz6mFPgOmxb8lk0OGkvYqZRbtPW5RSVwl/7daLPN7UzVWx7S28EW9v7FUAOS
ZEs57f5qn1ztCYMG2nlogws/hNbqbjiMJ33hASxfv4ajO08om3IuvcStkIpJ6VtA
u8YTi/dlWMQs3vz7ATkaEAUYF3DTSDoxg60rg0BCFRdrw3A0afbqKdybZCLfkzrw
NCBtGsZpKb7eNcFu+487azT36tM/b6vmSUk5c+lxDtdeHr9APj5h6ufyC3xKoBZu
U7blB1whiPsblKoxEy6bJdbtYnVTvU0X/IgHVYwWqHctOro1cWb69roTjrM1azzj
Fn9E2xnK4h1+JutsWI+UhFbGbwpLasOBFwMl52W/kex2Vmjsiwe6ZVR/bcW4ru3w
nnI/jHcXQ8nL60lYMyQH9TWRFqkgNp90zVBpqL55eLfJrrq5oOuEqUFFTk3BK24Z
/qP/AG4gi0D+u1TPlWAug1ugt5+JButxLD3NMPk0ckmqAy0pPaexyjC/Jth0qIJW
ABccgwQ3TcNr21lgIM4xOjxYh93XmkuSW4fYduCO1Q1d0XnsvLoZrgv9hn1Hf7Eh
86qVZAr9cdqmVsGJ8gKp3A==
`protect END_PROTECTED
