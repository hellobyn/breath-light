`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJYSuNAX4/hoAnekiKg/Rzjr0nTVUK9bL3saPteEEQjvPLV8+0PSgSaMfcWKE2P0
SjR3F/ZTdZtZ2soLw9YvxwQJw1PvnbKQdo6XCtvdvOP347Dp2hbUifP3JAkZomB+
GY34D1M7kYbDN7cGKbP5bBLYn+UxVCvqNBVV5mDxWWvAVb8cEc2B3fYjn8FpCeSl
PQhiTzqRS82PudwUQouZhusIm9NSMPHaIXH2Z+PUe75n0g3DloSXTCxazbi2hHim
vaHMFCtr/9We0IKCcNVW6cenmJ9oqp2oVmGzlmxbwG12u7WejwE/nJLGzweKHP1U
QUtoluF+Annx8wvICpSPvNbW7zD4x29M5OQub7A+ACrCnBEOZK/UJUIJPvQDjNdo
6tQOoTuQkuxePePhjioQReY8rZZRUptppEfK5UaNBlGmmQrbgzyYIymroxijAVTm
WjO24D+DVTPsqX2i7+o4YmjoC2j1DyzU7wZAeLVxiTly+DNsJ2hrmfLNM2Lzts37
Slcfake1nyLKC3rRryE/QUUMSKHdqGOSteb76EXlKZ+uFwIuM6okDMlfxOYyvh3Z
BRPb5MX1cwYw4qfFobsns8ss7F0LOnhIYeinBmyzqyUcd0VMiMMj3XFJMLi1Tcnx
1bbVoP8HfoYkLroH7Flu26LqBlI5zgTei85FumcpO1XgssdfnxXCy0iYcEDf5gQT
z88C9cgS/IFieYm8tt9NsSds2GAWBIAgvo24kKlfRvPg28yFdB1rjHGuL198FgH8
EDgKaMub7PlL3HOesGe3/0i1Dr0vbTkRuS7Q0QBrG7UNd4BEkAGVTcZEn8DYpooJ
HyBqAUMvv4MgZSx45e0PxRHXvdqwkv667XT/aXsKu5g=
`protect END_PROTECTED
