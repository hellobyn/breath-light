`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4EIBo0XgDZnu6E+O6+LWxvKmQm0mYC1G608dFb9acbISXj4xFvV5AOd+YGBRPep
qCZs+F5ZBf4iCaUcRLEw6wIEeODU1AlPLn5K8aDpeNizLngDkqUdQXqoxHV8d02I
4wLZXTS4xCncA5mYT8qvPK2Vxir5R/2wStiTStUjkGxVuRjkijuicYWo9V9zUah/
CQx8eBNVW0JUIqyCT+wdFhQVqT0gJLw0Wy90ZNTpquFXSVLjQuRHLVoA+pB9N35C
h8soxyhzSf9rdegVHaFvkKrRubxF7pFQao2B5WwnH/DuK+Q98GXPrVS8hM72pCWV
dx6qwW7cWhedKsjJzT0c0FIWzf8Gt3uukEe0GLNCmRQ9vMmeSJFtMovrwbkbTBf8
Oy5vGq3QpvWBt51CdZ08NmP/yWNnKuKe24Ywpzwzc8o0Unh2p63iMoDgSEbUV2TW
CZ/0kip5ob3MPMcPoG8jO/6Hrp1gqs7Ng4hi/RwvzWi8m4QiRIyvoHZ3HgMVVztd
nh7iyKVUtY4tkw6favoCTDSbFAyfz7/Xle+xlgrv2YkGYqCEUpmFLU34UtC2LmlX
yvX1jYxf30mNt49T/UofqUPPAuJURJESQcR9Zcy4Ua/tsATxsYHbCQbR+n1RboOJ
jqz7a97hjMjVrP/9ftfo4HEETFoG/fRBJlBBAMEAyVp2+df7zTMsIiuuxiBnDJ6X
6ymaTaU1PA/gyyPby95iBSvoK6sZAgkO0athDR2sdgIPwqVNMBOe6hembfJxBT1t
S5aVfhRDByBYHJkLc9dfWLweDFI6MawJXOrE9dUmK7+e6mmhJDfEzXNgW2E+sGED
s1hWLO84BpzAXSFokafnch0NO5yiesT1sQ2D8H2UP0HlgV2XYVoIT28VwXicdo/i
6uB7EMCNIJqTjVfUzX+sp8Xsazz1aKLJ+tSUOXP/q47zUlq17nrn+yN+IUIkV1NJ
FKhSLRUYcMPVsTocXK5zAJMu4DZoutX0sWTXJEC433CBdF4n3Nzne1P6T7uTY/z+
HXxe8nQZbs6M0tRNaVO7n1Zb+uMyqhYyWCvyHSDEOEt7rZ/fZigtj/BrqwboLYgT
uekcw2GMh/bXN8zBlizQTlsj6F5iPL0Cru8BMGg5CDH4EC/dh30Sa3n8Pebl5vm8
4Eay2xrRgZBYXU9Tiy7/mJlwPh/J1dXCl4CcOW8zSQVBhCEyCrJremq1xfTE72F1
dDIfQAOCw3JsLHxctraRlw2MYDg+pVbsqtS4oq7ktysVpJ2No6mOsQlOiepsZval
XFkvk2SvD37qtNug71X09Z4nlxCGOo0O9CAteJHSRWrluHQCOw/JcsbMsXixptf/
j3+IzVScyEp0ne2+uWg8DMxXfoN3hTxlQtWamPjMOSczuOo3nVZFGhZxxNQXxuEg
wSJYQWuVeXpXLD+JUyxxNEwzRdiujPKgCuSo4il3Bi31Vt/IKZ8dvzgXwr9LTKLZ
s86PaHvryz2O6/Oe6suU/m9NaQSRV3tMZUe0N6w1myhe7/PlGeB3jvs5z8XIR/IN
/VoLjFjFIUTI7M5P8qHLRBS6vcToirjNEtVa1AtUrL8FZbCNk8fVoIQKaw2SgjP6
OfHWmttP6tvEs+au7rVtOiSQLbgK3qVfgE9GCHkU8eP9ZIwMx4fqcMrjPJFbMmGA
I30xvsKdfVJ8rxLQbkHw0psNUZSI+GrO7s3MQPx6me3kU3tT7ed1pSK/mEqZ/fDE
d48Y1XVSyud8dtGRPFr4n/VZPB8KfYHNYlyTFEgJUaILB/VzJ6KOVKlGkZGkyI5R
KyBUSbDLpPOmUQTJnEFp4PZV/XxuIVZtjTwMMb2KtM49PJ1y4c4bBzuNoAvA+Kzf
8CLZB+cqGrTREiX6hJKxiGaUYqZML+mdH23aO+OJoQFGiWSSce2duQt7NhdQbh/F
PMIOp7+TNKNb/c3GJoWXB4tN0iLHQsi/QKr2mVk2PjMKSJoHMhGWjI+wN2v514la
mGmF31MXGwYOqwarZPwkogT9f90Hm0rLtLV7Wjy9FdIVV1b8xDX+N7tnmmz1x6vx
/ucVF3lRkInV86cRRStyCToqpqAeOCMjRq+AaErirQ1heFTc8q1vzLDppU0BAoXE
UKbxR+ULdh5eJQxT5zoh4ww8YS3Y+dL04oHQahbnY4hZLebVn88hX+nCq+uRWKbX
e2vxE65zmMg+39GzraPuEM8f7cWB5yf/o57X+RfTvat1GFJi1OMobKsLu34FKV2F
3pntIaAK2wk7g/577JaJwPXaXtx7o7ff5rk4uz39xerQFSZtByGcYQuya9wSWwJ8
0MCzIL8kCL9lDRR5dJmhazrIt+MYCXKCxSR3tqCnj4pEd7VnwdDq2RHc99vEw/7u
41YljG+X92S57Fl4AAVJjfcnpyQcxEvvgQz1jrY+/lfSRzlSmwZEwH/agY8KiGth
dzp+IWQ2CeUt6cJmweaDhyUNugjG3fT/LA2+HFW3SXAqaNE5vRYDzV80tgaFpd/P
CBY4+P1A9rf/bauuZDo6TzfR/Kqi9FOcNBJzx72ir+2sSYDrWvFu+yaTgr6L+yuq
Rs1w6XMFUJFmET+/p7lxAHCEbuc0VbCo4HVAr2ORvmKTG9rZKFPQX+1b/+ivtZnB
1eWfe1+3SmuRrZh9cBh3sqvSWF/KPFMVjvy03D1OGnNIrX+wdkMbCmh8+nQAwMpN
yq4Mc7bIKNIjC8gG6l0CAfoJgNTIfJTu2GkLLROyZO/OEfs4esxNKBfty/GhTkWj
wtdrLlIEPiRZBIef4ONcxQ==
`protect END_PROTECTED
