`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtWO9L1Ic3GoL88UTf+fTrZHEA87SlRuzVfGf0FnpNbyVznbdX7BjIWeVNVtb8Tm
kW8smjfNawrn3acxy2UgCqC3A2lNlj7jqAYJW8jLWH/aEaiQtBhbHb7CptfsnhJX
jsyWBqEKK9awVr9hbTQUys5/Dl/zUL8G8YVNJQV9lM4mZ8lQ5IU4KOfmVtSHOTrI
XKXRsiq+QswPn35IrT+NK7cwkZKWRYQXUAbq5Thrq5ujCzEFA7BIs3DWLtYj/9hB
+YdfOTFuN4UCRuXu4yAwqIliaccaoKmCXpJ7Lm+Lj8H4gqzdOZD+//2iBB0/WozD
TT0Gp3w5/rn0RlK2x4dieF1l1TtWvIOnj0IPpsWfbxw=
`protect END_PROTECTED
