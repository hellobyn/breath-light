`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8YpZejmueX5aAjNzMTFtfRT4VFlhvZnpHFSgQ/6zL7AXn9NS+/ntSsVoojLpgFD
nhxpU43wglowSvFk83zAoZ5UeMzFdd286ZcHiuJRWeCPl81qbGCbKFeUNteoImfV
PsBjIJR/T4R1Ro3GiJv2tJkGdFVxDuZp5cBuF3f70/VM4IvKIe9PAHDuDGPDt+1r
Q3XeHyOoKQI/y+bfDwGaytd2f5nF0BJIhHe97ML+hPiVmAsgpXaTze8h9Lfrtyz/
fDw8Rz4TVOMeQOoUwO7cucH7ugq1+r0C2tq5MTLJ3iqHzCVaGBd2fPltE+xCYeDT
i7w42/Oj5gleiBEscaHvSwskNoVwG6yr1znaVKiOZShe0G8b0mcoM2HRkGdPOD6N
k+bqWmzsJWOY25VFgLfh0eLyaT6BIWY0ebad9oB59NL6LtlBEpg6snkNaWlvDDe5
lVWw9KfXMtClF0G+CCcIX0SGGHwucY2nYt1JvF+IY7yOrwhEuGaZifoM+seyfEJx
HNBWCooLcXzMLqBDnjS1X86lNQAlwXJXi69+LTfICObI6ylDmHGIfM2wlp7AKN6S
4gNPtf2pAMAxwiRz7Ftj+tr4G7055uhLJkMv3v7VyLcfrfds1tyOeu9Zr6Tn+kQq
fCUqzolvf2dRdHVp3CY4MFdFxP77yF2/MAgPXDnjl2lIwJJg7HUn3YlW7pUJrE7c
gXr4ygW3490a4m06qtkWWkopudbq3iYrhdO720OcH4bN14hvphJqf5FnhaecHM7Z
W4xYjyqhE6JoaUs5TGuRiDrm3znBeYB3RELUcLqZY8kVrHuo2tj1A6fA+F+OMDml
1wZb0exdieec9B5TikqhVN++eOlrUaUYWQw1aA5DkuZNWgqg+kDSLm0hFUhpqgk/
kpMu3yjJDEUeJl+JBBWvAJbVM181ZfRmGAk4H6t82O87YLQyIP1vldU48y5i4QZG
6uIEm3lcvulMVMfjSGfW8tQB9ZeNbafQo5HzBjjn9EW/e2p9V38xMwQUc+aFJZqs
i4ll6irBhEiZEvZ+bXxOFw==
`protect END_PROTECTED
