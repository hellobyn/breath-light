`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02xtSHm4zuIJStD0fivKf0rzHLJYbf7oxAj15AVwwQmlwbDSltTCOFHGctXZtZCG
+XIz0OF0QMsSwWEP2X90XZOrTmvNd0hayOPn3iVhj5zYtqLsN07+FqASdV9hS+ey
pHW8sY/4MdrV2QKCcWC1S6aIG/Dj+paN823hBFbJ+N+JBuO83uiLOc4cNSIhqFdF
hjqEfc5UTaQXI9BPbOfSr3fMTbi3HgNToXr84LVlbkyopLWA0qP73fkOHUpVu3Xw
0LUR790vloqysiKWNQvHK5frG0IuXSxs8b23gS1C419iOGWHANQqKAGJNxTVthWy
7siKOiO1QtuL2KaIgsGzlPlm2vMat5CDIuiNUYhWQ5LtSqLz0BI6IM42ZctxV7+f
RWp0B3MowuXpGgDy+Z8ET5h0xpHdA5AxpHpC8S4jVDrDp4p/dgiEuq9X7L7NPX6b
mRhs+hzpJvWncEKKroD3und11dMYN+uY7KPjdCJ8ZaqjqL44JnYEUCOP1AH7l1pJ
gPA0/Kfe4hhvgpCPVoNPv5mOW9O9I7RVwEpcAY6DoNHJb9Tl8W12HU3fR+BHaUjF
4a+dMGAf8T6OFSQ3MHSFlpsxotxjV/kRiErnjVyoPOCqhC+ZuMoJDOp0IwrBpNBi
fhxLP/eg2JPXHVo3EKRjms3WGoo98s4fawwCDf7lgSdrASe3mizIFrmClnW3R15o
jtlcPL748Gt2IJLsYmkVrleLKkxoyhtZc4ITT/sDV8bEOQBOF6u/uG5UcZgjoZam
O/SoESvx/UuOX1091fNw+3cYDfxeAWpDIp2MqbdSns8zOR8KnaCfq9SUrkBMq4Dl
65/9EQp9UiHtwtPE59Y6E3Ow/VBZ8FU+cl7FoxudWI2LtNjVTf3SBJziOoxZqVZF
rneiTvxawKNsk2LKq082tFm1by9vHqB1WnjB+zXVRUF2cjuNfT+GXCmbaWyzY3Gx
fhonbndIEwcxEE1aOh9Dzcf+Rv5qy+3QkTYuXlNKwcy3JBVBCNtmjWvbyQlOxCz3
L3cFH2ttOI7LaUo1AYREqYbvnO9usFjUbueSxxlwWaYnCtaynwqBJdLr2eibRlOT
ZiSmK4AkTTEAkf35MqryDkwvMI01/G+vX5l1/V6fP06x2cmqG3DAQNeCBgc0xdz4
YVwzW/voMTdyGJgHHQU4dqYrpzfxNzYkMV4FjR39OLze579Dmw4mjX8csd98pc8I
Xr3ANkjG+9EBO0fIpLl8hfTcF3ACIQlcaDuROt2XEIy033h5RkA5xng0Ubm2QFwQ
hcpxH+/+SzX0HgEHoCBPJ2M7gq3gkSEO02BLNdgKxFatpqoUYbIC01fR6uS80tGE
dC1l6qid6sqr8BN8s4X2Bp/YgG1YZPaZRvzEPd4lUnjM1TWlE7sg/KgeDk+i0R0c
xdMmuZru6v+T/J+RWzUSJ4ILZaKXLDI0io4tIJAGGle2dk2thrQ2Lheh+pu2qtFc
p5PlG5A7A9g/HEAqHvjbE0DiLDMBIMuW+X5TWqxH0cz26FHRLlvmFJ33+Tj1saJj
W+JdBeXh2qIzi2R4VnZk8hwK/D8vrbcPVWjCvJ+LdJHbq7CcDl8xZ0XG3ZRfm4uA
NXFcKTnH4DVYUoWGtCGlYtqzhs2Ucr6TNjFQjvmMSy6iID5vognQwkJGWDxEMU1+
26wfycSPN5CzXZrxE3sJ5B/Qn9ri37nN+MUIodpWFJsIRA1JXiWE8fq5jw32OghR
BBvvE9kTPIplgSKfGla6Li2VS11e31RRkHTSnd2yZ05FewkNC3aqqAuwciuHP3Yp
qZS3/iw0eobI+Gdz/jbJr9RYaJgyJKvENe59rGHRZ9bYRahTWzZUhLpKiOznsaoz
f2d2m622d4sn9mGjr9G/8N3bQoKT2mMGkgPP3kJzcCxYrjNc6ZkQK4LI+8hO7CuV
ldFdG0D2uHeFVxNt8erdovSH7ngJz5cQNSxraRhyV86hfIvXYXjs2kzic88oGrvN
J1tql36yDIYXvK+jJRgvFt7//KjPdB1zPIHk7SNjDy+za0Cby8lyTniH0k9WI2Ks
KVF1qajmKmo/fq5glr2OXlZtznGH1SvRDFewqeP0vZkpbOk0dzQVZGCuTl2aFXM0
Keo817dl/uFif4pdbjw46RzbrIGfX7uNY/h7A8BS+140DzHjDQw3yccwQYePVCl4
E3fOfBWneyp/IcP6Xo23duVXZYkVD5qtsCkwP2ACnvNWhBc66K6K3WxDE/WmPXfv
gWgBkYUswteOzni5AfhSfx9WiGqcmBo0gXAZkyGWEqt1OBEaPcM2FzLFl8tgolPI
dryTeABUEm7CArSOLho90tiEZTLMG5ZR7RFhCvx8i8ehDYR1anPTG367/VLpO7mJ
PZ5qNsJh/HXWeKvaUb6lFaFDzTkcgE8D52eB299kBP5911HeGL/MU+OosjT4tgZB
g3dbTn5J/CGx2XHY3ADEJU8BA4GxKsUtt910xhQ+yf08y3YgcOuwsKt3eIf6HW7Y
3mx6pbOvH/3k1XyM4BPURsNpL2Oufa8n9ZxvDtgviuDkcECecZuO8fU0cY7Ixtkd
TDyJ9bSxMnOCCdPrB6OUK25EaYWelJa9YZ2rXc145kXrozA1GIUI3KrIIizh5JCE
OLrfAOWUs0PeVvULdB/yWc7qL1G6SxZA8rSFy1wNa8NNkIE+vAZoy34EMxrVmtYP
i7Fp0sUit6Aa/MryLpeDsSMCW6d6PAQeAOpBmpmp8xJU0wNOWXLYNCMC8pXOtoXc
pAnbW76WZQKqzqkJgtgn3BLSa3n1IqcGbfVGAlpL83bTqzJgE2D41CfqxOSVpaF2
Oue4p5Rz0NLN5O3ip+HoOy0wWWNK/R3iw541zRL69EJ9hVFt35X1dOzol1fEIx93
K6YYp/ycLxk1Z1OqBbjhnxiYksh2w+hpF1wphdFiCRkpjLvAaMKwtMw2TXFXx4hd
uSTMVXgsyPjyDAzYLuiPl6PSIXcRiyCBVZBM3s7sfixJElS7q9JVlCj3x9qp/ehU
noRfFeSNMECtRzRK/6ZQtmJqpH25wp/OUaP7KEoFYXNKOKGLKevrbq3PCA1TGKYF
jShFSCYUI5zo/weu7aCXPsTCPcYH0hAuoFTLF9QlxHQlfsrb+cRTcd5Udo0TsriD
di4RtoZk3eH5d/gssnS2bParVTxVdA/2MJFy776dsy85Vcw4ShB0pQDbSsVG5eoZ
NLXzzasCP0olVNBhtryLgWWYBf1qAmTsU6j1ISoVp/sGKbSVLcXHoI3HRy91XBQE
Y1matIonnN6AblhLTRbqxo4MZf5+ks1AzpRvOUH99hy7A8DO9JFWLckY0s9Hiq05
PXjxucHOOhaYBeJXZsyHtQC5YKYq1eJMJUo/dburEmCSmXjq84ocl3jbR6qcRKou
I0Zmep/0jFiySo8f5jqwwI/7UOpQwijnhPX3O2q13JEI8e0jIb3wgn7hhA3/9udo
eMpT/MurwAnTaASou6/VLc4Oc7PgOyg++J52z6en9yAkiTP+TgyvOIX4zQ2Y+ZWN
qp8uOtKJkY6kmT/lRfkPtUlmo34OEY0X+eOFPCP5AGeXWunPcHCpAbPjLk245RWN
9rAz6Ql8a8pM9dkaF1KZ0i8DQMw7zRv5G1KBt9DLcIEz8+FjU6awbQ9wxVeAtm/f
JvJgT/eIkXs5sSg02WDViqvUp1xrl74dd6NRdq3FGqcXCo7eS/jvsQwhjRcX4ckZ
scKcReAscaeAuKPLq2P4qiJ1uupDVSlL7l6rCv5cinZXKBC7BGCPVVbO11QxOyAj
4MtEFYuRRL+3lys86O/FfiIJKdbmUoBUdKvZ6yHIyX6c4q7xIi4ec8Wmu/Pd4gTq
fquFeh5r6D8ju1LR15wcCYAhqYe/Os7mib+rXwLyvDj/MZaTUT2CuXF8QC/YjHXp
fCn3dBjL+g88QTXE5mKNpow01FOg674rvbvW4QZQlyVW684LzFWmUvyRdKqG2S6Z
RUEchpjo/ep7Wf4J1seyhlFQqtMsNbpysJl4q8O6EAjP5En9eHNC6FqQpbqoMO3y
Qc4xJenvYGAXLxXHs2ZIW5CteweY0KdeRs9jslLr6byh8odtMnndgFM5ZfKKjcrp
axyImBKc3+Ah7BQ6y8EuAjj25eJM6wmvy8bEwp9dHSmeyfZs/SFb6g+oEsDS+2Nk
F212UNkvLdc+5eEOCozM8MC469uPxHX6CjkjfbIwjXEnkkLQd1AHgF7mp9j0gHmQ
PyDxtg3XS7O5mib9gWH/qlJu5lKh7M2Q6qSqA5mrFkDzBLfeplQr6hR11e5fJmOY
pPA969keo4z7LIvi4VnqvltB5P9qH2MiYoaZV1cHpWckfdCQqhAFmLwnVF8O2foB
2TD/jhe0SOT5/jwXBIqI4FF1ik4rJQXR0j/D24JHjf0AfjW/np7snKufsfuRA91e
cqcGQsm706llj3pdRbQvHYrERoJfB3G2xWSMssf0PvNyeNScbRC+1dbbHmqLC5Ld
5AzI2MTRH2pMalzWuOGPYxNO5Eg1H0F8mxFqhHb0LDs6WwDr9Pjj2b5PkgJwpOQn
Nxh99brLwWrAEJbImfaARygEQLmlHHKZ6RN2OxN2uolKG6C0/I5R4JFWeM0ntLF3
`protect END_PROTECTED
