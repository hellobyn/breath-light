`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MCxmiISQd8zwAo0OpOHSLhmnNblqnGHzDSj9CzTZEhDjOYggY2vg+TAEkkvVD2dd
mzgoTygKp2MR2H2RFjKLsmv9Y65Yv6n8gr+vSX16vER0gfCzrNgz6OCEq0KJN9w+
pz1x/dWSJszhO0g/woEWtgGj7sQMlfHdZIFiqgTAa7CD8izEwehN4k77gOaJk/nq
g3aYJyc9x55tsU3qFy3w0ovVMO2xcvbfNx4GoHbsTWPuO3L7YrgJKgeUaXPxaIOX
RaVt/LtXm+p7EkkBYwXlW4CRIXZ/Eb0BIjpGqaf52s81v5Or4qGMLw+IQ/x+WgoV
mjm+ro84G23EX6BmlD2jrFUI+b5xml/FmRtg2YfsKXUqj7mBeCWzPcZp1A2LW3mI
SBX5/QHj23f25dCJGinaW1N7Cs5oGZ+O9Ia7s7s64gNDRDBZ4u5w6iMlQ+p6Ve5a
AwIg6yxOos2eQVSMcGZ85o+cncbRCwDL+fGv8HQIZSqrNX2Q0QeKez4OCblKCzV7
Kn9sIXOfacR6DaxNcfbS+BcuA/weKUW2i7vKJh1qGxO1tGEVCSfUkJ63wyFniOHg
og5240164S6wsgh1QmGQncVgi8CeG92aC07AW0V8l2SRXAvzajCepVLSm0cSM7XG
98sVpf+NWigM+oYlMt7lsi6/7YwDOCVLlUDKlbOcz7qPQ8m4ODUm3lVYRPAIfzGu
IBqJZe0pmYAIhcvHQYkD+YpGpDr7XJ8CVEcqpF9/MAPeXTDRdFOOVFDeCDVBVN47
zR3EY26gS0N2ewYr/wBvcCljKGdJUlFa1R+SJJwq2+Vn2LviWZvebjMkQhy7f5+j
d1FpZR2aL0P1r4TnGEgoaM2nUbjm0sPFD7E3fP+aCYosMiFLqRz5RCu3A/COUP3t
l1+Rs1jti5v7wmGyojl89mb2hLk9DSH3d1Po/7PptMv8l1GOBCr7m18tNqtfKphF
gXXtGhPo5trHFpt/et9KO43DRfcl1+zwe7s9pfS196Smym7rpSl74NNShV+S0rmh
9yjMKC/acYZuJ6z8AkyvTAQ9+i73QlfMgFdw1zZ22Ryt1BMvpJdd/XgyK5a7ik1m
Jdhs4lq9iDQNwt4nFoRtoo40DgGScuFJ3CyzkER6ttGtSVPvzqXnZHsPSAP37g7A
wsKnDfRaAg+zAJT9LKTHv9U0YAiY0g7o7vu60stt6aaNjkoyD4zCu5x0CaSV9gng
cWWWQVAGmUvmhk7syhURG1NX8/YVBC/JLuRQ8U75BW1NwqKqGc9VfUb7yXMlEGIS
BDjmcZ/UhbBwq3o4kOcIyoX/RIe2V8/IBsNbXqNDEJGG74P7lUcv4Af44kf7yJ5K
Jvk/YOpxBRKz3ZO0O4T69TAluaG9IuGITZQktAQLLpPm4mGbSZFs4RdXoqa2FtZm
o+eXhn0BYmG1obCxguip+o7QLD/Y5jCnQyhu/K4ecPZ39Xi1wKjfuLXNX915Ua6A
AgaVjYLgQAlwOL7ylYBUfw5ey655/yuiUMyQFfvTnzk9jj2UErt40NIynO5bD+2q
5FfxbAQrVb+Awwe1+t363Flk803bcEyx1ftyYmOgu+Umufezr27HmJ0aBS1fO/e7
vqJIJCcxJepaNSNpUDCLnSUs1GypoQ8feilFBcsp4lTuWNDcrlcrn+Ys8btcxung
N7omvT5UhSOGSn1IZAlt5i8tkCNxraxEt8NAKZfqVMdVgI78c/ultUxyVrp28vq2
BrlhiNN8Y054uW2cYQi/UC92jJEUsdvSmo3HvGfATRMOs7Yt119LFfAdZQFd8ukg
G0ft8NRFpsduxNc9Jh4l8amnEmGYgxhaj7CvpD0mJPcwPJEY+5DDdq6s63BdCcW0
HP9Z+OwKVQoYQPlxmfQJ7KpgZ6JbR/MD2z/bGOhTFRLz0SP9jw3wz4u1c0AH4OVn
eXUzMz5L925MAuAQpJXp+fNUQVZUC4GVwh6wGoR9Et/BF0U9TzvOJLi5Nlhs2LHH
5CfaILp2wrEbipct0ZjCuG06hr6nmrtBEXGXssHD2tVovsLURhtSJTmL/wmbeASQ
wOkmGhO6YtqU1H/4UKEDI3f1aSM/2xZhJtX8X8ffRG1Bdvth/1XpJt6Qc7/UnOQA
PwwUwI0uwuAHOvo+HaZytYEw5J665qMQGk5g1VO9gAAmEO/qHJLIbSF9YjEoW7Nq
hbVtbeSaTFPFlvZGONuBMnN6JeduEnGGu3oGM2BKE4m9PUfbSkQt3B5B/WH0i7kF
r+5uSON3qpa0Hqoq2V9Ph6P7DtUM6R/WM4EHfY/KprA84UislAB2T7XhvTAp69kP
Ys/X5K9fD16UEa6558TRcaMMjxgKbY7KbtN/EHY85+ihg7Tc84JzP715FlR8SXch
Eb1TWUlgtmg+pz15glwFyzGzu51gatI4Rm2aqh12G3qdYkyA3yt1I+QS38gYiKF+
0Mhx5IUq3/EJi+rg9QthaFZO8dAp+MP/6TGAirAwZzl+HVgHHud3ktVvkPrEzInW
pPV+fQh92GvzR6xv6GV6JF6frMG3W+FhS0Kyj747vnQEQejnyYlbzlDkcpk6wtNF
b5e0g0kHx0k19GP1hHgj/349cQFyiZvZ1KlBKu70NW1iOPXwb/Sn/opBsL/b+WvM
uWvuTLYgSszMNadWtGxfmGsaoTl299fcoHrQGNA+FFYvT9ESgZckDpY1okHKJHUq
KhYiF6g/GdFTwcbyCUlL5aeDDWopIUa9TcJ0wFerxYdJJIKd8tLqTGv8mqZxWMtt
7a+PLbsie1JTU7wX/3G4gfW0qscQnOuKk76Ps6A3M58bOdFAbE3mD5TAXQnGqdvC
lDbil4+3LRdvxiIVmqT0+FwnefVaD3q/jjftdT6d5h/t39a8176C/SX1552tSnxh
HKhgqhiff6GZZr3XkX4QK4l+XynLs7Sh8x1jaPiJGurW5LdxMsmSNP91tBM+E7S+
qMbxYlL8aKtD8refsxpSHZDVwxkJ7fTQUERVyRCLQYQvYvM6goNCnMScRRRxD+wj
gBS4QTfNxbc3qeStinm4syP2ch2lelAvsOauWNwlbwAMpxYf9FV5qKf4+xBrWixS
a0lTEvJ0y/HAU1DTGqvOFY5x+2Q9/A7oAzXAzwmTLgPSN8o06FuWnIeWd3RBZWd9
8IGTJQ783QOluVRbKWWCPcKtK0n6dDM6mgmP0ZR2t8QS58BBe1aIegvyskQNeuF6
uEw/sK4IAt1k2nh80n5DlP3rha8ozKvWslSvNPMLDsAIOjndfRVmEahwr3fBvWVx
1MeuH312WAgBe1jYL1YZmxXrBMoofsKuTQONYCDfjrndGWq2GZF8d+PllVl4wLZh
9SpG+UVzUtDngNNKjz/uPP17m/wUDLeBGTo27Dq/q5wDCSyUvmHhjGLi5s8HUPjt
9g426nA/o2Oq2j43BtxLWGFg4k2oUMTQ38eIXKnDnc9on2Qei8IyEOQD2A5tnuzq
/uECeEDKpOwVfhxEEN+sekEOZEUP7Q2b/C4ov+hg68im52Lx4H7B9srYwxwhV3hi
LDP8h7bxvfrpKNPK9vG+9hUh129MLoFG+fA3wXHCFh8Z+YK8QFC5iQLunVvgUmL/
+5pNbN5ru7ohHvWBmDyfoGcNlghtJ1n/fK9Bd6tKpjBkdrVvliJCcwsrPSBAPBE0
1tGIiaQT1zSIcGDubzczifywJsj7AeNPzxg8ifV2wA05yAcgkEYBxdjlfEpMJ9kb
3RUwH3U9eP9NtALP47B2hfC3D5l5ItYMEgTC5NcnR2Pmu3lisRELjcmORv5C1Zvo
Tn+M2M1DlXGsFEHT4RVBQTm1042MDiuh+TdXon+FWC8Tajmlxa2yY64xsWyXSyXz
kTqZxqABFOa0howZSTC7FWMtnVtuzYm6zwBmm7Y76UrnG0FVMlo0PsEZ1YEt79t3
mpE52f/b6Wrsj01Xh3lY+j/ZpS6+nZAnWsRVikDHniwAHaXwhdPuvt7k5D6QBBkZ
7agY2s9OovQ+jpEgIcF14K766YpK//H9lfnRDd2Bq4QpfPkOcNrWlsaZH/E/39kN
GspXH/o8UAMSDsCF627ep5ntyfE/rSZ12Tzu03CNTvdDP4Td3vP8TClI4pidkV+I
WMNe9akECtCFuMXaE9PtgXq4zjP7bKX2KeN6ylYZbEFMx9Idb3l7t5Dpgcd9zXsz
E+44YShXyLUZaCsT1V55EGWSloUqQQrfZMsbvDX4gchDq2vNpTZ6e7rehStciddJ
JtAI1qw+YFl4DcS7X86MDCJfcgOVQg58ObOnGVY4UzZXosXsHNAOKm/Re7lRpSb/
pB8IO+RZqZKJ7IgQZMvX/ITZ29iWlUccPv4cvCOHW71ZSOmmsu9PqI6kbQjO+1cY
H61KoAIrGGqVugFXJKg+KOBsSrFwqi4qMHVV3OZTIMr7cTsVNwUV+Wt7xlE+cYHi
BfYiUI4re0vTdwZFijiu2KUZzbS7jhaqVqTLOpWzSIJiuez594QuBvZPCAMZ/xdY
cVThVCOtXRhA238ZieBh1mQ4pcfRm5l32qOsai6rOCqNXEWRvIX9zMdmtjt4e1v/
zQiIYAG+hEf9SJamBYK2m1OrRg+AOov26H4Zj3J3v0D4LjXb8eBF9z7NYSqgbx4I
vrI5aXctfdD3an0eJws18PqEXysbdlxQlGf1tiL0Np+ZpjwhYavxO/h71V0wK7qv
X2oeHVfG8I7LFj6jup/LfOQmTg0TiqWONZ1r0Ad6JL2gHp/aRnlAyNugbwosm4O0
aw/nqnVEUh+Y9/ShXyhHgR5jy8s0UXjr4r1wSD40dFsxc6YsKiA2kbi9v7N4U4i3
INUVzq6OhPFEx+OyFn4t5EfLqyLBh/Cyi/UstH/7UZA5ATsxr3zxDs4A1HetBr2R
9I4idcCFP2QsnKStqSwF5eNRkXqjfW0XQQCfjv6mBnSN4m0a1k+S8i6dieTB7WHP
Vfm7iuR7BPju059uFO2BjNOeSDmEc2P7jyXLtt915Vab2QOikYDcVDMo/iMfp/I+
+9FoOdBf0wJJnqgaJTBoRvd1ptWP9kIM089Ctj4u7MVR+v9rT0B9UfKMpFAZ1xCe
k3M8etgL0XMVBj8O12HFww==
`protect END_PROTECTED
