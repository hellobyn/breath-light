`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R391yUzk7eJ1MhLurIbWmHOii6T0Lu0iZrOFovbjEDL2zEal337vW6c2kK32qnkm
9VsJ3Z8wW7wBT5T8d9Sn/t4gApJj1Pcd6P3i06ireSbAIGys3O+O/79bnfN24cev
0ozO8ykWd1NLYMb4Cvugaeo7J75F+3md4lZ7Z8DP4kFAJecxqmK3BIsAURNbkNdt
qyWDFcVKRIzCUpnJSo7BFQh5SaFp5e9xWVmJxf7+CCIOu18banM+jqQzHUow5K5W
PjfWxSp3NIXA/g2D1Rfyv7gW5yq8Dh84G9y3wDaOXTEy/Rf8DYXCUKxtr7jSG2cV
oVGn6u/Xccfz8NlBeLOfhxzIQO8sYiH+KSCSbuZiu7oo8h8JK6llbPOxOgD19nfv
wlZhxeoZzuRYvYRTl5cHjD6FBDYo8KUWL5kVGasqQPn/2acKqKSWn1mWTH7m0r5X
zSYRvgLsy3EML02MSSVXlLutQLjpfEpJ7Jm1KzAZXFq0AO4tCKH06gcUFjj9EwAo
PPCvY85AzSNSuQ8+cX+dri3fsAWDB/PvDXY250kZKp5xnvwww29sFRhFktM0/lL5
Q/kgOJRUzdfx0SkKK5zBohVL7U9S728vVFxQhVOkFI0/U6pm+sKCPtzIV9n9oV36
5Rhfjcon4e2kROJ1xRphuQJf0uSKjbYijCVDBJAPl8qeESJzWvnSOE29Z0RTA3Wp
yKTCE9u/YIrAga02vF0WmUMttr/bVmGvxZaDuhNLBI8Nt6AJ9rPOrDGJmRmV7j5J
atarvJ6KaVvEnX4SzTz8ayvKXCg7jY9N0wj+RhIwZvFgHz8Ssy8DBodBXZnaGP4P
`protect END_PROTECTED
