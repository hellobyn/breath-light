`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2bb9U6uPBXPOKo7UR0wfikfqqrRQh2xwA0F9AXGW24CEk3cI1wjVRoFRESFQN6/
Q1PoJoi0GhUMKWE3AJXDSp1Ej0yZFo9k2Ud3SfCfWKtkA0fqGvSAA9lJsc7lf3D6
uS1vg+RXn1tqZBnPRFN66JagXpe+ocoyyfLZIzIDZphtiycnd2QIARipjyNqlIoK
TFaJ2TtJb8ZFqpRFnCKWwbijOysVpuINAIbe2xlhkSEvWRwFDTNXheOVk1EryOKH
53yfrpDydZz+PuHr+IkmxsZzgaOylA4SaEU+RypRJy1F+RAUBFtLQEhV9CGbg2n7
nLInu7B2pMrJaDC8//unfyx0JyAJ7Hw+85MXDxYDMFHdy5k/15PBegay8+KwXkhA
D2J0tDZKJD+zhNXTzNYXNGhiUhL/xZ/ibeIJYsJFVXNmbGQNLDgwDtHVY38kcSvb
wzkqil7JO8TPSzu6z2ita7ZjeCpSKy+rWAtWoP9rkREyF7PU1osQ5dt4krL62MHl
kLElJsxYEPPeGWoAyEvY7qqCUIorm07RuXt/dYufQqVRsESE3JVUn0lRYyKzPYI5
yQPY88w46YPeITUVYMWomNY+bT0m8MnAOSHxi9kbINTOb0Mb/YNY/ten+IlKbaJK
hk92b66IbMxJCKI2Csoi03tnf9DLVt+9wZsOZd0mf2seatJqqFQZG/W6CRMoqo1R
bnPm+uRmwFgdZkvOPY3R3UldYLz/H/gwVHzhJGTUlLfSTAT/aRuWK1KTG7xBDO/M
rqTuN7GVR28+gwN+91GOEZJQlglUgbQIdIt1uiw3Dv4oorFNEr+1+XHvWDajSyih
fUPJTfXydsGcoZ+FiwxSDfUP7MBEN4yWROE0GS946Vw5WQoxWFX4Ksn/5FO0ikRp
jkyh0wUFTtlIRc0S+ftReSlNpJLgoa4J4M4KZPI/+e+xZ6XqThr4BcZGb7/9nqRn
6s0uyeRJ7zA03IGX4n/9Vl0hSyRSXa20zigtBT/+F+jHwDizydPZY2ycBEkcD9ay
LvS/J8sTe9qMdFzxDa7KQGabdHKr4yK7Ono7f4TQJ6I9OGnr7ztMa5ri5V34QPOU
QGurWezliPhTucTJ9jerfko2EhwYpuk9W5QHCXPRP6nzhAYZdtJpTbFiwiVhUQp/
mOrD1z4kpiVdCzvKFxmnscOIgmHfrE3ggXd+jqxtZ/3pr9VxwHGaKI9aDa/g1PDD
ZJ4Wi4M3NVzu38QVYbEWu008xDV4x7Y2yu93L0wRz9NChOqr8dC1o1KgKKv98Kdj
dwdmoowbFhLQALkwQtGYBh6w9ziFEnm5TbRs1h4hUfU3EX3jYmhsC17noQ+v3uWT
QNylVgRTGsmpwWUklPa4tqBEVwPv8WMCiIWhy8XiqPun37W8dHDLAqttzuZIn/sR
5UYT4G7h9t4blKgENjtFx2krb2Fybc8TQacI6pXeO7d7IzNFkrm6ykK2ZpOwqmCW
5sjdA7TvBlYdCwagS2zeBt2/Fykphk4vrQzl76fqjiueo4nSQZWJygMrOyQF9Sp7
aSmKEmx1urcKrqd0IysfaA==
`protect END_PROTECTED
