`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICm1LeXWYb5fiIT7XJp00SxBLH9f/uRs5EdnEBRbgluZ5ehiI7AfE4Yu5rXNOfbw
eiJGlSZp+Vy+5XwWmAh+WHkMayOp/54Xa2QmM1kZz696I7W153RvH5okWVovoyQx
ZZWp9UVCp/OuAigw9kGX06kH55K0KbP6DfeqYq8i7cdaj37GASj9wbo3cb7sa4ZY
Ks+GQc1qQevEAep++fkjWHAvjyopv4BfJ6AnjNdgFUMIeeH2qCwDtbqYPHGwXkol
H089VoKPbL3Mov4aCQTtb17F34pUhlifT5B+551/ejymoeDEIMxV7h7tv/zsqBNQ
+e1IIwFVOvthee/Gh0aL/I5ZpUu831QDWfQ0fERpdkHwAqIt2KbtQWahimtjnGIJ
JMNAyrLfLtXauLMtR3CidCWEcsBs60kFAARKPFSvY98yYerg7uzlFMUUtdSgwuVz
XlMDU1jQxYaBJB5bmxdqim1CFKHVAe7RA8L/JwQF6I9prvH9UR3xVeh8NLZDgtt8
S7bp8AJwkzkAo1b+bLmrDTrfue/W7q+EnENnJ8s21eOoAhsehnoJY8ZRGV/Sg2J9
dbX77utl8H/kZosV9YhbklUiHniMfNWptjNSkJgIOLor1cYVmWAW65ZdH+btlkji
FrqlTvtZzGIAR+0YHHvCfJvxmY3UoyOJSnFlNELSshSYD5tArJEOvJvYEexiGF0G
g7txAAs1xAYL7/YdTNGMOtvZiVLf9/JoSemFwBeIUrO5NNjGNfyEfwxDbvLyCxYm
UxsacZGByAQs36sxLRoCL3Oo/hxHh0BNH4IiohhqwrUP7plOcajfJYNw9n/liPXS
YX4awec+R+OHoncXwJpvzOK7HCtwwQ2RTC2yRcZ36E45+eU0KTwDgitHQjaJ0jNp
18UtFNvE3A0r3FRrxx7tVqF3jyXdq5fN6JDZcqJZ/d/2LrxtvtOaFMzMPxeGajx1
NvThJM8OhXi97jvY02LcB/cKsydZYQRS1jZrfTJQ6tdFa4TCuAcy0MnlWjyJbVss
WZpM/p2FZFPUYlyU811gAG2dkDRimb72pZG5cfBXvfE4bkE3zEE9NBJ7UbJIYPZm
VTsk6Cs+8/jB3L4W50xrfXRBDwTiWQUq3GvCAdNNsYZf34iG3cuUgUlH6zklhUUP
W6wbmzTVAMyb7aE6t/HhtYB+n7H6oU7xtV+OLKFVQAs=
`protect END_PROTECTED
