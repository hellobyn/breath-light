`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZC4+kGIUoI4tw7nWTI6D/FgQxAYaGmYO0V6hdZB4GJiEnrHYiKwO3zcPuA3jaU3
Rerlhbh09aDA4+eQUlufpA0i5NB30sXF7hduI7jadPWTumTgiHb99rd/Q2RbvqLH
l4LMbG4qh2mUgQ+jYV6Q2iYM9Pd6+3An8mNO7Db10/rhea8VYbRRi9OCoOzrutA6
0bhsdOtw8VjXS/6d2aUeJIztPk1EN6B4nIhhCkAlGZQzmSB4qtwzQ+qZx5MylOdC
8eq1Z0Lq1K/4U3vEqxu7BzL+ET3RtRCwZVjs1ug0P0s+HT1/dU9LPAiulwVczaAn
bK5WEhjz1w5u7/BW0X3uiSC+0p/es76rsRm3d92eiSeH0I5VxAGEe9gD4zYVaNQD
crTCtpB931HxYNUZOt2FKNPlccROOEd73Xn9HXnfEOzGWnkk9tCoQ12rWSVmvehz
zcSGi2rKuUc4gH7JTIV1BHXbkq40vYnKkubFNtEx2Sh0KYooYcUsLLflyTlMeHCX
6p4prVl/GVL6nhQSkNSkGLLa0Y85kf1iF1OcKMNXT18bvoYlyIfDYDuZmslnHUDi
P2Asxz9bC5L9crom0UAIKtLpvbCwkiDDDGy3ESlzVR13YgVnBnPzTw9NuAGQt0t6
qq8TDpyriHNmKsO/PQGxjTN4X92Nhlt7aJlyinEmxBHeMYrMk680qmPaXZVLtpYm
B7p8triBtb1Jh0YyVzwfY60MxU0SCIjUTR7+tgG2YoH2DA+itPxdMKhH7nH2xTkv
5ta0L41IZMjYJYVy6ffvmahcYc2VP1+l4b8lihNrHbPA5T+KQMlXa6NMXTm36XUP
W5lgbYlIZLFYc/zgTwIn/RVK2Z1PWeFoqhgz0WTFZwURghp9irfP43WFL+OYMDm7
rwh3HoaP0NTS4wx+zQv8opBWr7yypSjnz1cV9z06bpnX9mjZLHP+Ao3WNG+nVDnk
41pjEwiRyw6YcbhK1Dwv/woTIFRELKFd4T7wSJ2JcB429wIuIdJYL+4U+nYhMxG2
NENqCanMDSRnSOljYVEjZijeTP7tVad4TBUkZnsb7x71NrDxTKe2Ni5AQ95xZCVj
+5qJLtyZrO8jjakp4f6mqMtIKF79VkyEfnbn39lBMGyP6BEC6QojRVluZ1rlNcov
DWEcFXT6zUmx88GNIi4Y7AeLXJlVarelRXromModUMJDnnH5jbrZKpcrtlztUeau
miLBM+rulfw5hx45yBEVePVXSSWP51+F1dT57Uyb9Y0=
`protect END_PROTECTED
