`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqHkr9rrSp3cHJUtcd8zlm8zyNum5JTzGfcCLRFHpDNrYxSjSJmdClgFaoiQtoUE
39Q3UnqpnQdDt6qyUMIRZ5lnryEJArAoFWzX0+0QWil5X9dk67pbipB2nwctV607
oKJnoAWLBg9kWcY4vHfKpNBLrRTzX59cZracrfairjNqdriFS/COHY+2Dz9NeBcS
KNq8nfR+UawaVG5A0IdyDZAR0ewl3K8QctUmKlCiwgbb/Dn8bXpKxUfyxQZIJAMA
q+Cbs618p5Ou76oUBdwURiGXa9BisE5bPuIIZWbbziAY96Siukoz7ejM3+Zex1n7
QmIrMb9eF2jdRGQJnbAYvUgNvo7JLeC+fZ5Li0EUCyW+ovJk2bj5RfKQLlnLok0e
`protect END_PROTECTED
