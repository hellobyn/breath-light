`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Qm7q+8wag6Yh7QrYGkxN/TkEH30l+XwXFsHnizQ3mCqCZdP7fYebzKH/qyIXIww
LDxG/YdPeWD/05zE+YhjdH9lFPgOMqfd/ePSQEG60RTSH+1ukFzXkbTCREQ9Bi/h
siZ6ksPQ8fhRxKx6Lsry7nLwIiQYCj8/4nPCcxGyLrhhy6dC+X6C0tdGi2+/9y3r
fw79hFFyQObG0H0FRB7nLUyW6MjdO480hTLL+P62yton57nJXDZyNGAhr7nBGhve
0zke3JNhjpF5kqirGZj9Ggxh2PFYA23g+OzyekRTZpn5THir2zZTCx9YONttnuTt
q0NFOtMLtegNY764Y+Eim6NO2vD2iD0XypyweWwqBWw1m7IXUbP48WYadEFBuPxx
OwngKABbSYvecYAbs+Xgdtsju+0rcnKFQC14ARhxo9cMKQhNljjL9wwwKpck7Ym6
hY2W/2sVFQ/qevBIu33iH9LIXmEYAygKHsf/y8gL7qlNnZ/AjEWB80VRjtiGQYui
dHqTDnzblpM9HGCDiOpSpas5wc8uRfvrPEWlv5eUVdrn58/MSDcYcxJ5bb1nQuZS
H38e11Tzx7t4titfzsuAS+uPgGokNZSkyh7p5Culhjgsh7FcsZPCYOAxlDmRlfU+
Jwda4y/ZztQc320IJu1y+CGoFPvyHjTRNi/oxfSF+rGZiEsOlaGKkJruRYzRmqVg
jcBBI8qeDrM7oDr7c6zwSG1cQgowRP6l2N/BL2dYlKaq0bSFTJqcpL46k+PpHM2i
/ppJk521bdEeKOiXxaKmKFXoyO6siBf8EILhJHwCZfZRk93tsFZ5GM3m8Hnr6kIR
k+7V0cRc96MkJajI2NZWtf6/XgoHvFZb+VFf1GxBa+Q1Gsb3qZiQn11aqwNFsLRt
vm8d6DQ8Sys4p4OxWZIQaEyX4xSmgbWVpOBkM7xzi7nXNeIuVCSbhwwgFckwABdZ
ByGqwoX/hpSy/SOkxgO4UQAioH1tHAiR4sVGmcJfOT20C+wGHFK943JnTre7z0VV
pHYA9U8ueaUYFj7TqfGYryZyULEJT6qayCFUg9ctcIkW6ovRdKpIx/xLTXYcSiDW
i4jOlPtJiyE4JnaHHjy36E2kwwbR0a3UZuKlNpWzbkWbvYYkRxzfMhcEqzYeHYvd
Bkp/necgP1j1zAzaF7n1ptfsxQE8anpA7R/6zk4kq5OCnnMz/zHQdfDJAFGXwMP6
jVi6gfn6Q50V/HR/PTYSQyCmCijCl9kyy2en3ik1+FfSudL1elP1RKj8R9GSx2hV
oiQUGWSmkqNwEMl4TQtof8ZHxxqFCy1/Y9dgzQdl8TahumsPqsMq+Kjv5kwmDxJM
ojPDKl1y/Lm76tsaSxbotSyR7mAwrcn6OErHdvmY2rj6ttEhBCfQwXnOQjj1QH6j
FD5sQwIcK3odvQO/vO0Y6N2a6Mkxj16tO5zkp/P/TxDsaNUUyrVen01zD2ti+kjB
cCn2EZqacXP2Fy2cSdsgaAtM9us3cBE8zNc1EstDp6knNElaGNHmbcSPKu5XitK5
XPObb9Qyp553CZ1CVcBYmnRllhu2V5f6kO5QMTOvf8nrp7aSGEc3BXBR2re3g8di
2DO+q3QEJ8f/6qjTWZVUV3yP7BajuLGLXW3icWp9kf4yrFS815oXndCcz4ewMhVr
0vIRBm6PovsAd2opAcpYFFmmmhgERTIyvpJdc8kvpf3m4C9lWwP3V4eKC5pbYBtJ
5FO6kycHlDhkPHFpzwj3lByqTsn1C3Co00/vpJMAkQvQPLNM1ELTNn2A6uTDHSWL
jTUhAChtV8WeNqnvBpChi1B+IBYLFXJVFs53viSSzbyOdSWYGfK5rgLKVfRmWKJV
cdIGpgW094LvGzLAtEPQLKxqbpCKotoJzrivI98+/4guUUkRaX9jlbEp4iiRz9CB
giXuReVRJixViXBcqt3yeDJJqc3nehGn4R3L4CSBNl/fEU4Z2TTjmOpRpErpFzy+
lO9W1sdAVqWVQung7zvp2s5HhRYSfIMHfaHHfMNp9/BTPdvOdeSHY806u2D1TBPK
9pd1iDRtoGXKjr5gAqu106WkA/nlaoicmseAuPeUfJ+VHFBnElY/nQvhnDhyrDkq
ulj8k0uEoyTnCFTwNcigFlfPcyyBOoLekoVIoTYRc2GkjwXO1btYuzO4IQ8VG9wp
dcwi8Lqu3QfbaYpU3uK3eEF0IuqArUbfhMaucmeGWW+VJhN292236Og14tcGibY2
sj523Fwu+nnseKjjHQrIo0jAAR4JAf+3WN/uXb/VYzhlIQ9CDP5qzMIObKQC0qpB
GvoQAujszXd5EfW/NXLPvFHh7NgdigztIvZopWNS93tpiW9R95sct+Q7zRHYmwDr
v9ndbIqhUWh+hqtYCFhEFUkbZQoKsBKpHC53Tt2fzXSW+MZPyGq5R6fnbfw6v6rw
0uPI8kdcGqlKPgtK5oXvgIPtYsxAwIMxXH9rTSYxwJyu4EgOorpNtT28IbzG1eGC
MhS+1iA3Ooq0Op4PtL5jGBZ2lKVUBqltRbALjrFNfPlpNYY2DU2c/iNoTVf6uQgj
ngAAfuK8ietWlzCyt7HHrZx9+bmE3TGSn+7odlQXTLKdW/Nihx287/5wi2o0LelS
rxs51sATs3qkjtUew2knr0L/dD7abCgVwka8wfjlK2Onusb65xG+WdHewoUZunWn
U6lFMioe2Zn2oi8YitY9WK48Jx3ASpdvBtC994pISGflDM3NkssoBVUZX0hWT7GE
yYKTMxOJEZ8AYz1+J3scSCGCoCEgiTX8frvjmtkqrhsvoonNuuRbiTgfrvDjJnfb
8CEQJusoT4jHGkZi6yGg4oVa2b+5e4kl3wGqh0MZTb7cIOeZCsX9J4t3K376n0+/
9NdLsjGu/x+2jXBthhvXGitNcvptk5oQ7ptFlH/vzHJ++dcCDolpWB+aZ1qV6MNT
LYkBXSN81wi6R0UZox6WURzjHBeOfHVgXGqpmvSkndAJa4Z8kV8/aH1T119x9v3Y
HW4lH7TD24h7TNTckX7TMenilAYT3sGC4Co/A//lfpTm6ToVvD4jX4cdFgpD8iyZ
iyBAmbS9Fxls2QXEBinfTcMPuDhRqeTrjgYQEafutaVoCTrseWe0ypLlTp18NIbm
NXqjxHBj6J2CSMpr7UJvU7yLtpzfhQTBciwMyX5cFDAPQtGsJAqOtP5O1Gso/Hwc
3MeM/ti2pLMVdRY2gyBQAus7ZGQqTSE7/dp1O+FA++JG1VbjJY99NjVvdP2dP5xG
4E16DdCXbxKF9JxPAU9D/V5cHUe/482KaA5m+M2y0tpuBWTfjOD9Mvy07+nSAnav
WFRYnB74BKoGzsMl0+Dl9mGEt9K42vWwlFC+9zzcyat8YlVqmG17lh08UDVruCJq
es1StBapULB4ZtRbqwHvTn5i0JlGpjDUJPUa9oUK2fDTQW0ZzTXepmrpGhYW/ILn
QdNlIBkIyrkXieGcjShDNQ3Km/Uwjdn/KdKkFoMWJ+qDES6qwG9q5io8eqG7I5+Z
EO+2Lr5d74+rj6G1qttZZ4hohqLL284wjFL4Py/r88Af2X1hXGH+tbRhL3F9GnwC
ZTeN2WpQQjQuXEP4t6G+wj5zHJVEFTMI7MT1iYFNvOANCKpGiHMh5WPewGN2RepC
U7cOI1uUF7kvLWuWxHaCLQn+1tGDHdkDVy2O/GTC/hy6fr/hbgAYRg6ew87yfvHg
tKKFChHDKx1Khf+KioqLCaNw++Bgsoll0MmUFuN1Q+m5sCI/N3Q3HBt0pvVNG4EM
dkTDzBYcVxe2ANwFNPdgMClIoQaGnu8Q+xhCfMumI/jQHQFtHaqnyDlhRwAzsnB/
X1CeK+xdCXJZs+TNkK5WrBDRUdZzpOmvFRwzfVg4auExM1RV5OZ3NaHJj4Ke1XCN
LZzx9T+hlL+HF4YFncbH/pFOigB1uXG6up5Sy6wa7B6rSa6km0IzICl0/wRnWtN1
KpWSSayXBVio3u8r/GtpAaY96FdywQS7YnUCd+JwJHlRp8OTqt5/md7hw+ASJEIt
tqm7Ga2q+0lQ2DbyeEU0mJLX8oF0I05a0yfjsGtLyBdao7CPsOY+Q0NmO3FbQgvl
V3ow4vGs0mwwWNdqRD8+WEsoZ4cyO3+3FFBOSdQF8jdxSx4FK7pyAmn06xvgCQV9
`protect END_PROTECTED
