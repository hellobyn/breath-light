`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrTvOcptNtVUuQsyMsdtC2D9zx2FOW+c49FWMfY0hLN6MPRPt6ZaDoo5fzek6QjX
T2RsT4cbFxHJPINPWf97sdE9Iz+zJ3oDSNVIjAkvjlhFEt2HIrNIONJv3KVT6uDe
6bFiOo81l6+htoBp/0b85u+OSE5j5tNTqDEvxQc5JK/LL5c0dEW8Vf6DovY8pE+p
cDCYcsc6hvomGq6pmP85wsm5E8sJ4XFrpuLkorowIxbeYwKaY84fZl7Irl/4E7e2
8DJJR8W4g8WmE4s10JQ82q4ifXekHTuS+1otA5ymw8m0Y/YVfvOz4C5Aee5qjVBS
v2+MXus5hBnh3kKeGVdAjPrqqvo8hycxofUmKZ50t17/BVdoP8kyrjVkDMLCPpvN
t8E+NAix9H7tEAP6IpPGnPe0SI9vmuDBmKv7ZAbPAxPcnKBB5ubyY8WdD7VmKlz4
3hfdlA+N9acG43SFu0iOsAoBcs86SaoUUhif8aSMUv7AMyLIwIlaflDcGhgU0KyD
oqX3wxwvpxETEJwjPDWXgp7I3rzEt+uDD6UXNpb3c61u6xCozp6Y0DXYevfN7SLl
ylNQDdLvKM8yyermpY5fP9I1wnKnKJZf5hHO1M50DNb/2cOvqPC7lat88FIllc8a
0C/uB8VoEfdWgS/UXTXNSOzo3JKVmZoP7omXAn+cbzQWesQq03MQ6y0XKmikiKYB
qk/DqBZ8n2EtOUWtz9w8Y0clt9kKYxugyfwuO/Sq2+rde3Mm/HHrCP/4ybTPjy23
2Kqx4M0b2GbEaXAnSlXoOQYIev4LT+coAhGRSYoYRhQFgGdQgwB8T4zuIdOyQIs4
mZ4KopcRmcLdepbW2jAS8g==
`protect END_PROTECTED
