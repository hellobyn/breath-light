`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBypteNI3rEDBaFz1HfdYn79w5/OHIddCfZHj9RLDFkMxwy8CWDx5P1PiuImVH2w
LdB4lhTEe/Qe9UZROm7KWReIYvbbKZ+7ubIAbGNK3Kmhzi7/hL5KxjdAfVrLOYnR
TPFVRRWyFDa+EBArRcgJ2V+yTjjZdwL/rDc+UKjUMYbKPXRUSe2spwDgt9br/xJ+
Ct3rEdvQFyExL9GO058bdYySakhFGh/MvjAsQTYadp960NZN6ol8fTxpQL1BVCXe
RhwgTmaMhXMKPcLqbcNS3QGZuNGDzsfxutTx/jfcbunJQUPXjrPeaa9AtAKhhTFC
nW0msjiL/O95WmEu1suqjTf31leu9t1ff4r48OAZd9BfAvjDG87MiuqNfagbyirJ
b/RZiW9TVlAyPpp1Wzke1dVJ/amxT9u7w5grU0n5I5KCTj3bo/vmI1HHtegMTqNR
byEQXVWZCBrTOAyH5ji9CY3sx0cXN8Gy2D1VddVgkOGl64WpAbn0H2B6PoUyj1wM
t05hF07DHdZW85D6e1geRef8wAAUhQiYwMkRmnjtoNZMQnBsgpFz8zEI4z/4Bf+q
skzBWAQ8WmZ3sLwvO6qxQy42HTNRr1z564Sx/rpqBUBAwScFm+mCJzZfoT1eaNZU
sP2alcQfJehVzLRxIjbUb+c9pUwdDrG3B6GLfOkRCdFQaRP6/414caTfoLYKW1z5
2w3hpx1wBUDUbBsodGAEWAb4Ey3gQkarCPADRuC08n/I12b4ba93Nbpz8p8DQ468
i3+N6JT7UsyvCjTZK9nbyLvA3XIYkFFEAR2/kPC865uwJOx7h+IeyscBZVhsIRsM
QvBc6/hGip2o0fnL2Ecvg+COsS2jgAzX6+hyRTA/gbycIqYEAe/vH5i+Nc3VZMk1
1c5jf11c+LPVDCD+9sabgO+hK6H92tOBSW+nq7+vDqzk9ImrW3W5fqHXwP3FeSPX
qWrpBH2h08nR+ESgbladU6A7Yfs/iZ9ZyaPEw1G9EBR3w93lnyrpp/VHNkIgMgeR
JfLdQJiXr6IWOsAd84nNshZFFtXbOEKpfiGQ3ro9ftP9JGGtrpyBuVyiQrsj/3bR
zce7t3leguvKwbeSSGI52arHbJELoMEw9+q+WxgEb+kaVObEG9zBcifEF4lZ8/KM
d9BZnkOg+tVv6m5mB4W0DAX7uVuS/iDPyUycX64hhISQoyxx2jPocBBLyd4tHzYO
ZXiD56gORCPZ/F2KPJMl2JOkrv/xoRFB4yOJSjNycINNyNnZ/RMz+A2QhS5XIgbv
CjRSXEzFoIZC+eWnmaP8DhQjFpLeIZm5ubE20Aayr0bsdMDNHI5f+YLa/wsBQFZt
tCIS6NDjIuB6JBD46vUOLnAlq4NqpgdGw/I8BarNo1RwMUSSN9QFAjUHUggtBQDK
9WL2X17q0ksavu2HKmbQY9B0/QMZaD+L/E/WCo40xjY6adakFE3sO7Jpwx9te4kd
1dbSq2ajjN3qZh+StZM4OWjUP9A+UWjijZQH9hzzQP5ZTIptD6/KQasphnblCvan
o2Gcp+vJMwU8NltLW1UTFzHA2M6+MjhXxzOUSh5EHaBHhzATiolwFumoYzOiqehQ
ss1BIQyvAnwXR0+VT5/Lh00F1L+mTH4eGUemWuL0atVTYXQo3qqKEm6YAPOIvn1g
a2MC/Z/GfZs/5kalhn5y8cik9IDkkKA4uTXOIUR/6JgNdz3suVLFV6gcqyEfk2zJ
ow8RMtkMSOm4vLyZWPtjvdLHcRb6mXJWZxSyJ5JxlJyH1TNcEE/H4VM5ZQcdlZaK
OqCk8fFlRpMJOxSC6GsaKnUnPa7S+NSVtvV40gSU0gMeydS3oBodyKbXyCpjczqn
Nh4sTAWXFUJrii1BA54VO/NWSWFn+ENQZE3HsJPCMzwjoDjpPR7Yny36itRZNeKP
HnZ3+1qy0XBsOjfh5ZZ0Q0CxahrZ8ealylZQTPNpZA9ZKlS4zU9VikwtkE10RZyo
m3umMJPKuke2CRdZsLrorUci6N26eETccIgu7kvV1u8qNKiTI24opxC8wYGmZWYD
E/Jov1yXHzHdyUmWUVFeGjTqQvLuqc68xAjklQpTkQf4HJWh2JdNLUB1djiPpm4i
uFbvAeJjhOmTuqPN9PdXBQi8AYxYsY5iUJELz1BKda0KvNX5VqwPmV9EH0AqnRy8
9CeKhnxxr8HTUiupJceCWimlxQsW/6vEM7ernhYaFbDtrWRDDd3R/n1gxrGtRUi+
ZChujj+M3dFAxdwo0WD5M4Kp73wWx6+jrknyuloD0aJjWbXfc2NYySOY8NGREFO7
4dceGPZXqyoODJ9GQU0syL1ysWl91Xsl9PWgL8+StucWwtfi5VyaK+lr2lhy55MA
ossk+DWNSi8iE10+9wM81RZ0CjJI8JQpQeM8sDdVD1a7roI8HANGVmy1LHkGfI8V
Et8bvrvO8YS8GvT1BjU0uCy3LOFlsYFhTOSG5/37F89JFiL9+/PrMPH+Hl454Owr
urYRf1izA9xBSNrPBV78NL8J5G6+3n09Nas+or0ORJCCYm4TmvDtibTN7jGfAWSc
CDWhp+1JDuMajvquKjxf73fV9U9M1nyhPiE3O/PkNvQBLN4Z2ieF0BfIFnb0ZD7/
yDlU5QuQplo71IEdcX1tmEfeCu3PMqZW0x5h6Yph8z8PvF2jeXQ78heLobHdXtbn
ElGhem9YCKT5y3vmW7mROBcEpp3RRJ+iUJEb2wPWDZGsxtwHWAZzsJBiu4473XxR
XzpHTSyPaaKGEAsiFrdMZuIFtnAl/dWuNjTU5f0EGaU8CVIHHyiMPjKFVqFmF50r
UFFpLKVBTM5wc2WTQlUUUjkdigAECbMfwD3Snfh4KY2TbRwCuwdweVkDgZc6iufU
n42io1n2PHE8M/W4dnQaxZOIv5t7sjDQYgdzr4KynsWggjSgyX0Hp5I38U+VobQN
fFCOXEBKCw3CU8SOVh17QejEbYO6PEMQyb5mXxVxXwU+jlXkekZvTl+fEm2Vb09H
MvwMy9yfvWZOw6U+vuyWf1ZgpiXFVSimbdr32mSst431zgU9PHWTJM0+Dq1oiMpz
TpYc/LVyZ/k1B6j3ZFzQNtKAqd5ndnLmkEh0fXvwH8txsd09k6FU1FXF3bQrUFBk
A+KDiybATcxtsYQfJzsKb/tyHuyw4xTYQciYZdHNc9yY0mxy8/OBLpAqzUNJpl3/
50mOxUvobDzW8IfocXIfRi8zfOd3aRL5nNT1BvR846t3b9ukug9c6zY1Py1ClWCc
h3eTdcOD7Vd0GEz5H78rlPd5OAnuqWiw008j2D8CTNlrnDbxcCoXQKYwoCw4vEuH
mUeWNOFSk54beQxvfwSYDra6RPooc+Tmk8wa0VKK3V2Lr4FlERCfJdiT5VGJh1cO
dlkexpHKnazDDiXlQAd0Dbs26xvvBXu43RvyuZ+ahJvmOxra82EhP1A0+1CxsczA
244SY/xAg7CzuDeBq/C2hNjWpRCX2EiZ9cJFB00OL0fwWiUxW9fIBmGRZkz0zCZq
xKCSI5lTTFdNfVpOQvkgrZ/6uNyjSmpOH6H511BfoafdHGz8vqwveZFW1dZbBuei
5nzIa/m3hw7MEF3ci0xgCrOm3jogIB1emiy6nfWkQPnb+KU8seIS8tTC0r0rLoBa
tD3b7rR8Vc9XZTRF5BAiL1XRARKqjBNvAuO7J7LQsDUhEuVwrK+kLxqu+7RSl5+n
H3kyP1G98Dzs/P5YIGKl0dU1Jus734YL88knRtM5GJeqUQ3zUTN4ruc5872Cy6H5
SwjSBYEPuFEGH6iF0sjQ8zKJ4xJ5aTWLTlJR3EYWwbgXKbUplC91sTzk1itgNdaJ
+/0yrSqv/X6U3mRr2X/08MUCiRUkm8FBKJ4EEVeouBDCJnzAKN+taczAqWM7cc6/
LYzsN+4UerKK/Frr7w8E6UZQxZvfYHWk2FznnLBizMBrvtdRQMEvKGHC9RtE/jKq
yYNRn+56+rdY2CD5xetjGQiBf/JaRHqVsgma93U0gU5eu0KqFaS0QoRp/ZR8gDsX
bCHzHbTzsf/XR/q4uKjt5kSl3cKlzGtdf0lMXbI9V+MlDFRXNY8QA4pAVTUnj5Nf
f55ocB3irvgoY5uHtjiYMbLcsM6BUMbD974ZJ+NpBNXgLZoL6ID31Sr10Ass1Imm
TYJTAI/JgSmDqIHq/V5/F8xcEqh9vOlSw7e1ly6cuZ2Wtpm2aXcraz5+Kc8xTf5S
YSy+RNE5piTxDEHVy/QcSUWKCxrpGGZa8fJkzWuamk7lVa6lC2CrpaHgWid8IZKN
nKJYakJultOP/XZ80BGegqO4QbtjJn4BnbfOCE9zLjwR01NCwRXUYOvsa9WX/e80
GbFrmGyjyukjxy+ma9Crl96WVmuYDJ5WyYU9ZI3yug6XEwcEvxqU1D3URMxitODw
yf7jgmEN3PGmGXSFnRZc/69i0cziq6fzS8d8Tz4pQV09Jx2zOg/tZXHVz7KGszKV
JUc1lLr9fNY68PfdpoVU4R7gkSf3cP50AI+ao/ZnQ94W4LFCJa2IL/8Xin6Xp8ly
59BkTo1xWnvmpMoUVqmBHhhDcbt5PQkfkTvOq1v9mHhoDTnv1dPn34gmYqbPo1bG
NEvv/XYa1JZfF+vLybITP/UFFCc28PVWYqxtzi0zNnTERmTN/SCxZLV3wqE2msJV
xqer/yDQ7+5S5ouRrBtMXYS+eyOe0Ip9iISDVytnlzBwEzwqi7FPGMKjXW5iBEe2
UPcAOTqvjDiL/2evlpxJKmAXeHpvGIcQ5nIZw9b8MCDvyMHn4sBMuKK5PzbezxgN
fu/G9tpl9WEAVuyK9CUoKGXowYzjnbDaoTy/2F8bea9QbJZpBzU0xRetNJzb+nAQ
juRYm7mHzGAe/FatjCxf3xIyQyZXUTXbGcA4RsXkgrnLYwxXyEPy3lCx70S8uHdL
TMGu24wgE3GtRPXx4i6FM7KMDl2i29NcJ9PmezYMuJbsjPNHM3vNLBuAo2QxipQ/
9IbCKD00XUuNYQD9e0RtB3EiypDqeU+DrM2CagI67aOL8mBPQ6ZuSlBvic+sIh3q
2zpOfu9vq4NpDTdHQmR8ndUfJUByXTQAjv9u+OV9sGyXzmjO2ZSIvguZGQVBdnBy
LupFDpZOC0GckzIyT9OrTS0UArpL5guQS4p2kfwh46KzoSkpAYCA2dULyBsJQhj2
PUtucGfMsEY8eZgQORFY1NJ5UiM5kJAFfgbDgSrt0xzmQ8kh56LqI4VVjP6yNwWi
+qY+0GiXdnPvzTU2ntQelraoYxg3xIe0m5jricdb+nxnK+USegihrqTPTlT2Oc1n
ODzN1UjuTLa0MpvPFvy0WPVbKDQwdyxQ3LPa2RkMkUuPPhNv9DHy/s5S/4rKidym
6lsNKPOoFlLPGgrq6CA2nqEGAoC6d/BCAv1DRKIcdAhAGmb1LhJVl5IRUa0AnLcz
0L6gp+wkZapb3RKsN+6RLE8qmqBTC0I4D0OD6yeMpm0kcinXXGcue/M2b15bbQRj
KHBnnNDuOWSzLl78mJnqVXiCJt/pST0gUOpiZWXp31C4hwhboHukr04CFdpa/yho
Yx5lixGz1VsCu+bSBUIqhgpw8njWHOfNeOEF6a+lijFzyUbTv6AmeruvLY5ZzCDI
MKx20htyPKB/XSEITKA7QpfYlElCDn+Lp+Oz/FfYqXGiw3tVUwYkREcDI1ksuOGB
AiWif330TQ8smfI2d8YH2n3q+KtyF5JM5GrFoAEy89zUGHdCCAZDJxuaNyDr/g1K
WnwzjKm2rHKeFlwuoE+kCZc7ow/xSW8BLN/MJgTeKphap94wHuprTQPEyvXpE5O/
vEP4WX6yugr40Pgu05PjliRFNa44C8qz0JGud2/Hm1fA3FR4go8/DhtNrTfHIeuI
M2TgWZ8cq3nmcYgF9ZBPSWI68QdmVCjt32UpXSZoRM4g09I3G7qaRciWyWmRT7IX
es3wiNf0M5FPYoFHwZsInjrC3MDj9AFPn/Xz7S41KT3/6MQj/tR0jpCvPzIBci8y
eEk2j++45qZPzrCcXa+/8EjhjT97o0o18T2aiHTVqBI=
`protect END_PROTECTED
