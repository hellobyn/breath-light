`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEkyhIrkf2Am+8j4WGGNLDyb2GLVwQePniHJ8lXXP2hL5oZJjJioKlszM4EbH/cU
/I0nr0FBVYWadRIAsM4T+rxHwXyIjatG1zTtsmLfG+Cb8MwnUnYvsBj6DbccfGFe
m/Wvee8DuDsu8TPbps6Y9DtynQjHwyHr5I+bAhNkvsmeBOoFBQWfOLjyXZPLris/
fqUXH18/kX9FGji/LvHeIyl+YzFL46ORWqTF32vMl7gYuS70b98lXTzaVgHKPSzA
ioL/dYYHUUUHij/wWQMt9jiNleALAFpzmJlPlIgK9hWhFZnL9NhiJp+qInKO6bGI
NJBPNIRu1QAofpmxB4V4A6dJzMkSCMc3Mw6jSpcqQzcpg+eEvRJZqRrvA4F3E/GU
fBEj2wwG7tVaok/y0vJNA2qpVbWW370XniJwMaJOPGApy+wfQE+E5KlZgcyO/2sD
0EJWBs4tSnm4k9TdkCR+ntRdaBDziMymMgLMeoB15R5gOb/UO8HxGEKeKY93mcsV
KoLgxgV4ToneUcAwqz0FBxuPq3CAa400DJEJYI89Sho=
`protect END_PROTECTED
