`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSy4jTig6iQ/LYk7cDIVmUKZ0+uqp9KisVClAYLJYll8boWitrApL+F8sl3xAPX9
UkN8oU8AIyFwetwXaaIeXJrQ6XuHNQ7fX+A8hxA1X8V3iP21YSGhYY90QUxPjeHZ
wBovyMLMO0vazAX4P5nOlWfM1EoDN0b8ddoIeFdk8zWGbUpJyEmSqTmQB5gj6FGM
2aOiz9ChVJn7Q5i7OI7veGEy926FJnWCCZuMpBKDZiscvbWOrygspPMgDYabjXqM
R9DWNQGKmzLT4D3djbh90CJ3ejek4dTlwyyaFtz2gZq2ZYBNhqMOaE9ir3tQGKgq
1D1OIEa1gZtDXJ+YStlKEXQ3KQxnu+8e3lupar6KWvu/FuWU4Rnb0OJGN/BE78KG
/4vD59mHsjPqSTLn5pqlqXonHyzhMR07hR920IhBvPM5SWRoh30hicYt1qY+78xH
qRRw1W/btDBJ0N8aASR89DMFljoBEtPgkAXJgSFOQSe5nDKG6OvKHnxvt8g6Tntz
lf9/J34SBnJEQbNLa7q7c7Cn/gprex0OTICnN76RM1VX1KQ6q1UVcZLw34Mnflfc
lSEnU70vfzcTQwliaZHG52ezH+QgcZHXk0DOZ05Q1MNzw9usGM/dS5z76HQBaKXC
Avb/k8MIr7pM3pDOgwhm3FAeGc531X0xqGsNtldHRnGiWRRQ7utLOLBAr2tqY6Ic
29TdbqUyzy3tMoJ4O73JBbMXB11PLVrE/00IFk7sZpMtIHtBRnAPveGBZnSnACD7
gr0lM8Z/T05mUtYql0HxDcru6m5NglYSPtPp9B0YZ/Vb4a3hIIFbYIecnprSJVAX
xtcqY1+LWFrkuO5y6yBON5pCWi+fVDMe2Lc3UzT5ZInxSu6lUusNYaI7ev61mufe
2388wEubHvyX7lZ/p3W8OYdIR8FfW1zUZpU//oItGZlg9rUQ8BzaacY1jt+ab9Ib
Lk+yj4qfi/kZveBJ18wVD3LjcJnXxFHIiB31be9It9SzmU6CO3yeZdTubsmTEe2g
KBU0gXE1b6uXYwTJKhKI9oDCp6c/4yTrBjQcH1sBfehcEZQpO8Pgimhf9uTQ2+O1
tu/aV393iyj8kZ6ZFrmvh0j1MQcBzw0JQuLb0mQMQ9P7Q2oDYpm5K0sGQ0rbDPnr
WQUN0CIm1mKCc32EfmdF/kDMfe6uZiae0tdl121f4u9Ad3Ne8EwqNKgyypguSx+o
CreMk7ylTOwmmFo6tq3H9AIuA02bwBgbifoZ3eHpp6WvsYkwhW3SVMnY3B/vPykm
GZJrjMG1i4aeAR3D34kVok7Ahl+bjzrtnspH4zhmA0BhvdDJZsRplv+miXjMAG9F
gDwE2ySNf4VWHMcv+s1ptNQ/nxu7Z3kcj25+e2pevhIl9N1WJcYaapoP9nXXmPdf
Qgnt1oElRcEtUgOF0iI8PCS9p2z4MBRZztlR/SR2pFVlb9jt42AKXyvqPiKc91TG
sx4lgF5Avp09eOsMYOp6X6zfVYsMtPKMDuEhDskpO1lLtvn19VHpNzDx6mUZrfRx
v00mwm/v677F7DU+qMcE3muE/KQt2xKRIZsiwophDwIinQTxsZRqpS44hr+j4LEg
TJQt5WgBkHi5Oq+BbHDn2EWqR8ACmCcUOsZbiTpuHgMOLU3qy38MhnBF5o4q6Zj+
ytvj1CBOL9khkZSKRJt7QFw102+NfGpehJF+f88rd+O0nVOW+laOvhjB52RonEXY
+CbTx4s0ejxQSDl4FDEN9FsDGX5S19wCEGLj+nSRFCyaXaVdZCyRX2XStEbiIOUD
wF7p0cPDBQl2Zj29aykhhGTX3Vh1CFiaT16KYwMxCD1jl6/g7ahD7cr4d5F+ItDH
rCdAV+YSEP3z+TC/4dQYYcqmFZzrnWs/dRsGe5NmkSukgwhyy5fHsE+82KaBVu6a
cBYvusrMVd9S4WL9rq5h4NvDZ0h2nUL9gcyKbUnvsKdNdsGfUEAJ35IceRlnhIeC
A3m+LKkr5kUw7iY5OaSDMPsSiP3o1sHYqxzsBFawhS1FKsrVFOTmzRA6euy6cYqM
lafXX/JIHXx9lwSPVG2qdQ6blVqszDQjv59O8YA9vyLCV2UclCZdkXHWoYqi46eL
cciERgZlXnxUFtMHfybpPHdpxMr59ALjllFxiaiPNkPIQBtZEVtvulJ5Wo1dQY6s
bQTxEqeu9W+aT0/od86JHA7sEQpT354jP8eo9e8bnJA4BiIO7Z7Se+bTBcdBGGWe
VKDJrO36dkBRrnHnFI08ZaXHOCI++xdLGySCRp7SK5Vpn3h8dq9BkJPKfwhCENiN
piMJ7lzixdPQTjYr+MGoV6WATm0T1L3X0zyEgUUfo9V6E+trHuPaAE93aqcmUklF
d62r4Vd0TsB0zfGvMx+pkajHFUtsns2zehmNw4snjJ3KsmM5nX2nI1nt2UYeA6BR
kft+x/MRHkN5Q0HkUBZrV2wCguzqM2zTOHz7vpWJJN4GKXK2TnhA+uIfxqJiN/S0
cSPnh12oXslzxvsexldIQMFhYZ+agNISlfYCB0mga5mKcQ6Q6RNDROEzrBvIoHTQ
NOOzNyu6GPlZFD1dIhahsDFSyWk1NKbY+VFyQLBHpE9gZD6Jr9r88BO5vk47hwAK
s8dYT+cRcw9Jb2yT8KxBFm8PSOSkUpR8gURJZb06IsaGxnOlenyesgFIUKtEVViy
o3DrsDhXY8gLYZTUpdl/SGwlGy4PiDZK9aSnYfFgaPwqve+dtJl21tD5uNFALJ7G
TqSil4ldX95qPNpkipdZY8xTAO8n+f6cdFPqKY6owkcWnQW8udjhoS/4Va4U9zah
Ty7Q01178jdS9ciWvt2LYEkIcRb7B0b7gQCTORvZciZO0MWKyXECX6C+Wm5v0/FS
YtvFPJ9OsH9XX/aimr2CPR3QfiapYcYz4bN6z16TAn2yiorInlwYa2EsumxTSY1I
qyKwtuVYeB2pfBDvNoD/qNrzG9BsW5rwOq2j0gUGVqYe0yakzr1pFMV8s/IzdcYo
IxqPFS4REW11NnhJ0B4EBxbS7NpR2drHtufXuYUVUwwBrWgwkoNyGOghLNeDbG9t
AhQMp5Yhdd0ingID6F/78Hgh+JfmYg+Xy1Pz/mn64O6G7NZsp69Kco7eFir6Iyzn
tZvCLEf4EMmNUFUeuybJbgDvaTC89cwBlFgdqQEKKs6aHZlhszNCrHMExNQahzfv
ZHqPzYkkn70CaKBdx/Z7Ie8KTKtJExpp4NPeGC47CPNcyO8J5gOg4Mpr+IJnfwcI
+DtDoTPIS5Y/av7ropmeMwPXlU44aAWayO5FOdpnLq5TSwH3ap9PAWLIUGlTEisK
L+2AQaaixB8J5NoQYc+mNle6cYMYe9f/kLsliZrJj3Swh9cXMzmvLt4jaTgVawZk
1x+N+Kd7ksQelNIQlV80t3Ui/WZtXqCVZTkBfrJ2yHTF7GVfPS0I5yJILy3xeS+v
1zzXGJb/uIGS6DiH/fF1JO2X3zf07rGfQ4R5Zwd8rUlgjsy2vnCMDgbA8XnQeKjJ
0nk/595y1AjCRmVn5I9l2lWt/j4juCno0z2GpTfnXKD05vgK6CFLQE5k2tkgcB+I
mjO5Kg2+0BYFLQYTA1EDBNaoLFDfOMglG7MajgEHy+jrbJIQYCkkw+6mAktTYx6T
5fr3Ira6vWMK5rOtEUQFhDYHImTMNpGN22bW/u4tcTwK8pqiBmazwMzwhMj1Xb7J
MjIS1XyVn7/zi85mTdU+ucAZmHRhhiV8CXQymPfeQnpBEqvLoFkPdcRFWifpWMvc
wFM8r17QcXgR938ITisBZ/VXdz9VWHTF5DpKfB++hbjkKYn2k1SH+5dqDuXE+4j8
rixqURr9dH9+0Rl/UCiSGHtbwLNXRP/rMw/Lu/ksGw6IZrBvjuEYWtxxRiol7Z5W
21jFyn+5CsuubpZyrEYm11jVyiO4DGVJzSfdOltkswX9Opec3ytYg6YozsUUGPUB
trbRjA9GahBHZKKc3sz9XmVR/KgoGHErBvHWTKZc5LnIzdbsyu3PuUKhOXU428gv
fDZWoXdgEj0CK8jcnYgQDtvBEKSNmVjkYQzglhhxI76jAQV9BOlvYTSJzx1HrO6k
xPVYSWKnwTHTTtTKFQhPq9+huA7p0qvdYR6DE208SqDE1o0W4xfOLNA6NZhdX4mT
oEBkdv7URyeSV8Xu5uK9GIvmZ8OZIDahLPGdvdUcYqZtC8XhkNW2LCbR8jPU727E
zpEsUp+CTgo2QE43JM/Oo0wjpnQ0EkjWLhyE+R7CMMlb8siMG8zwY2waKSXJ1Il/
mxZ2jvm4Jv7/C1N34ZbThrqiNgYR5OAOxGcnAUG5B1pFPIaHuYnRemH4JHzGMRdR
+YvVgUEd7O1banbMyhKRQvBsCJRWEdBbe5lTFxZLiQpu1iB0zlgeMbInjsTmM1P/
lkKbEGz8aOVO655cWOy2RodWmEsOSAtOz8dfHSdQp8twrkUxpwEAicAZRyW3VvNi
lLspJNETUZ+rN2bSy9iywBPhd1jKFnIkUkYWmCcDIRTL31/rHgq5SUen3+1wPhwD
JZjy+Kl3AZ/SzmKZooswWscKueJes57cc/kVpseTrajs8LXL14ZUQEKl0DjGEEve
m36eNVXIdaZV6ir+xA9vLkmauyuxeRSpXA6hEtNdwEVyaFG1VBuDjOobC7X1MDzV
lIsVpAGoueFjTi401kUqMxxvnOrrlwb4fx7Ur9x/X6id/tcwbblOCQC0o7ispN10
KQc0KN8NdJnmfP2CynNLDh489fyM0YxxEyepaoOAekSn9G5bMi1FKrj4MVCMWcgT
mFk2n5PL/JxsMMQr8ZCrTvOV0bX68WhEQQv6gaOPWgaROYUk8eLakMSgnGdn3+F4
o9YiZPE1HoQpCFAWtbmGA1BWeSHinK2W2MutAtYykdBEYSGeijmFsrmUnewITrD9
dq5vs9Mz3nn8xa9dJ67CPedhUVP9Fcpqq7yi6KYvfXqbSjbWzS8ReRzeZhTpRNzv
Gkqjs+J8mGrQv6XBdLr0z7zxZf4qLiJh1HzA/5+Qvqou6ecXO6Vn4xq1TlfEmOfB
8qp7VXu+uIsWBadyI2JTigLPLiIVJrM4gtDBMl3e6WFakFbMsTG2P0cnkYEHNfM7
IGFgUJnBci3WVwhMy5n9bEYI4kRTIUGCAZk3V862PNeOu12vh21TbAHu+5R9s9QO
dmad4Gp+T+xhtwIM4XM2eb0+XtTG4JTnswfxA2sesfEqUnvVLEnDnv0s+m+1dG6n
IGtCvdToOZJ9KwtIa46iFbPiBLkdrsTt4fvhiLzQEDMlkHLprxHdJAKEfzb7fzRw
RbdA3Agmj3nJC1TDorboOvHzmaNuCttUgPpohcbtPtN24bq9Ajmf2/Hp0le9sten
FAorAG3PRlaSGGSYItoGhzfr8CrwrXcE5xPoDLGA7qxAnOa5khoRfs/i+2uBxFdv
YjKFbeavEKUfLWCFVYNKxCJdcI1aex5p3mfWyR4CL7ud0PbKrFPaplHlVTaQURKq
OoDCUHSNQsWhUHZ0MnSyEJ/c3hLu4LgadVXLvMXKqnM0EktVJaluikBg3XnlQ4+u
Jd7TEvVNDPOzQlKtFnVFxxFWSMM0OQ5kA0T1+1Tjrvme6RYKS4wXXWtYrl+gOUTg
Qx8+eC9mrSjBoA4vSgAD3cV6MhYTjkcy0IbwKKjA+X2iG9VHBACAN7upSXcpsvTF
8Xctk9yztDIL9L2rEnLizN5WBA6YZ/8j2qgsmwjb6MGXMqxvGG8qq1iUfpEOn2n7
5/f0Hygt0T0pniKXZqorv9dhR2sCR1EIrW628/wHDd7RzY77XQxuZRPR6OsEasWA
u068A3kJdjaL6cTHHgy0U5S7bXk5gaSu0GdgybzesKFv1AH63M/NiisomAMFPOus
cyDzMLAki0Q6srr+lmYpm/HYsp07qjToH2MGyyrNpuTHP3qnZvvATeZVqQFvIV/4
Ok4Rpl3bTy3NQYDn+b2GLACBxgPuyLxwhG3F/VlnMvRxTtsWI4CtDT7twk925sIs
NCM3MsRKmhqRDv6+x9eW8nHDcE/AtgU2IoMP3RjN7hJsX+L9Jb3lk0SZLLr5dT0f
TsXG8xf0BQP8Lg5y8Y4ezK5I5P8i/K/TCaqNMKE8eQIUStgb/KArH3BLvMPX+S6c
PvR2C7uGuJJw7aztH+oR1S64PMxASO23SZV8B6qsZSZgR0/yiRJEwDXdNMm4Whuj
SAD8igrXmxwn2LMdCtuEOvS2LCmw4gZwXX16Cfsu6cpti3F7urONyQKBk8DgpUJt
+YCOQ4j7NYSldTwh2HtTcnc86YZu9s0xzqqTrkTEbI+BO6E6a3Gc8qnI7RagrMO3
pkV6XFLrOrCAGgkm9PpzWJiAhQyDYNxkqR6wlFp3Z0krz1J2GNzBvwbpOZ+JUEUB
fhODsQt3ofqg2qrtJb8MKEDmSQbJV8NUAKZSCh2y2iOQfwlmjdlV0tbKSFL8+f0H
9UqZnBE3KxcXbmDZyUoRa8pxtGgNjGojHnA3U1MUNPm6Irgkv9zcxbY/in/+ECvb
9A+rqTEyokl7izS1w3iO3w3AYxVFIsKk+6PtSCEr72nO2pYLuUWJqTL5aNkyKGlJ
D3bNxTeUtBY1UIZQZP95dNWdwAgZrgWW3dvPczdzH358sEryNwKkW75AYE9oPfEg
QxMroQrSiLL/ZUZXs2L5v59DHgj2HFSjHCQBzoaMq9gtd2LE0jtG4+ZSKu8SOIia
zXkYperAA8KoQRH4+boNx0T9mjmzkBLQcbc0nbgMka6Bsim1GfQxXygQay5XPK9W
je1RPL407r1Y2An8ahIh+hglNR+Xjo0AV4cKicGh6mBRMkgBFLzhQfmLWtMOY4lu
1AvOPGbFQQAL4EHBnG9rr5ncpyAGYk+6g9K30OCNvDZDQP6QF8hZ/074vE1Il7xH
Es962+flAzLVHisZqUa/2Vf/mLrXYtIj4Eddto8i77nLbqdnTVBBktjGlkHjyl8T
KPt/Tf1mXtKfSdG2sOQRYbUenlqdMb4Q+emusoI26m2NJuEd48eFOjLed3qMqw5q
XmW1nEQRdQNOWK2/0/jIB7dB3iXlWRnxhajtSNN5rh7/l0VF30FeTMGXEGmBP/fn
qWy8/Szk2e3/uQKWBZ1Ie8NCZ1HuCyBttulB7rN+4nRahifVvCU2GPQvGq255nvP
DZdtu+FrH4XnIk9xnn9U6d/uUQnYjQpsouDGZybVDZB7BFaNmFHwIWKt+reR/LsW
8PPi5kBuuT65XkYYkRkLlGtbH1LqY1pWURKW7wTZerPnG+hNHo5G9I8KEc9/L+Qz
vvkYs+mrZnKYQWrXD4jn/BtXedSdPaSB/i+T17GgyliDDIj6/weHkMpvb0IkX8yX
V4LBVdL/8VcXxZJans/y3gfio/bTK5Lhb47P6fw+Olg6cnWXh1D5Xd/RzpDDuzAY
LVZO6fFvIoWpN/AkHh2rCQ==
`protect END_PROTECTED
