`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8AnAq0jLI89B1iiY7tgwzWShxnobzd3krQIi7u8VXiPng7m+k6mlxX333rDmp5dQ
/IO2TGZX3sv2ustxn6g/4m1BEpnwLcyaL38FnPDewzXqT5OhnsyvL1p7K04gTNzQ
h7IqX2MlmDKn1ASp0tyBn4/jmmsB3OZmr2uuiTZoo7zSGiCQ/ltwqJLVLP9ZF2n4
pM7BZjm+7iwTXGFb7tra43fdcwOw6CThXaXF9jR/x/CYnR428iXRyYTj7ye+7b0z
s6AvkVB+c0S3ABjFIj/ai0R6DyYCkjHmtNXP9SPa2eXavnn0gpohCCQDNNil6XU3
tSmurFn5kSuh+0QOW4UEDHCIChh83RoyiA2iiaK5SYBkdZ1tx/ETkh5CCjsf39+o
Qed51qF+ygQgAYe2GuD3fCFYMOyjE+TO7fLivoeMwV0PSrmZuC2M9U3S3USTtvW6
2QaSlmAEqnx3ygW66bHIaLJANVkdEqa7iER67mkLCdxLX4cB7egVPtBliuotYsJ7
BcombWIdBseS5O605HFplGJiiahPmQuaNKpLyEJCp7klK1ZBXmeLdVH8vsCRLfZr
0i5JMaUiUzKnyzzW81QtQl56R8reB0hJNu601fPqCvrIGQI7Ml0u2Es+h0vUIIr8
Kd6Tr4SUcGT1jGwADxaVRp+Dpk8leQ+ZZtyKgH0fx9i7iF5vVMGEMTOc+pY/AjWo
OBBO3yZgVOjN7X0YfotyaR7yie35Aa9E+oq/rCCvymbypnUgfMb3dBPJ7/MEaR5A
bRJIezvSCA0lf8sD9a3aSw==
`protect END_PROTECTED
