`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4Zmd3bKhL/OIYJdcUMqGbgdXxdvqqywT/JjIzhmoyJB9xtaDsZeO7Dusquqboxq
9ivMcARw/aHqP1emTuj12+aXIaZR9x3g47otK39avVPxma7ksHJWjb2FNwN0v6v/
tqrf5lKb6fVTAX5EraQ/H0uYORWV9mlSWBIu22d6ubju/VDZipRrJbiRbrAvr4cf
ZTFzXnfUJFOoq46TdQFOMHi8+8Q4jjZV3113sl4xLOennw8O1AVIz62ytP3eC31w
8ThYZApxBgUvcqKLDcKXS18CkpBn9vlVHBejZShNbSjNrsDcef3a8sBut5kJvtu+
unnExmh+x0mSF5XuINdluiuwbLuNY0SCS92zaDYsETI0uECTbOJz+B7obByz5CcP
fG3NAvsAsnIo/pI8HMvGCXplRBgc72kPLwRkFL8WPDVzOJhfpaqLv6Zpl4rCqtBg
LxI6lqNeLg4vR/FN+gn6GDu2/GbdbEE05+besouzSqZr2a1/WpsCq9RdUGGqossB
kc/mu94Hh7MLLnDlt3vLG+lxDfHTT9mQ+3ErTh5ABR0WNEOlGf8DQiOtQv9iwgIg
ZoQYV/EZb8TIeBBOMoBBerzuQiZEbAqI7Sg5OHRuEnhgs+7WxAFlseBASu6wpBls
3PYr1kKmfxrxWxypo5cmBmLbS0D71MhtkDaEdQTrb1Qre7KlCFdzzfo3Ko0OP6A3
XFJqyrGebjHSJvAaxDVeJiYHWrXTbCz5vdK6Bi7VytV2okuhiZJ+T2K+d/B5mzWT
kmgGICSuP7rv9fq8YlgPe/JG71ajwYL4HR2IKP+A7caAaROWdKNdEkQ1g5yMlv4F
xuv/gzwzZxAtKzuiHpbhT5xHRNUakD53Qkierwb+13IYlf6So3e0oUrXwYR0RNgq
lR3SjpmzQSTlH5aVuE7syklmAmXqVr3lW1tc2VPQPFTfrwcXzCy642h5HFuoRyl+
`protect END_PROTECTED
