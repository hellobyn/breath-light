`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QU0yQEfnsk8mNQGJsCojkePLf90VhtO0+NZAgaYaipee2F2+hLgF7OqhwBVagipI
yKeRx5rVbnQ2GNIIO0l9+ImFgShydIPQXQ0wq5OlfyToKL1pc0x/JWRleQHTfPos
xsRu5mZcJNZiNmAuwpxr0hcqtuRiuwGGUycWqzUYpoMRuJyBu8jN0byqVk/siDw5
DISJiGdo+rcINdIkV8f5paryGOot06k0GhF3jIn4tf1L7IGqb4gUkzE0ljLxeghn
r8jpn6tnU9BbNPmj3HIBtyXwp6R8d8WWVoPoWZIl+vkTKOfmc2q7mj4NI4coPqxd
AGkrGPY4m/eY9tqsKxDg3Ab3peI8yzXQATvQEzZNK0S9b4QK996bl8udn8FE7P7F
4vKdkuVRLlHB9k+cxw/zB0B2FktnNyI+S1NhnwF1HpmFr2lm7hk/0nFNoUyWYcot
9sYyWUm41gZ0y+DqXACzw4z3PLA3pFUxVtg/G51QUD0Zs8k3gbedcMyFQObXYe8l
9tcxZM1070UEsUG0+dYLddMcOBntKd60tBWOayP4i1IBKahuoCTcaM+jzPwBruqZ
CUJ5wHwdn/fqYyp9y7lD55uANNDGQbYTw32yE5ClVfA=
`protect END_PROTECTED
