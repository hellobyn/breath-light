`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brFJhVnQlDq+0Azp2kaG3m2PJUWr2qGU3X0DtpSzsp8GCAprM7J+ngkKG6MKATDO
e9r3VGwn/cPhcU6Ar5H33FtXLQmhYWmFOUa6odbF2WqDOqp7b3YvPS9dKfKAPuck
OAA/kJ3hMF+WE0COKyS21DbLYhGHBeBWhIyVdbcCmqrpVCPYqKDdQBEfqWXvwYMB
Jduvfwn0B7uKO+nRIv9rP0xS/JWyw5Yo1mbx1RRpzVE93NoivDdTWFzc8GM/mtuz
lLiSgv2i38If/rjxF7HHbjxWOlGoQsv2mIZGl5KnKfWmDvRLhL8BCe5H9njLctuI
ZAdfjIb5KEX0Ru7khTW8JJI23M9uE3wXmYu1yJYpc/XLMOnvXR5OdkoGShHi1GrC
0pC8Vf4H9ZfNCgR95DEFaWMwT5YfFxHL3ZkrrHPFkdCI7hqIOCy/jg1WNyEjwkpy
pR4b4YUNq8v6uKo4sV7sCvjWG7D+7RNK92/Huh66j8Kg568nkznIZaEdCy4tAEYr
GbVgN122M2Nqs5l+EY/ddLV7LymCnsk6QTl2+fJRzyHnri8GSA/1EjeqwfgjcdR7
vCbUQafH5JTtGzxxyLXu3/qTnaQWY+DbTdYAgZqCLLRVLkG0oEhuVo1b67oPyMaj
NBbHQah1ehqgcXguMniBUg==
`protect END_PROTECTED
