`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct/hMj/j1Adrx6ZndXy+WFvDa6SpqVt3Qob+91X+DfIGMBjNfe3uHqke3ZIUg5mY
SQYr9wKwNczAPfs7nA1Z0gof5WkjIKA+ZxoxxzontjI39oc7NvJqWPxJp1WZTSp0
jQkmjX8Kbxd922h23QTBYP9uoQYsJTVfdu5TtI4iDVjVo/mGWjAuO+OyZrLCvfuE
pxVRK2GggMcChxD2RoZVtJKcEORsS8oNcqu0nsqehZHosCBIEeUhL79tmMrVwS1q
u/HMjWbn4Xx/coJ4HqSQXPcM6zD2cL6NDZG+iobqRGLUlOwoA9pDr/lZHiTL4wYr
o2ix9QlJOsN0L95tFa7JshOfsCMM/0mJ9Y897c/doV9Z3tW4MdAReCT1z45JgSAI
eDYAJR1U4kxh+fMVvRtWNt8IzLkCzdxz+wkGRUVy6ETT3IdXU+sMitYaCbtix5pf
6mu/hP0hQ+j0SYGIfRRTw98u1IggjZ9f5a4C0UZRunD6ftGCMh6lq6ypUxHnb+IG
8gCNT9+AOq6Z8B4ijnCAiaN0oVuuXw0LLyYKu6nr0m39jjFMW3D+RC+LlChL5D5t
BZy5ZiSzzuFUTikYzbPx5RMB9WRrTHjOJR0VIQUCMDJp2op3cpUjabDpWeJe/3JC
iRK7mwRLnh8ThizMNxu6+ozSrvI0jXDi9AktvVCV/etmR163xZ1unnmKF9OHV57u
FUE4TdTmP2IWtvstkiCrk6XmkWUux9fXw6uC5zRTL7UFmrso6OGQOwabJ1ZU1z/o
71h7I1yRwpiHqhW9RjIgxvHrheEBp5jE8kjp9HgRmIk2vleyG6tkQctXFbkuVuYa
Q+A25YDwdSyUET+2zGjYx+uPCbLXbL3bbMQaS1ccI0WrXT901pmQ1Xk076K094cZ
LYpfVD+oCl1rDmMcp6e7RjJB92e9olHdW51DpUtrOBlJzzikk0h2gXKzCSWW+W7x
aaNVpUVeJf20FZUq5GRc9uCJuXCnV5Y5MR3a/HcQgqw=
`protect END_PROTECTED
