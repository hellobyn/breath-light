`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1oxsLlxMtzojd0ad+qb1SUIwKZpvZZt8Yp5kvZ0cvHLxTXr+WWxoUpCvakj/3tM
EydpJaZVG9XxAZTYpr+A/z8YXoBMWOXRshzDMG4hYuXvku339X5R2Ouc7yGudpa+
hbn0JdbejaOxewwGEDxCQWClgABmS1e5tYHNWoXiXhMzD7MdbeShpXgkehmFFiVD
JEDlqd2jznwivBRlJJLEP9nzp5BKF/IfBNuyXdePsx5fJAz+k4eHvQbr51L4RBcT
UaUrgrYtTfbOOa3Rgm5etLIt4/yR0EM+UDMcztRYAfnubD4oflISrRxLrzHHCuCo
jIEKq+MPnMREJqHtXUM7cypTpn9sT9pg5sAUcRk2HIVTBpyEBfYefAcOtPw//7AJ
W6zHf+Jf8Np5WmbC+oLOIUbnBqAFDk8WVanL/ijfeNxmji62xJtjp1+H5OjHaQ8N
prEifuNpcySJ31/UbI7SY/f6M0ZagQpBTmSiiTptdiA9lYLsPMYcLPxeZPPf4X9E
7nRx04KfjT4RJWAHAwoqhhR+XUifnHe9dMRc33ayBt+Nn22zlz8F0oUAalftmlRy
S3oBA5kYhz+iQbkJ+oJRIv01y6JCwKrqsIcms/Bhz2AGVS8srXOtzTdvkU4D7Q6a
7sEt2gcQ+ZQ8z13YUjKwYh1y8H6Lz/tUmj+Yq9rkV9XFv3t/JiiOzYN8tGIGOYkh
GxDZxHrBikqa3UgS583TzinnEBB2KOn/aAkRT19QNkucdqPl9/lfMQdXqzxDwPhi
2W8b6dKAuP/FSIsqp8wLQA==
`protect END_PROTECTED
