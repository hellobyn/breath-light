`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bo99ZyHVu8WUUUJ7I9ir3uvHG+IZhAZS/xSLtzAevOWVv9z+eG9EEPKXCuujrRRm
tWuZmo+VWkcdP8ZaIWKAtvG13XeL6//PZOO5J/e4r2HJ75MHn1XOuavw9y/Q/hYW
qLDnbPYAnAta7+7H4ye9PfJ8OP7BC7UTtEQ3tDokYZ6ucRzY0WonMh0/eKdp53ue
zLvpQeB+gazHunymHjTIdZ7NFogDxE972tCAfPrhb7WHeDk6C1NLlNzJd42YB5LH
JebzH1AvDShgLT49yAUirxK50OKNgspyYK3OFFql2LHUiEXyfDxG0GW8Fp86+7Bl
ku9SRRLCAj3wxNlY/uuZfLVrS+18UqKte9RIZn7MbnDgKXQe3sPt6lxDwLVfG3Wo
etFVILKD2zeJYTzAyosCmKVnmxY8d/op0JXdy/BY7jVz8QSkSfsaij+mSSUfyjHr
u1yj1u58LUW3Vk9OjswA2GVHdSZyuBQI7hdOmE4sfaJmCgssaMvIF5b04ATxUMk5
CpFKKNlufvQ1+V+KRcupX/CWygaiYJfoNiAr9HRTen+Qy9ZcZI4ChXUPOTdobfM+
ZR6KvzaOvim2uMGBWNhq/suxlz0ip8nazRArhBYz6rzLkjWrnO7UUtvvc7Y7VA0p
HCkaqC3Iu1RfbeyX6JLc5cjUKnglQuqCfhqVLz0qb5VTHaU/xLWz1LJm6zw1grWD
8Crt7nD/BkFPF+dZHMbRmCBG6EHweF48phoUOevjlNgWXBlk3fNONPaYN+CLsZX1
tv8qRtLqU1v3ejcW0oo4VpjfVBUPt9P6AkWFmvwcPY7bYcjZTUAbKx+VXFGDvYf7
CRTIY0AOCTfw93OUoIlTAvdvUBqFtWZuOyB0RHwcTkkdgRnzTSdHDcjpqkvKhqCG
nmucEDe4zEUEgU0DFAN0cqmIgc063Ifah20Fltq8Ke0bO23zbjenU5vVot0OIOTX
StuUUia2psBpFtZuoF6D0TWodcVMT8a40N3X/umw7XjIEmBJe437Jyuh76ru7UQq
IGDl809Dm/B00FczzWZQpVg98fRZ3AUGuUR559V+thYm21yCk21xGYWxnrxeN5P1
Jszu4YySO6PzeVL5nLHejnu7w+BQjDAxDYO0yglOWDvBi+9I7Rp0StHiIGC7VYNV
/fuVghc+ew/Ona9S+TAt/a/qQqH7br9fr5tuiuqTcpaHyk5szjhP4GMcxa5OQ83J
XLpXc5LTlqmWCFAYbhYH7mqSm5taEy0X9DdAggOY4Hg/0AWbvUoHjxIGYQGHTQ8h
p/1YYGBtePeoSxfXP4OfJrZtGdwqXe16txo+x1C8E2dWWoIoYu4vgwAYDIV4wwP2
cpBBb1DonrnoWzEIBVK97T2F5dCTfpgJ4EmkUgz1ZO/8o3gbdJS7UYiKa0iCcLQd
p6VQ/uidXdlE05rDiuaMMTUIzKJl3q61oZiCoVkmEj/ncqxt7OVSQlLDt7O4JWQk
PxsOWLTL6eFSKBnOGkA1k74J+IF7AXJifNfwk1/GOdrifNCssBjof579M4tNPYSF
rEbaWKPiwJUl/yMTL7YLf+YDElo8u4/N+AmuRZQPNJ268vRIColFGyvXAd8tA0S6
2FLdVmFACeCZr0vV3bRFIZE7zdHbZ4G2w4pLO1O7+uoRetJlDY4NxGEqDYLKg6Sc
0fGF50B5ktfwOn4PBrfdjGBc8aR93yzeFX6s/BbbmX+/9p6ju/5+CBnW0Z1k2+q9
2hZKT6z+wBAUGieRKSzL7k8hRAEIC4RsCfjd/8MS8CKRQMtL918rSVGkApuuCj+s
lmF1pE/yJGbO0vie5apZy7Lni9qttYaXsDd/1iJ37l4k2YE3IRZXhmb8OgQunW3q
jO0KDNvFFTINt0eA3fEcMji+Dr74fxgFOnDcGqIFQ2YHe1o24fkPXoS+Q3wT3LKg
D35fHZk0R2qWakK0w87OpxBfSVb5cRvtwgYN385hBLP1jy4ZX72kCKT3nx/J5Vgx
u7mc7sn4Dr/vzb5gVkmXQRSxjWpzChcGcBeNRldN8oD3WzY+05+dRRj1OifgWI+O
RVpJsV0INTcqUwUlMWFKsS6xWzmmSB7C7MHL+HqxAlEGPKQElQLFS9X58ZUWCQGA
uoHPLwNC1izPGgOWKEyFkuNrzsNm311ksZlip7zMe89Oqhehkh5/eNMVZOmvmWpS
SSrt5vjW63RFtfa8CcHir7to4v7Hz2q6RujEtdx1ayCGCZvaCCkGn2GqlPocpr5v
72ynOf1NParwHmwl8/jqikSreEgavrQSlww5hf1TEblUAdg9t7vEFFmX4pTR+VzE
nAyTe2OCTT5n9kZ4YM7RssE6n0BehxjHbhTTvr+heTW3Fr4uqfLFWAFm+AvEdseM
VumLcx1N2oFyS355gQ+sNwl4VuNTkKQUbxcERjMdmkulr5cQ0FI7n/bPWjD/kWzL
KKKA97NBrpdR3exzyEln/syLkXFGQJW71AJ+gjVMU9iHTyFiR2rYzHow7KCucfH3
5YXl5pfg7IM9N2usa2LH99PLT3dGmO/hZq6K6spoH9zJWzw/e1LDHkaPp6L2vpKn
gArstjPJS5YGu+BSlYtoTPqyo6QHffzOf5Uqtp/ov6ioyRyNdhUfOlH6nU1sLLce
hNgC623D8sFeSS69Y/roj0oHkKCr3iaslOXLOcFF3j10AVZ05EIOc8i+uFDOldwT
rybCJ1PYsh6QHHuNN/ASIIkIumPoxOYWasQj0xSRre68VsEtpWDOMwuniYArfyJg
0pWDOHgTo54fb85DNXAmjWGGgFdzrmvwMYlc9EGI4JxcpARxfZrdj63KOeB6w3tA
zmnw6wj1WFzy6MIsyAixgvkj7FOSyVS7mCzr0giw5uLaXgavFgutCj/uXEcOUBML
BKFKvoTAycvklHTdpbKew0DgVCwasPUnLgLFW3Fp/LnEmd1awIQmFsVSfhsmEVoa
a4pNzQx7zCAxQ2a6wV41WKOUq/k7mBX37fpamr9tPbU/cxp2hcFax/Gb49r4tsZi
HgLECJKG0wlWs/fYlJXKL3bqtD6lUs1iNvue8jDra/F6FnrKT0vaQ/Nq3qvxvZLM
75vVXCn73RQSxstqUxXGbhxP3alUrF9OCS++6DQZXPD9nhNgUl6092Zdi0Z3T9ga
O5JDndvEV0iBwk5KMNwdBKAWd5korIEvwzXywRMTyZcCZIFa+jNA5KBkRUVP304C
n5jV3R7YD6OyYw8aFvVLXp22DEYH+vbUXghWHYlPSq+AkdIGMR7T2c64WaAwJ+xE
Z2qBySwxeWV4MQliZ3tYkQs15yFdpTVHkEFkzI636LKf0gTo2L1soavIk0SpVD1L
ZE9/hGuxQoWqrT9JRdB3KM29VlTomk7C+vzpfTWQB3hGN6tG40PjTQkWEELjkDpX
/JEMDAYIeE/cxZosuwvQI7o6C1RKlbvC2HC7XA2FIVnaVsyNxxJMmfj3pTUvQu9g
6c9Dgg7/GFJ8e8r5jmAH/NpcodV+SiEKnhWmJ/IeYoB0IWNBz5t+hB4URxDvXh7D
s0JyqA8vi/9mqjPXOZtkwsR0r5rYK4DyVThrQkOCsMUIZqFpG+u1dL4NKF5XZvjb
NuYT4HkdkI3RVVzg5TPeZ5epzNlmqCyETRn8ysUK37E+mOeUn5hxw4ia4wscWwN4
TXdtfkdScAH1JixiO9xggNQOORV+Z04zOZIF+KEbe4MIw8IwWVlSuKt5AfgN+9xC
8Luz2nboO5YmhvNcF2pHekoU4S7waJqpz/QqJT7LZKMLBQFsVnbhFzvBmPN2FxC4
Xw5uZHA6tu6ATL9d20JtXowwj1DRVfPJcQvyRC7JFTqVNcyfSbAjlhstgDUQ476S
yPO+LR3yAwM6Z/DOE+ps0JUYl76Yo6gpT5c//oeYbH1d973T5MintI4nO/E5dqLy
45tyToefNh+2H7aMxBoifIv2EjdyazirtkScHcBHSimu8He50ffkm8U5dOnVKZve
0UJy6nqcpHvQhqvSDUVRrmpdIU+plngnig0K1ePpn75f7uzZDGgxLxN5axvJOyio
sU5g9+Kd6ojNVP1yS4iQ8ctbUKRCuX82iDc1k1ysY5hqN5PwSOG2H6d1qC5wHfQ8
1vwUEIufkvjC68Q7266gpmVKRUwJIlFQFUhqCUH87t9MLCeR+lrNxQXQ1B0C9VrJ
hgG5RPbh59AtDhfQlXRzfLAkvnR33jpRVpdTAQogqABTIbzQgz6eC9bkfK9dof9B
9TgnJlhMal3kD3GbFYoJLBbU9cwQz87w/9aWd4EJLi/fY13ruGNp2h7nwCFqq8E4
d6wlw4SBa2T410MHai/Znz0Vh7lfInrdT9a5EkRb8NNWAjplaoLxqA92Qk8htt5t
FYnHB/s3eT0fZUgrpL5SYJi5tVj5ElBYO+/tXekDqZEuFvqcstSpHzE1+w4tZHFM
vEWKQjFtjIw1SBfnW4xBb4gZs+1KbhDWPp3cowxN3bWPEhHiKoTiFa/VTNb4ns+e
6x/1jjbGcow2hu0aqvlLtp0um72r3TbboZZ5ZwOSykIJNmC/RJe1GL9qS2QRhAdw
fCLfu4gjeZd3B6lyzYNrvkqeW22fh4Q3hIiNs/qgIrWhH8Ud38kLxPnmx9RVsmV8
87JlbIlbDIw/j/nqgcS+NcnMPEj6sHVc2dD0+KiIXyv3IL+VsLAZLgLKX2elq/wl
NdOnuUb79CM++jE6vYO8yq4kn8iRYT1R8sDThVIeFnbHfOhZwqWFOlnF3TVZNjem
WD8qTV/LpiaxIfZ3qZQQOl0zjuB7NEUH5O8gq+VBv6waGqlgvkcltRWKShzmPSOD
tlbStg8VSSWuaqXg+2CObWRYCXgVSk1wvmmT4mvDoETQ3HlF1jj87PZtCFWNnEB5
hKkn6zXS7V/iFZ/zMQBX8OFfH5v60ILe3MYwwg6JoP+cVlWlBM69I1v3NLzlBYK2
yijNo7V37AXAznpbDYKjC7f1CLXKFKXUpnGsjExqc18RGgQpawSH+Nr7/TRDApnv
`protect END_PROTECTED
