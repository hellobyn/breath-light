`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6dMoe2coIhr2Zr82QM+4DmNWX+7p2VoBbMtFSbEbIndqwQwt9T5BbY3b2LmPByi
bG6YrVg7yxWZzDT51Wa5BE7lGMujYMlJDkz/EHxfO7exV8Un2GxCzWrrUqb2lDMu
V1tg8/yyCXb0/J83pLoAOh2IphPwlSjJoEnis2qBizVtoUzjwpu4M6bCAES3X7Nd
m+4htxWRqnb//vnNxVQ/A+15TnKIQwp6FhtRlFasndBwlUosfeyxjG9PIU2/5h+C
SLsk7HdWVnEmalm5tZnv+BTMFAoy1ujMqa1EdjcX1yvmyIY7+zOEHo3CTyI992gj
PoloTXg/iM80Ew7LEimA4gfKKAmsfKH35DegEdAcws6KX9trtqlHeZXGrA2XZFuA
D8CzBK28oMhxtr8wILJKy5/xEAK2HcEkkjgw+0AU/YHEKkGsss67JcgXcFoXMCeD
i1AW3Kl+8Q26flOeTAfbi3pihNjpkAb5UPLIHb3Jxmtc3x+56Ku9NjOE4wlgD92i
XO6w1+MEwugp0I7ZcEaxHcrQ121MRf3K8+BSNQsJ+2swYYSEhLj0KKM5VxuNAeAP
AI6+RUIsgQGnNvkN+df0tHFD1iKcIJjExUWe/+P3xYevJUnLbzz7LIRWWK8dQ6z0
iSQTx4k2V4Mef6aJOqCU2enKHBTmcCMXGQ132/FWzbZ3s+OZo5Y9B/pctS6Ddr+W
ZiXX62EK2zVKKCNSsay4RBDHcuCnRnZHS0MAwXFKQCoi6uIYMxpsCnKP9cxJUA/r
SJZ9ykrOu6eHmtT6wO1GXzu8wPjlz1oN4OhItScOnZ5BYRJRlkXyHGdsTGNv3ok6
T2qVZHL3RzsvUzUE8EcGrT+XwOwL/XTY37myHDazTDdp5rpBw7sJ1CKZ+2LOOR6a
qEVssyC/RkAaTsxc9HgoS2Ekq4lqFrWE7oXGzO33t9bOJViW9NEC3RmmJff2PjJw
`protect END_PROTECTED
