`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kMacGPQxoynE+SlI+LLPgcKaozuwDpSHxaVvGDPlaNi+h6zdVidHoES1lLAda4c3
6J2ifWjnrccPavkBRLS5OAhUZFGP+sk6zmtxjSa6jaR+XoveVf/2vMw+HJHgEKMk
G1CQI77/4bL/zFLFvho/ShVyN+3N0ob7vPEjJHSIErMG1ulFG5Z20uccRn4gCAFS
77lWDnu5c/yl6JkpRTeCZ37DXvwCgi5J9F5lY+CCsOPZ8/g4RxFFJDSA6TlTnPD3
WiCZKMpMtsF0F0UG7kBkstG8InZeMFJ+Vyq7aKGV+Rbjs+8vxs4SWRRr0K0XL8VK
9z271oQRqgmsZY8a0AKpKTe2HdDQH/pkMQ7GK5xzx6mzZgT5n9O4MCmWbznXkVxj
2nrZy/5oqXghQQUD1DjBZF6bWObioKtuQJqpmqiwIiVgq4OmGkE0unNvg6fJ2SUC
VUDokpn3GsLNSHizplXZDgUvqCgTZxNpwEDdjEWwcIL2Ga8CEAuDvi2PGLr0g/CW
zsvf4W2mcvvqNynbPymxO3XfnmPqf0Us/ZlxJ17K3Np7P+B3LmigQAlipgkgbjp3
+TI+gPWSrrLXZYCNjOdN8di4x28+1L88nxHMjiYsmjUnfFR1v46eOiCR5NDBnxG7
Vfy6gR0knNIdx4skChWRCF1LX9PlqOpXj9PQwjgSw+ljKZrNBcDoIZZEaca5A6Fp
PF+kiQJVaroWEySgcxCyMwQARwQ6K6vMehm1CtPHhvAcQWQvDDzwEc0pm3ybjKbk
5Uy6qn2f5KnHsQ5rO6qiIHHvohzsi28WPLbsElnfMeXR44pKpo3Q2YVl7luVrw8m
4ufPNAx1Z/LqMnGIM7iye3DqIhrLRMv25/sJlQ7YIJhOOAorzZbSxe8OD4iBPOzB
q8vWHpyUtmWNiiywxs7vXBWPFPU12st+AG2THB+J3YK+zWLlX63tdQcy+CSyigAK
MsrtnG5cqLyM6ULaswPiQUXtoT6crfNfVUAUh+39ULZFvlLoZg3TeOLvuRIP7d8r
ukhkGI69UNMyB4lTZ7qmgXKhr8+z/UoI1pUxig1SUxqgf+xHb2+4CZuY6N5nMFf+
XTxaJbGTehQNyi9mKmkfYJobWFGAQT4hLfXzu4FO6PQ3je6D//bg+7gCDadsUukZ
HGO9y/qmv8kg3rIQlYYnEtj9XC11rBe8UhEH75EKp8dmPVRGeT3MYXCqLaBWXyNv
xkl/2M0Xk9klJ89cw/PUM3PjzGQnlxTybn4dlsrblqrxMa/2WD3nUQrUbECCLIjN
wSzZhIY8QgQpC8HI2WQvIUsVsdXUNSLqb8yUsmDPSf5CB040rH9E8r0oaxsE7IUj
CZhavDLypOJfnKerKzFq7iExbtX00eiK//hLZslQqixYGyrzjC4Rz2l4/wlbTwPH
n2zGSeWJnRzyIsYM/p49rxDhnu5YeuvrIcy+T+Xskz4+yA8Ly/As7IXG/lOYkio6
u/syLCtj1ILu+QGPjti4dpIvIEtZaX55znMWhfKIiOpG7o0dwKY5jKDvvAClORcc
DwlUS9+0z5+1ulkO449f4uetHOIRdeTu8iBCBrprfzGCFjXIjBy5i0RiAEqKzPPY
tbiAG9EfOGrjv40LDPmmIjep7UipbwmleCCU7bhT2Uoy8W4gZNaQhcYcwLjDb18n
0+ztFugJ3aP6emgp45a2WL7Kv+5rAIs62iuUQK+BiLn3wdmXy0Xd3vBtzS1FN2Uc
SaJsb3I9Lo9Yy9HzPIJkwqo4xs4BfqUhWnDc/39hrVTljqYnXo6F2+B8KhjcIx9r
0Vsl5oyLBPEcRqj0EPPaE0+E3EEMBaOIP8Fe2BEyj1d9LF37ELH6HmGG4ZsE39oW
Cf5us+GiTNJEWqW/+UdvdukiW6iQotu8y/NSyvqPcuNKv3+4hUf6Rjn7y6a2eWIM
SCfr5jpw0LDw+qlPjwxs78jx3jbFGKAsLfufOuRskSUfK0X4rUONbfhhmpWGBRR8
7p8oTEdNjYKsVP5IvIXEYSrMIuAjoa9FrTAu7Awlr787tYidh+T2ZCWRrpzBfZfc
GGUAYothfsgdVR3NeAz0ALhi1ZGj1Rh0pXlzHzZYTB136QWcSFkOeDoGWRnsoEMl
EVD6ln0z1HrnvRAVpPb1fAHuDtmIE2Fq3GJd8Dpl8F23w3bE9glilE/eh1qZUpO8
l6nKryYhGa8FUkoU6uBFKsimxSzQR8pVQkv+8JubOyYtTGcRaILHCE3J3VVhN5P+
SZhmjCReC8C8f9od5wNvMqbANAuaMQPH4W++QPZWXlciJ/zJW+YBziFbHiN/Thb/
cs+3WtGjcz3ylBTZGJKn6iPmr9y9SmWgqG54f72yhUrjnQdePmAX+xNwlfX9YgQt
0JBj1wfewMBcOhRbwaHJy9DqaWtacMjAD41Adpdv5lWJiu1luDflOelGTlOcw0wg
pU6WcKEK/W+mo4syGDwP9fH4Cwdkbg6f+bCtMBSAw8dbkaStggJgOktXXXAJoLid
2pDQXmC6iLFm0ndfp4Va7mMTKCgMRVLYK6gJYxhsmgZsG2CxjwOrYm153aiy4ATz
nJPfBZoYVVME8kaYCjmOPBkOlA1SYC6zHwz3QvP5lCDr/eHjPMuWk2R3lvLwnLEK
QVuCPHPTMDweQp1lOto6RpP/4jPHNX816nMwG9MiqPYIZMllvxVShoGEJ0xohq9c
8uUHRXWizdv6qG1u7wNdpZ2Ky17k2q3uGfIclORCAAqydixTncEG66iY4CTiKO6d
frPhesRjCpRuK1w9f98xioS6EhzsNXkUaMKpgNPLzKOcUT32/Dcr4QY2gBrbK1Ur
bg9ibhE0LXzbqUScGRZUQUCRMh9+KPwWyVCfV8hYWY3XFjPhRVbupieqIQDDfOGZ
tCLNXT62i92KWADT+O2er8vwoyASOXhcRPSq22swO8sjHZWYGLdG9+W9Tf2sN0fG
KJKA3cEKmP86wptNqFvK3G1i3+uynBNLsJJ6a8dbUTKfXD54BCH20gd/ECAQBFLm
S5eUsbxMowBe3wulzuJuErbcdIHXcYc7AghJCDOPiZ5b5+G913IBNpazV0PSpvEF
4vxavpgQ4vsnqBDD6lnsH9dBuUCccx1jOfUU9DIHurRJ3uGAd3WzH1LeoQbq+vWT
q2BGxgu2EPdDwIMCtgLUUOkCBb2pqToNAnxrWYIhS+DBiCKFBvSackU850wE3ZCp
5odofssmtuxdflqpmvGmf3V+yMP52a7ImVkoOd6er/t0ZP3oqnDJZJ+TrHzno5sq
5OSaVsmXUvOcaRumMsuDjhU9XWyOE+pniReLm8cpugZbfpXpI0ouJ7kvxSyltW7F
aqkbZmcV7XBjuEQs7IF6IkxU5I9wPDEZdIk+/ZzTtrq2SHspRyfHPSECvBTLGQ6S
C4Opt+XeCrIhz9ZyDpaWhFPN9agdfKVCok4kf5g5HOJEzzvAsCEkizy7vQLVteD5
eqLNjG/1aL9MqYuzp3QfEHqOhsQ6SejQswKBH0/UjoxjKx1XHmEGl8hs6vtUgMtB
tMUSV9dG5H5+a+SEyZVHRX8+QZidrV3oUkUjpyJLl+Bv0GDC80ciz+cEjFHsaJE9
6TLar+/j70sln1FuLfh+BYe9tGR+cXQWLMBU5Py5aEM6t+yRdiU0t+PiZWGHnQHb
hFuvJ7M8pFsesVWshhtw8JJtNNesCYvdgwGgmEPzS+Gzcf7tAF7TCcggGO80T9F3
vJQ47BEar86V2gh4sz6HQrLuSwKJXbZom4SLfWhjJj6d1wzG/aWbKZHkWO2j50aJ
A1aU1xsXmKiz+4XWrxXrnC2GwfKxROshtbVfs3dfWcTwySmetah/D4evxuJsnCG0
ur7KoLOWtm6CpdPJKogx6vrVQh8L1yX7kXupWGs1sh+Bl9qj97xvZxUCGLrCAaUv
WTp8Hq67FBsExNeQts7hMuZGHsd+9xtzUb1T6nD8nFQ+tGUCxFs+rYPTOQgvtONv
KVl0LJbqsX4+q1toPa2wnUaNVih00drrDAn+/Cs5X8AUGwA2A9BJFBo6rR1BCKS4
IimP/2e2lSrZUZOtthO+EBTbPpyr3z5ZrYQnwSMa9u10gq0z/DltRdyS204EVDla
KH4kwOCaQHzkQW5MeIFFM7F3Ai7Bvo0gIzFTCdJiLdt4F4ospxzcwfP37z77psGV
ra841sOFZc60iK7eoTM91YHnq9MEakOzcGFckVSGzCW4yg3bsed71yhqh8xaUvST
yJWcwUfgwL4rhAFY6jTjzUfFq4OQezovSPamZnW/DxF3hzyzA4ImBH6CNgGyRmAG
hJpJYl257gkBacZg0y55s1MWG7BzW/WD2PpnxqZtcFYiKQ2FQDTyiVl6aT9UdEJS
GBagOo0SWjpcjpFn5X58HUJbtnawABgMfwBNF7JoROkFZ8cmXbYssc/oSEoBaPX4
XQ31s2d/c1KOPph6nMJPpZW9SZWR5o0M7Z59hcd6oVLR2xXNoyiBbegdnGZv0Jon
`protect END_PROTECTED
