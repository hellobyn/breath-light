`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfiqKhVMBFenkh1bsCWX9FP5q+U591UCmAirLSUg4yGmvqmFiNw37G7lkDHWHuwb
8J7mXL0cygKos67O0/sD7ohUQnvUOHukdHipb5ou6L8jn4lbtPLjyQn3Rk+pkWNv
TRwkn4K8Qthbv+sgSt+qjNQnUF04b7SCH+/uj5WuF9MNTjQjYeCPHt/ITzS4czl3
+HVj7Xr676+kVraqCaobnAwb08wuhtDWaLRUgePIIhIf6s+mHpCNCm3pkrYfky8L
cXoJQDS02nXe6jO90e9zRcmNmd22EqxGrEhZpI8t/kGynmEguNUlTBaxw7cS71tj
jpQOyHWP3XtSXdAu6Ck7KbeoU3RfZr92PqOt4RU8rlGEB/RWz+pOoHZblb9cGaWP
uOZrIODy0CWszIHuoqmASC8MAnDkiHKQp1oYZfS7WGhg34pRR3ug53RXQjoyLLR/
LFTAlJ/YzO/CAkYOofxvC+envDSPsAzAJQbrkeZPguurw4Q7ljFpM2h30JNOW8zw
smBJPpg4syJL8jDkt+96hzhVojq/p3PZ0eBBZdleNVO7H9+7aXsHvpZGsownH1Es
bC3uBOZrSSinwk0cFsxn219SBQZu6BnzhTuM2L5mgnOnp3xTklUM8t/Vj9P+fah/
BDOqOHla7MGwxdUPOp3TUDzdWoidsZptNpYygGlbtJLg1i1V4eeYSw0XrRD4EqHx
B4Pafpq4aUjqW2mGKnjD5EFrHQSWgQxgI691HLqp7vQEptfKCyDyBxwxDusFlfFt
GvOxmUmJGbUjQaEQ7/X7t0ewCzFxHUQQr01TmupkP1TdxywgSH857uv7DsFQaX5V
4yxrvcZ9MJ5jvYfPiIAQ0VumOHMIDQE1j+6c06r/dnQsYJO31Z1EYy55ymzXK0Qi
WG04eOmxejTOnSgqv640lcUFAuYzE9l0OySw3TZpz6jSu/lj+G/+WcOg2tCx/xgH
Id3eX6ekuY3xjLtm8fC9TPbP3baSSlcHOysX9I4Wy80YFVYHIsonU1RdwnuGeCH+
Nh3nYKUwcKAwPC6VsDT5vfiAfSMeKYriKTpcUocEufuDzdUVoYzgZql1K6OESTOA
6leRjn7F2weVjOWNkZymbC+xt823qZ9Ib/GxgELwbgnyT+HNGL/c+hPM1vr3r4x0
itUMDEDue0VeFTK31kZ+xWeni4Lyj3brQDJCmT3bX5DabpCK9dQkuyxS5R2NGeK5
Mcb55BH38ngXZP2eoS5TYQ==
`protect END_PROTECTED
