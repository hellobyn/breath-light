`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/QSBpEPED2yIq1ImBz3mOUfyCBhyA/5bTXp1Vp06KD99SIBhjDMmwk3m89LdVDC
2oDNxSte+vAzGKSykh0cl3AKYMMFXw7Q3uyIeBnM5g5pAcg8NVIOUUqxdKjaZA8D
nGPA6bN83ZwC0Wb+FxsU6gLVGizZlrHwC4DRCSzFLLWcJrnjidhIkqyX+K5IEse5
qXCrbrd38SJA6UHWsnksjCcdblqxv+RvOhjaOnjJmY6XV2BevYPCfJXPKZo+e6qZ
jP7h5LHSqovMT9T4Gaa8rljlkA8qAJosCDFm3Xfnsh1vZXKHD4o7htqfXYJRne5z
fZWN38wO6GngbgTMv57zXgYBOuHb4WppSiNHJZwXWMcJriC6DcXLZiVfyLWvM3q7
S40s0JGEeAG8hH0N0hGrSPSfRjVCOrHU1v9k2fr4tcGz8bCDDo4b3HaoqN2+E4qi
5e8qLdqtPsU0xx/bw4aQTE3w3tc26uXewLQQPEub8BfXtXihjGrq42yQBEU98Xkn
GisPSeCmL+3dluJHC4op5Yod0bjJX5p1Ql+lOfy+A8aRREXbPsng+53+zO740rGi
Wu5p00G+6OULH/PIG1c5TnLs1lToBUeleDZNq1pkUbLqDQuleIXJFzhc1BPYvqon
wNbzlug1z0I2Hv5h3djOK/C+ZuP+zu4Q5xfnlMUgDvwHxuwzKD/gCG2D63UNe+4P
1uG0b+HUPKtNVggDDjsfCPZT3Jsh7iQiROEU0aS+qwtpuD9XB0wUn7DTAE5f1WPH
kjmoILNrg7Dfh/v4dDUntUODGhOi0fdxBv45aXTss8trDbZITKymZUxPFgtQEc7p
5aXgNF2Or958f4GoUI2vzlfJwFhQvUGCZPleYsJC8ITK/HF4IMOoNQYLOfU4bi8w
qVhnSDiS2Eh6Rv4ZUIk9RM1U9phB78MLlKWlvE6QJyIi6RbrBDWt1RX4Zni9/dgh
MpWDPIvHLw47L1+nDEpSn08onAlCh//t/SM35inf971I8tpzEYFT8WtI7bvImSW4
9fglaRMnHccgA15EYsz9Lieby0/qJbkBcpzGsEEg52/L9Eng4RspLlwHdcxCjKf+
ikSYIJ2NCFicVx6JYpEwuqLNK+t2yJZ5lGQpJAgdCEvMqJSILTzCXMXa1FDHDkqp
M7B3iJ9AdJYKwo1ATxNXuiHfPpf87PbQa0RpsdeonVMiyRvxZ79BX489sy62+juy
T+0W24S6BhhnBvr/RiJjk6uWbeFfe83qLXGOVQJMgpWNQ/4WkQl+qLRMd9c4o0PA
ALiqOj46DJK2o+DBjH54eu4Jmq1hJGiFqbMh2wUjrzgomwujsiPQRYgwC++D+MBn
zKCCMSVQazj8sf937Nsi726ZUdH4A+stUqyG5npFAXDXj1FTGpIVsYrU9pqU5ytk
HOGBqbduK5h6+V2O0UsAcSS6WSgE/IVhfYQr6GhYyCQp0TQfW+ox4CnHhZjN0Ouh
6IkVvtX7yLn0S79wdIqihWhQtsy9P4cXMKkpa/WDJq6ek2U1C4Nq9ty0RiTJIhR3
7Pa3WtBlXEBUcTIjKraluEkNL1c0Dtq4jzECD0CB2O6xIuVVOimB07EiCnGyNB6J
+5eBeikUQ47FawJ6lEm8582zEDTePP5Ms8kj7YbbXCKbJdFFeRacMM21CFgMPiPq
+iecVNgd4TaSYxw7jaaRsK51G44Lo17x7ILqAiQ4tgiuybGcZehqLCwezkvsjEhd
e/b+emlE45MoGTXxCnuZcdJoVivkwuWvc2ZzIzc3M3aK0rOSC8K/Bns02KjHjnno
w7GcZh0G64Nog8eFVnozwZY3NSjKZrsTKiRJDt4CLgizHzTN3eCQUGA+tzsp6vhD
rpECEa2A4ogKVI3YKQ7BGwEhRygfQaCOszHDvXW3isGaKMb+sWHLRTTnO0ly0iKb
yf8UR7qw/xy4n38KT955iJdgk/iKOn4+P+NFhrs6DZ4p7fdCaZtQCmZkGqSuBk9X
gkWRKm/GdifNEYGNkeISdAX8QAzfdJSk6DDxsIB24owVn5IqNQSGoqaiyPBvirIj
NBYrjKkUuPg3rk9iSiqiNKQrfZtpQVvVqrd1LBYUIMfX906/TogTQXrqLOAJL/qK
s12RIQhf50QSUjcjjrw4E9ghsCbq2Iz9paIuxtCWISdIJe7RSLCjHurU3CDYsO7c
LP/kMGUXir08LauJaFMP+XWYFv2U2JkfkbzaOIsO2RExkdiCzM01K1tEQga0+e+D
KUbvQ2Puolb6onUEBeiNa3Ad6P8WQoUBBdnBieDA0KzVnarEIiPbJG88EjzerCk1
yZEHJHIMr03wptaEKn+wd4goYrJCm153liAJkA8P7VLHXYkYlV5JAodFEFpwqcGG
RxaYGKzuhEVxUVOM853/T8yXzA7V/0B5Ju6/2GaYmmzov6UPyC4bSBjIh7f5lu9T
4wWjTLAsQzaR1OiyTHiCfN8e/JFdW1VUcP5AbEErVVbvrHh1kpIYOjMgHYgVwE+l
7tpotw27Aaap2XUCiSm3pKCxANg0qO5/AGdHcquJ1nTo6hKhiWo3uUZspICEgvvW
TtaU4eodyDeF0AeQXZbEi7bchCHHg2nnzIZXA2c64JrDA108lrLez/TMb+8w0Xg4
16hXvQ0+gN+YYw0b2DfTuyMISnjAXy29tq2OF+4Q2Rq4IXKSi8gKIB4MNTbNcMA+
CsiDz/AOKG25ywfkP6h2mmRaLrMVxT3IchQLUIL3v8okBZF75CwhH0e9tM5W6kEB
Hz3LWbNCwI8vNn4TNo52tJcBTsLfCj8uk9DF1b4RC7M888bLpPBA2fcPc0L4C6b8
hCRHVpzBQXhrKyTsYQsdl+fDmiUd3Bd7QgG1eGsu0gpTMO5NPfsJT4pqVROemI9h
dNnoJ1B6gNMd691tXtDOYb1eJpFDVj/H+6BEoLkeKhm5cLhm9etNhcibwxeu7Rfc
3xBo4DwROkZ5Gl4JKVvd6mosYbs4tTSwK897dQP+MQvUlwhN6ncQbqFQ933ffFyp
jUkwku0K/VkjwqL8DD2AMcybMvvriyyM62EVZo3nYNxEdcUQuODHE8K3znri9vzg
t/Fh50mXqEuv/gMGVq1hmmC1Wg77T9N/YG7Yrq9al1l3x6615wZenbB4GteQuAcM
7lWtOfH1qtwPX+odUshQ/7j2lvE2dRXmAMVx2rYwok70dtKZ4qvR/K3FS2JhQTUE
ySWJtm20RIRnzzjf+gR6EDBZTtVLWmtuj6GQgXSOqY2jCAkIx4keDD0a1RTrD7Sq
xtmYx4Ec1JpUdXToQZTVf957DDQNW/nIOFf9jlE6rEzEWfXzzXlqw9ztGGgd7x6c
Ca8CvBDg939S7FOCD5kjl5atJlVGWOnsCiGl3QU/YzcCiVUded5hH9yYfFF/uTY9
F4nnPEfQBRo4weYlAgBdydsQoYGF5ACmuk8/6QE416C9iGKqkIG1tQBOTm+1LxsT
kRtkqC/PjspWENKi40kH5w==
`protect END_PROTECTED
