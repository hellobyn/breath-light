`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PRgqPg7XqkBGjJ8rvHjzNLfbIv1haM9uXRP7vFdOzhzHQJQnCeCgBynUC4pfK2M0
1Ew4WJ4x9U8gmCXh9WOPjQQtB1rOuzSpMFM76NZjVn9G2ddLUdikg1wqat/hyqy8
xW7/g9xiX9tMyyY4vnDtrH7mpSZPsvqMTDhSgtwnxiVDw26+6zOAB9tmBZq091/z
RMLdbCU/fTfu5dJIBo51qm4Va3qoMG1Q/BSGuiX10Jnq/zaGyLWr/bsdNt98mMNc
Dzfp0tDP/LK7lPMTwpjlDg4j49cpwuDuagFq+d4pRCPWBrsGMGWqH4t5a1OrluEe
Vc6B+F1Hsie1g4EYMFfgGB1cxOgYq9GBJF5jv7qu7TbUsh1zSyIH+TO33fcMT+03
8L1sUxGrgJc/VnQMIJi9b2SUvGdMfruT60BaUUyZxDEqgyPhkFltCZvvSSd7QHK8
zecDQM8axzB2FqdisOVZcYgB6eY5GiIN5XhXEF9Jrp3Veu06nRCUYXBY3aPLmkXI
PjBPcG1JQmPWXpxxQxlfs2Olf4Va46pok0yY17/ds55X9N9As7b29lvt7BVwv/qY
UVS4jR3PBcTx1QQG1CGIEb02vboL3Q4M+LDzqxj4DYCxQCIEVR/n0o3Ef0LCm+K3
81UNpMfE84lSiYOr/elVTGFRFu2XZ2gHZbKHhf5om9PMT1/HeBRmg+9spDEHji4+
zKrqK3AI4rb1knO8Nuz4mIPT2eNSQ1OH7qgD6LbMM/f5WngQNNPmXcLyFugfk47z
5R7nkYOunODmChXdS3He/3NthZCqyBe5gxJllcC+/XiMgERDY9c4bvD4ME3bEP+T
eaNEo5dEx55OyRH0rPGQ9QJ7GbaybaeLk+4ELDCfkhFBPZAP+Q9dXeJkXDSI7aPx
43Cd1j7wXjrCD6+0PyUB8j6FFybbwcHHp9pu3PFUfqjJKEtZ1lKEY2cHTW9LW4MG
M7s5ba2uNT2DYuMPWeXgTyZ2/W+mCa4EHMjSo/tn5vk5ygqjvxq0wpmNPi9mapKf
Zo1dwL1qYqPbAn8cHO4NAEqF4/toMN5F9RJTOVYmJVfMgHxlDOqcYgzxi8r7bd0C
H/jbRC4Ol8/QXdHuu3Rhc0I5x6k7eVSNk+C2G/5tNDv8fLit/UUBLjcrruDxWqM2
e6CnW3W4sSkEZlM2lZEconHg4CdjObafQDCElYKyEIjBt01UWu2aAbm8m9z9BDxG
jXvKRaVWDTTQ7HdPXM9TFDI8poAmrfMLOmGxl8a2jvhqRNFWoTdMeP5BHKmvkjAg
LHIOK/9FLsWdMLu8umCpsEdpXkDnjpIWBZUhjrhQV7q4/3Sx3Zz1JXuieU1xDNkO
gQwML7aV+em++8OcTiszaZCwQvWWsuX7x2dbvAzlYBKViDEqB3m1pt0z9zfpQ4do
I2LCVp0L+XufyUsxpVSksO1eJfLyDMO9pcmpCq2mwYo9ySCcDXXN3IecrqKQpfCW
mR6ka12pP4k0HbF63ulj/hV9smfW/ksxlTwVh4m+aIjtLruDRp2GIWUo2+VRZ0ro
zIbU8ZeqdF02jPmfN8GjEWO08pklnlyVINcPMiO8B/a0WBpA/WzoYAMB1YXdef7Z
YeM83ChRen6cSWa4SD8ss2OhpGZ0y2gOwQAVd236aq1EG6O19mCvyKjnhHKASK9x
DwBtjBzAx0HOTSIW597xHc9oAzUtINJ9CIH8WzyHiRPocqKOzBbdwrxAK8Q8TjXf
xuTSnNIyw5P0gTXdXqskMZgP3pQZ8c7DXyfrzF5JHRBLJaYz56zI1/9vW5IgVNhS
TyZBStrhZcMYmUZWdujHf5euGvcpOPjE+4zrDi1soQ0J/W5dKbsWKNdGYMkg6E4x
EbqCwriiwEfPkT6RpeLCC4TXBdKUJJKpxvAfbaUyfaata6qRCV498z/EFnlx1upi
wPI1cIeTw6Of7h4B/CVSJeQ0DJbqlfIp3Py+y7lokEcdxVmft4Ab11hDmbEYVBX3
OUtGHvm2FfR3c2XjFWmegF2ozgtJ/QY8x76lhMTBNrqjc1SJpl7Pmj2Uqg5BVBOb
PxBtQcgG4EQ+zuPacUqBoEcQs//NGWJRwdxmxGeXDwStlUvGu9FM+Jf/gETQmXD4
3IyjU/n783gStbd5gKyQfZqtCfodL1vCe2Qu/H2O5I1msychHXT3zWAlvSQ/TFn2
r7L+M+piJrYAP0DPJjLqlsLZwuRKyZREFr+MXuN+WmXoIYpytEhSBUIFmDKcjeZg
ZHzJl56MfqR8gYLroJaek9vnLGG5Nftx5HxVvPP1Z7WdScvnvyHEKWzlv03r/ta4
G+IE5vEWbGuyyzefbUlCBWcx1fyA+DrGUyfh3OgS+egotVW5uQlY55QNV0uERaXv
lLNXBKLZ/2fBL2JCN4+8hT1SfYmjoPIAkJp2FeSNVV0wLl1K3a4AK4/2HANvPGem
HM4l4rsm7xO4nSA/JavQSUlaEtYwjH1cUkFLh/rP0dkIUX6SIjsMTW6FnM1Y4091
M9jSXWIBBP2khVqPJoKNk5M/VDbhEARedMD8a0nl1ursEPJI31A92x9FPfZtPvRf
2TuE42aN3wv4qHk9GrpoE1KgbOg5JSQA0v3S6vwphC56iW2V9YCIgwiSU7RCYCkK
W05UeZ6CT5Cwrx1NCiEMCncS+AdXUotQGl/alB4dBq5EY63c7mELjIjz33R2htNP
Xy58jylrUoOidb3Mnv8EzXWHH+0xqgc6x4gbyz78LZs3kHS9IrRwIp3veu5Md7y0
b0xkKtrox1TpOxfjYALMxXeMhEJZNXc39J7+Sl88g/3sw88O8s3YCMmFICIcQMJM
PgAmFuLSxWWMk6F7a2KKZLOLkoQbiVrFxpjnrtyRYoM5a+aBsW3o1naAik8B2w3o
MjvGioxGmNBTDLAHXwHT5EFAkXlq03eiu/E3J/4xZUoaQMITaMZLJsa9fmEuUq5p
Bo7O5L2jXR0G6qOR5Ghs4wh40E7lrD3M25tXLQmDMzrIJ8h5rg7oj/usMetAh08V
eqqfcBX8J8MxSZT5cx74XfP176BsS3+kbJxkfaeCjW9PMHzZzt+Yi0IX4tuFhH/b
vpZRNxyQo1iXsf326mkk5lqhyxngwn1xULJZIyEeLbD1qKdzJQfVHFVuHKW7VITl
FlOlVhrPNCAffksXHKih0T7RkLaEF3WeGQZCmnicEqoGQmMXrsQDc45FlZcwQBkr
efzM+6Q2o9Xuc5ZU4Sbvauh3uKXTGSgATodJ5fEX6+rutflrhpVOt82p/2cP9Wla
XdvsNGGv4L/wbmC2vg/MjTB1CgfMsrmGwEAxdw8s94LQbHSZ2iDjHfaE8RVZ00U+
sZLdEGcS4Atn+3sfmu9mzvzzzL8k1YSg1pZ6n7F8IMKUrd2Z2n4mwVgnzdH3mG3P
rTARRgOU5HFT6yY9+mupgZNnGzdnr+uOIcIcugL1M+w81MOYxItay34LjtiP88LT
1Xk3SOt46pW5NOE51TyhOSkM+ikE1aEuBBMrR+beOixJVp3WOxIisenjDpXaf+Ta
M0bnAKLgbfzbwF3+TWSAOft+pFKrK8q780vQbWroifAMRuLTwih7YHQLlFaic2zP
7BmsRqCXIoIrPUTobR+LbhEclhRevsM0hT5gWPiXGbsgYpQuf7uZkTTDSsodwoIa
V7w+VsAiOVi+a6U4VWjdNPzzP0UXf1WaZr9ZQbjM8H+6o4fCgGhMgLR5iauW+P1j
23/Py/DZipBHoD8WuZWVLIKo/a1oFxhE2vSS4Ywh/cwrd3UTjdf1GmYkrH6hhNgs
61ptZx9u85HBqcnBmTLHWKSFl0ZYueBqS42L5n7Ji3mpit501l6zBgE5HBxxEdK/
uNl2c+m4aoa26xfmpMs8DFKa8vb+yK7eIElov8B1+0VK5ae+SljuzLNYoH18zfdr
znoS/KvhdhuHTYoG7WfxvVTWHn4agSsr07muzoA4qVvS7jGg9WZUbCJDeUXP5Qcx
MPx7llnAyhPa22fNctqAJjO7giQYY1ghvN7ZjDlWyJDmMySBsTGrAkNWTU25jjrB
RT87itPYlhogkdlbZe5tXmnW6WGM2u0IpJIlKNZfmmH/MUXf8dN+HB+i5IMgPzWP
NtvVCgYeCotCZEqEUF6KOAEUkuDYT9onAT7hF3YDRRAKsB/tD0gyjWBNHHWFP3YY
boM9Dp+2ufOkMWqvy20nppgC1EUSkKYaQEj5BQz8yNRk7YPWGhju3MHNWDC908pS
4HSbMFsFOc5GbnC+FPbO1znCkch7S9a0rnxxJTBh1ld5uzzVp0y5Ut5cYxdVA9UF
wVXXCsS0x2dWuT1G5MvrGHiAZMjf5oRiRJ+PYn6g7O4FGsXnCcfdYtAscGKzIW/t
QmgFU92cHj21iNjP8i1d9jr8fC6nv7ApeHC2MDuco6vaoudOIvajoLUfz+CC/+by
A17Tep9WkhogmOmfaRxD9dUWoEy/cevzYQtSjczJ2QG2QvmtjDTbGYyWl0TXPqR9
X5rWZ5/2cROtp+RcmB7ZwJ9fypJER4Gu3+dPrRAb/Z3mHoqD8efU9BPeGzPlYM5x
ZPPIjjiyZ4nqtoDrZncxADJ9eHui8ntZwFppAC4wDAC2AluhSmbkjieyaoR9aTB4
oeLwXVk7Gt7PFG97bQBt/MQRp7+JDDlwjf0/sVx4O4Gt0ismfWF5IeJoE6/VAkl6
rrQm9BTiSDJxtflddRJMEO5j+3XuxnegGVGSMQVyU6Hpmj0iGYYlTLkxJmzTjxy6
tV9IBt8zBKtnXjXQzmvuwY3OuWMW+WVG7cnX4PzF+ki6y78mfz1Ciwl1Hn5VtA7j
fDrLHpxelVeKYBp1d9O1OrYL/UMPwdLEYKMIdny5mMSZQsZtqWKg8D1DlF+OZ6/h
1euama4mIO2fb0vSk+ESbC+6XXwKYV6+hrYtFDufq/xmPZD956EIzFsVXwbm71KI
8jUt7m9NXo0Jlyostc4kRN76tu3cwHBtTNE/S+ld4TIIxfznsC7basxCi2V8xGPK
OLtIN8sYYVNd7di7vf9U713l3Tk2FKa9uzoGWVMGHdZ1FjGe/WEawZATuly4Oq4n
2r0+7tzamVw+NI5MGSqRS3QGIrnXeOdCLNk9kRuLZXqyc5R+bA8z9Tp+CXaAuoOw
SGJfGr9C6gQId+OqRYPnWr8P2yzwCZ6JvWSMzHx7jEgTcbWD0cgLDoJzGT50HLNO
HLUlUQclKtlOCfHZKYmNIw0BK90Y/XofpGDr95AEa6rPtwG5hCf1luVXjqSs0XnX
kIxMgaV6dymNUDif8yZPFVrai2OZYiEXkmE9KYGAVGBC/ILEyLB0MhUZgcyVTHlT
JnWtATRwO6KtXB9UG7X0CzSIW9eCsM8cjdDusHvcsCzUGQG9cESTLcESaGOFQS/7
rQBLHRo0zxd70HkztrItil0KRUYIlS6TBCpf5J1BaTGqPv+HrE/CokwyGkEu+lMM
yMMtTZ1eID3SPhtzhq781htnXgo19uaAcwGcprjEvPnLNAIU0C30JVwXB1OhuSSJ
uOuqDEiIyUY2DL40h9yRA3fy6aTgaKM37sTAlbv111SzzBEXniaPofRsTrOQltGg
ULEN6KxRGydrQlf+1/qOybDYYyPZSlZ5JvoVlidRf1bA9GxTid+f5nH5yukw5u6C
L0zjlYLQOFThAfAW2E3VPQ==
`protect END_PROTECTED
