`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m27iVr+Y87OwvPFOWADDZgX9M68/oi4blmtMLNW2C5dOL9RfpOJ+rN9J6KnWHQO8
aj5vdP2J5FII2z+f7LttmmS7GD0IY1fARvaqZHBnHL4ddUB4hjdmegHo59aDKHpT
um0OfAiOLyGXrGb0+/IzdoEb8PRmSbUKoHnqItIg79M6FUlI71zQNjxvf0B5mj58
ULRKlVptp3v7yZGVTrLEkM6vMYyWJELMkLhfoLg+Zoz5xOFeF48XpEBij2F7gauP
Xq1uPrsFkWJlrRPxwZfe7IL+Nf/oPbmhwBZRId9ewWYQFM5QirRIFtsBe5EfD+j0
31qMo2BKrrSmt0ME3zdjrhtlkpUZYViUx/l8okWfGYzdPxoO9+XYi0/OH28p7ZhM
mQFdpkXF9CzQXqyX71mlyYLokUaG30xH1enBrwEhlfoSFTWWfJ9k0mwMvBLXPPbA
yd6/aQYQm+4gZZr70Vg+cutx0BC0TbtdHxH7SPYKJAVmhKGUjD6gUYmCDyb20T7K
1zO8666p9GK2XMd5vB4duUBe5RSfVlLemaW8B3htSQceK2i5S6KWtMjp3GgsFfTM
ZO9HDymQp2/EXhO0DmNcJDu/QakJjrBxtL47lALSm+LKuXtXbVf0wmCe8PEkTiKG
1CdmPD1+0AzmzwLfdqyq7Q3A776RIS7Qonam4N5gvqVVVUNUy9pMFU4ZM3i9S4w2
+vz1fzxR8/k/moxrwlker8qMrZMV9P9U22quj3dFwuOYQu8glkgc+UnTlORKt529
srAI6HW52pQ8hjCn9uqQb9a/jcouPRs73uTCK24ZgS3xtFcNDbB9a7Ogw1BYT5b0
nNn8oaSJDxWfVYBpTkcsppDcgY0jEVJdwu6zwQHO7iWDcrfm04SB4W0/lnM1nkl9
CgxYYCBA+v0hQGuS1NXhE+f1GuDyMII+xrvPdoXYJuCJh6FhZvN1VvFJdV6sn+A1
G7Km4/BsgcoAHJcikTBFtOBVL8NmAUp/FHBSwojv9IM323pyAAvonZKm91feXTv8
CPSU50lQH6j9ZasfaUrYFBOPhytD4OWFnPv4JR8WdQ/Z9qdmWc3ofFn2XNlYbiIf
zoA/QAorPe51JT9GAzrOOFbBztW7kBVKwmW1/1U6FZj76tcYBra3mZu0deG6XQaf
EDBz7D+Lc3kNcgVrYDgwyM7JvxLTeiak8amJntd3f5bQhQ7sjKVU/Yh170nK7/ow
TIJIY0TMbSEy52r268GrLIV1R3BAL4C0bnXodpdChe/xtAcuRIktccZNhfHOY0+r
Ix/3A+UBrTS0ZCW06S+5FpBue6G6QhVxS5Y65qpZSiJ3V3l+TK65VpBWkGh97fjy
1jXNibrrb3w/Si0J/uOvAZ6zXTJMNoSXENZ+qK79PTu7LN1LqlY4TA45EmL8lGF6
6oQL+Vt80BpF866exHTPp9E+MfYw7z2wOWwzFndvkGF8vk15aLvF/4P+1t4x3M+u
piOy9g0i08ApPqHfZM4c2du7NOeie6ehRobFYI/InGFa/ec2jRfMQncKYFrBCPlN
9Dzzy3BMSjx4/WJlj0uJdcw0OkgcKL3n4FfuFqaGtl6ReBIv35aA7ISxEdbcgsT4
H6cdzVWqPtayLDmYiv5CMiuryrkU5o9EWScNdkR3qme99wM4oJzQbEdcvT+Dsb4i
vGM8FDW43tgg1JJjoW4w3U+a5W68y9lmj4vDQItasd/B6yVZwV/rHMQUeBgedIu7
uH71sQlFmxzaPDmvfhrzXYzmVZA0PNiNOgYQ0p75qDfjHAJ3w3a2lanHn5YRhQHr
RsRUvNi8TaJviMm0f1EL5gTIVkDcBGa2MRSXkTWtOCiyG6OrLyUt/hMS5ENM6Bpm
zEbkXxXkDZbLh1fzar3f0MiKNVUtvgVP0rEStBRuz8tAymGdo4W2sgNY1c0kog/4
`protect END_PROTECTED
