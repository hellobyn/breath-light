`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKnWJRyBCBrn66k9dnwCj+Yx0wfupP62wCIcENJ/DgQSMWJF0xKplJD9Ez+fJ2/F
YBvLmcHGGwWPfuMBN2R+e3tFD/Wkw3rfDmH8Y5Vw3DMigknNfIYKpVJJP207pRqu
BC4ucCNlaO7hQow3mZcJBPZhgGmmqY7TV1qrKl8qwTXg7xWFsk0fccQCd/fMMKCS
l/mQhbZkXBGixVOZugjQhnoivd/ch3VyZQeUBmdJ2vAAQeJExNJkRZGEVKkEyS3z
GAH2YR/J0ACjrYgdk7aKfX55A6cxQ2mTXMz8dIDDXxZ+6wY1pzc7N5RiDC04GMsh
5F8+kMGWSmpE37xMGHJe61+xPKWXN5Qb/cpuHaXcf/DGj+tqde/vEnUrqBOh9Rhx
Hwm74PqvaUn8SyLHTFEXs7I4VN8PTVyXZRTA/90W2EZO7fpLQLocuQWK2EMZPZgZ
WUsBhWrBbvPUP6M8XwOJ5c4/A54RIhkmuqgsySd0eaU5ju0nJkxC2oIyRjB7T8Up
IjQO8/sblk2LovXP2rEAIbuk94IIZZ+g1r+9X1Drq7q1EL53T9dTuBVLq/5k1Bi+
FLis+UnRH2CwDjPZt/ka3Q6U6MAXBlx04nfxYhvEa3zm95XqrZTGOuRzzUpV/3h0
AP1pdRg9fb7SFNi41mEzytMGymfuIOlMS/mk88MQ2E1oAMAytn0jwdlLDkqI4Zrd
MQoVBfmtA+PCJSwei6CZneDni+nuAxGhWGf1SGbMogznQndUoGrXHFVKPMxLWQhy
855CkIPvBvwCBnCQla1GrTxCMK+3wFtvyx8yy+UDaVgOxMi//VGrstdQpybgAQ2n
zSJQX3uE1k8aBwPC9GdZlroF5bdSCBBD5aInrR0xoJ0RluCtprNaKfusEYBM/nlU
nhCnR3JpaxutpBDvyQ9vlsuPU5S7Xk36gl7DUA94vGyYk7tASM07HKyq06XVVgsv
UmcPgnYGhDXxQcF4tNk3n0Re75kfjsLzI0LLrGlhDJvHlAkvJ472B/BV3ebUdEZw
1YO/e+/12FjOdt8+2b65ZdwjholKtS4l71pNoG+wLjjDK83tL9ORsuD7jDEwT7cG
mIf4QBRx+ODJ0I/JFtXxe8JhcEAbqDLPti5HO+hmn8cZzaL+uMPTyGDg0a1rbVy4
2cupK2dM2jjAGYkBmpJpRO1NsSTfaxW5o0ITzVWkzm57qLDGFeiIUEJd77H+K5+m
iWvA6efz7ZPM4+ddXIWcVhKL+mcdM0WJ3E9sxA3NKMLCcsEht+NDSZpMMkd7mnaZ
PdbvuzbOFHRBxtpCXdPr+xYkideibJzALVtrUNAwlvSQD2K1FTwXXqdfGHBi7HAQ
9htkdrUc2x4SdC7EFrqzithrnUIGlv4PQlmYg/t9c/W+8GqHLEfe1TxCKq9LBFcv
92GT69dFNQfr4oLccnex3b6WR5WtfbvcGZos/zCOdF84OAXjVlMcazx9F2OAwVNv
M+cUuH49qG0+g5ztWnnbUxrI5RK9sKIQWP8BDznLX5PRGUBEmGj6eLYutj6/kNIH
6SzZ3ED+bhsfCTTXItaJHQ==
`protect END_PROTECTED
