`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vk4VWxQPc1hM58g5qQX6Ns9HxV2zNnGXbBk/hqSB0keasuFat8f5odd6J+zfzwig
ITwiZ1+Cudgoa0sH5BkK2s3HjW0NZwiOa5zpSTBRlX7pz8EglzoAFuW7Xt5ouXVg
p91mrO9svMGA8ybe9g5AO6j9e+i5LP208eDBFys7oQyApMvL/SArhyJ4DIShTQRU
AZEXwijtD/Si8uGSIy+aN3o6ZfdaLHwFRW1EuodLYZXVuZNdoTOdsrtkftYR18nZ
avUhPPGPaGzT5DgZy6i5P3ulMmDqn15EYheOsHnVAsPn7rF9p9ftNyEB2xKzg6hA
/zOX3wr+17f+NUA1pGvPCzTu6hI5q55gLIsu/tUzFXNxS7xzX9FBo/Dtz4RysWCU
52OQXOXfcmUG46QyZMqPcKnr2H9/K5Nb7A0KbBedwR/kz/9JXVCEsr1vMeJ95dXT
iVvEDLlm17xTGlYnXwi58RziLEhgdmPh8NiUN4fmV6VjaxhWxBLkNW8ZlKY5Yjsi
wVCPHwjEwzUDPGMMeL7PhJ9Yr3CZ+DXRkCh9HGpbyvslkxhjxuTavMjqE0WxuhJH
zvbxMB++vlR5Mou7DhDm9PlxQOEFMU93q93rA2xmXxv7Ih9AYMejVMOdNyum+GcV
`protect END_PROTECTED
