`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+s8+swX3ShLksJtduQClmv6ytvygrm1bdZvuS9x8NU6tMK/mF/bDZ87e706TGBM
yEoHtJUfwe44Sx8T6ZcKYOuTT5u30wFLQOWnsUGyxqX2Ii3mxpIzFpfX5BJFGNg/
Xq5gNJts9fNXNCXsCObMBjFsVuGo6Eg17Lqk5LRTEkrAUqjZj6mInkDWxZ8V7Pht
2sKfE67Al8WfDZnSadOSiIjNHlmiSunNdT3rEvjUAkq5IlCm3d+gquQMgbrF+bsr
PDvL9DOs+wCfjbOOfU2+9aBJLXrJ/M67GxRIIpUGd4rwZYTvMA4vah0XCvQBlLHf
MN6Y6X/D31uCooAapsfeeXrkVPE9PexNa+81rIs8IIEHTaNAzHVQBKI3hjjOTZ3c
uXFscq8QX54AWwxqa3hMkF+J/deJ1dqlMnOquMO45/MKpg8C7vyqecz0pii9yYHq
nGiPHxQ1N+UhvjAKUzBKLlCkJLxLfhTepeq81pOV1EY=
`protect END_PROTECTED
