`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/s66WIEmHoen6clbuoE7R8mrubvkh2cUduT3dTlf+/MiemLYMYHmKETZmjiQ39l
QtVgzVuVU6m/TslhYS8GDU0w05c+GRuEwS5A5HyYctBsx2mNtIJKJZCiXemJHkqn
cXgQ7+mmwiL+0EgcrqOKx7FqjG5IdilgxetNTs7MH5qqCnL4gwjWI4t4GDTHPVXp
HvvJdpMt+thrChfTwhmqlpAgoBcIM9REbX0Rf2XRvX+I5l4JZksNXxmyuPJwTGJ+
YsM58bD8ocQ1F8E0Hc9o+TFVuET8+cDUgZ/Yyu++pEVSrrM+n1S+fcW0lPHbFxru
U49qOzOz8ztQOMKzLGrh3ecMxd28TQSuSoIV1KvsZKFDExGXmz/7b3cYnNXXLzK/
ZTvhJlFGYe5EphuHU6HpUMdGL6aHze3qXOH0t9cdhVRFAlsRMPBplTfwUwNUWCZ8
4jgo6iTAvPgkfLEnpN/qHikKGKGX+mG5jmIj/apicn7m5R6025q8KmWJKiIQTAU0
2pL3KCdiQo0xLVFNaj1TzKUcEJR1to16Q0F0VWCMRGdokXl7YLDAVKkdBL8m54A0
Gl7DwOtF1d5cxLBHVbqGMkwFcSw/nsjQbkEOOfNeDNDJbDT392pPNsiQsCtDUDPH
XnOssPogi3dc9bPBfwmz6HAV5O5FzzcELFfR2sRmcR0cLeCBuzC1TEPcu2urolGB
s5p0Qeq+RYLOaxJdqszUjHsKKUpa2oEN62PgYVblZgYIqkJ2OoIyP0tTxXpdoW8R
k8WRNWpZpX0PDdgszV/lihIRGPwGE2txhURQuHxBQ6rCodqnt8avFXK5aNSsl0FM
FxI8+G1zDC5CtEGvaAI2bArq0qnahl5xo+Oyuj8nboOHFghorsSc6/4Kf7W0fieU
xoFjhaAJF6ZdGeCePXeVmDY2Aie/vsFm94J6oZNA6TNStv1b0c3s2JhvRNcXHAO6
tu6gLTIoSksNGZs9CIDoO1us+q588Odt7Eop3NtXjycsmeyy413Bpj0BlFC+pVLt
in1XjKXnjr2q8Ef1NbMCUD9taaeCG0pd8VYmY0EIbsFJW8Np0tJ2+4zycZ7MfaHV
bXmfhcIDMv5Mgy10xB6j0tmNFO1IwgqfbKxRfKRhwQevw3BVQhbv7frM0r+bV9nQ
kSaJZIG0TjbDFvcyKY0MeJFilt4gsXQUVskYZ8TA9Ma0cX0HtufuY+XyNP/llqDo
QyShMTezdtuPtPxA7Jxw/qS8kAnMF98fEdJCe/o9arXk56GhG5hsZDSJdCvXDP+2
bIYtpj4b8qtrbq/MiGEDZTK0B6b/bSWF0AzRmXO+WbKwVX2SMQq4CLdjd1qap+RJ
6/odb8HmYqyMZl3Ur0q3bKmCzLSAcOr90791wAgyK4f44DGG7VZ8diT7FqJsrZIV
T++skTmnLMiuCueFUMfb7gZgwrnXrhvAShhsVyR4UssK7FIGLT5IIzl+z8QJAVPD
EoeTXr/ZVudWIX4TZ0tT4dgAVl4RdwKDnV/EigkV709sktMKTA2UGM7BL2gy07Jo
IycJGa67UFT50BxlzusZ5oVjpkXKSDmcqHUAe32nMzmW6FI1Lwl5qkUXOh7pniZd
hAaOWtgnHsHkxD6BRCDCoDARPR1Xxhm8f6EfZb4df5wh3WkYEyq+syQemjO+k9Bs
lKZX9Mh48BYHOiWbTNziMOZxT8qjdMGigZLHELk05pxleF/iiEQHrIxu4oe2v5zP
eWkCe7JlAyqboIjL/G0NNO+WGIwD0SBHKTKNKf3JVjP4lm1Fpbhvyu9ZAIL6oA4G
F4dXdyX4R1/1AjRD9dPSCGvjeLu1l5vuC8NBJbKGTO841Do8eInxv9NQ2tMZNsmI
zbhQjQWCHRgYZypkQPE0Og==
`protect END_PROTECTED
