`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGm/+rII7gJgjOcyJOSyK6q/68fDbvhEykqSuS47YkbvJ+MdxP+hpkKcKPiIEA0R
/tdG4YDbILDYMxfg+E0aubOI5qe3rIQUXXLgzq0nMRx4aK/36dW53JxESWnNCyRD
q9Hk2stzss0KIMC8+A2PKTImW4e7+cx2rbNhzkxnmwGob129egZKS2BovcdWR3S8
NJMOI7fZo/cZHjQstT/gGeDaHU+E+QpQuTh0cNzdH4Vuic9WQtL0O2isLZiwhqpO
if9uyAUIFqwSaMYn/aonoYoovmUzFKSDPzHVbJ2KnD56Vc7S09kePaH1AwaY8gQs
UcNSGg54O3SSqWHtXm3CLG4IDybqr1fdF26U5Un9LEQejuR2kwJmu3bK7yG7pL/p
EGOfApdPiHyo04Fhu7zympSqU78r49TYUOcm6pkLTYH3nDaF4zYtj7Idc51oKOCA
l0FHQT3BaDOo0ltMUETvNvLN9gzuGhJ/2Q95bUpLi/D3AFKBvR0aiHhvvvBCjIYC
+5HPzcHgtH0/vFPUMNhCwxcudikZWOTTHkDvlSk9EXHINj+Ob3Qt5POHRWlk5B6k
TB7/+wXPpeaM3c8WCvzZuW72M/fDN9Bzbbtx4zMyyAsapPFpQcqarDeI1RTdUb5F
O8EhrIkd+0Dim0Mpk3/WBhZcEJ9dXOv1PYSC4JJl6loHC3+u9Ais3sSKL+i6oL+F
S3FXA77jorrcIHFyNQGPbkZy3vPOxMbe5TvWRdgy4rmNZQELnbUsUetOz3HIRL+N
ht3StL6mqz63OaO+UYcNRgWSDMVo1RteL47VU3eOOXU=
`protect END_PROTECTED
