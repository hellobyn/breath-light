`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zf6MzM0qiHR0H73MMA7YmfyLrFoaONDgRjvVCVo15TWKkhhPuTA31VfrU0peXc3I
iIPEOedR1VjKN7hYZpzxeK7CNV2iRRedXOIkRv6K6gqDsJsxzbiwmUoctt+o3j3C
DlCENUajuXbGCZXqFfdQj2N7fO2sBnc32tiDJ604opG1DZX98z8oiggVbTrLwha7
67Ap2ahqdNglZjMgbCCSl6UBDhbnObs2dvRbeaXd9+9cVSX1akkDMgqkn1hgMfpA
XRsAdGyHKvD0ZV8+6kc2dnSq5/tMWAW6a5gdonrsbc6/9i4noIZLd8G5OlForZ0D
MdfeBZ13/EBnjZP63w1qD94e66GW1GYiazawcn9yUeGpjyMSOQ30931IgdkRYDMX
ntbJGfqBWFFnCQ3JPHegTRSlzKZDQrDJMUD6XcN/2fK5BFH+H0aSH5krzeR9broI
cfcPMT5NFR+iejzaz989O3hmqaiS9mLGKUU94JJk/UqbXlnu9EuY3M9zkMNIn01K
EZkCEzpreqrsWsLfBaNsNA71knv/B7IOXKM+i5auUrAn5Fofr5O+0F9KbRDQ9VMS
kl3AA8gKngTRwI7e2QcwhoqhGwwDbjjHfI73vGt8taS/C9oBRT6oGUakWLsiM/p+
N0DCdh3n0dAprB280qI1CEicqliIHSfDxAmiTTlPK6CxIsYCad0EzLPnnTe6gX5m
YrkAzr0Lljb9RAy6xWf0sq/C0JhGzCwV+iQN3mP6soM0HZWL150nBPnlbAaeaTsX
OlqSqSYIwYbgP3qc16TDOPymBfNnkbnYZvSW1xWcIVEdxZ1JHX3xglPiNvALeLFX
iyKui7ImXicPshouHrPLcts9YEqUr8KKqqLZOIt3hUKOnAojfVcvMyquhOjNQ8fl
QebAIKY6T6zjXgkd0vffpBsbgQACcgv1OzFi9nbagDKHjY966ovQ9fEdk48ASoys
CnMo864buBdUYFmdbR6PU8wpi+T2ztSGqD9rpIyrFthsfrQDZ6ziqwvQZ00OtgFU
MZIT+pHdn0TxSbhZ3HODOMm2s8qqAU6+vxhP/XaI9mOHSSnyrCoQHWTB2GMjfSUw
qIQxFND8bd0kEvCAxQy1daXoSxn4nJ18mXcGaofKh0xT3YEtsVddgvdVdhtAm/kR
Rve87QKOMc6Z9YSqar/vweVY6cRti07QeX70q1BMF7iLg1J7Zs1cCh3dbkU7cnak
7IWN7keLeh7Q0SX/Oi5fYMd8HmAHh4rjNdhAy64Z0xgrwOk3n/gWmzDyAeQ7S4NA
jXDPjqsbikjwddPhsfCx4ZkwaOrx9vnP92Sm1MC805+nd5+e5g6nodyrMdRI1zGe
PqADzC44D6hEcXoRMR6/wMWuGKalSRHlZud/+Byz3zRo7A4w8N8Y6LHBfK6kUHEZ
aSCUnDfQRwrYS+bItFI1ZEJNB101sWytnfpltFUb1XKJPNxTQumY89/ZGxAXOaJL
8LxWa6gUvXmy0XLxSkZ7ayG94iEjhKnHtC9djeS/A9yFhqpkyHh5dUKOM3rTHtuL
KchKfyQLwvZjwhRtY79t8AMI9sqhTQ8Sq76B7ZbFd1qf3KtrfBJ/JxmREYTQ66zc
KXEIp0HRSEgbQR2LjQJlIA2DsdLoOKYxszk1vFHOTK+OZSrSGpT3thI/P0lqT4A1
GkN74SG63j+2VWqVHVVgr8Pq1VQ8KFu26+Hjks15AdKc9e2lO1Fr5XstChCXV9Gl
xWxBfS9NvcqrvAkfdez6yM+Klo29FfkZ06viawhn0BsqWVJ7Vboh6SGMGQP44FO5
GYMHJz4yWQgyY+gpOBAADs55fDGCtt+Pj4ftLpSRqZoE61CwFJ8UeeSRbbbXJqCX
Lsbzn8Kw1s8KlMelNTb8hzYskfAJSHBbf6FLWZvKYNiOQx4whVjhhhz9g2T3qBZS
AmpE9BnyHaUrUo54EYGODk2Z2sPlKAByodH1uMWtzes5TgAk/ZejXUV5MLuF/Xha
mYmTUG2t2G479yw5juwnfA==
`protect END_PROTECTED
