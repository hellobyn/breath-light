`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u9WweL3svFLdTYsLzDWEhq2ZqkX+z9GmTmKoenN2hS7716R9wsIRHTWtTyb0zCEL
yWyT1K9hP+CuwWsRcLi5a9VitBqmYGlT/plHxQxJldjttOCtNC5++qjy2lL3cEKG
RUFtRHjq4eufVdNncL3DGNsmbh439jc9L+Wc2y0I6HWTBU0X6rJ1QrF74iaMWcDa
kY+Btb49LcBv3ecqKkcxb8N6mSdxJmnHzA0AcyMqXnvxCOXFsd55jiHd/7WSZjAQ
Fl2y41WHQQjghNkrtCOTBxIrf2CkBj7/WEj8VDDUdlwIDqiokyO30vTZs1BwL9fL
e/CDTVJ+qWFtamhOW+t4Nt4ASNpG3rrEuZJ3XSI3A225BA8kH9EFNCOU8aWcgYCE
phy/llekox38tMajquIUlltKoKmk6/+9oU+hGMl1wLw7MtI1t48UaV2JnqKuOOIm
UzBAEFEmf7bsKmVLS2UHC2hFbKEjriWWB385D0WIOKc8zBi3LStJA4n8+gF8pw73
5KUu/WrfOVlEZru/AkZzuaGEfjyuF6k1Yhu8AB7i0AHBZRrLCf3Re2wSCRYlRtip
IDqQ+cjqFiWRO8Tn6b6iXGy11vfqnSiF3hfJ/SnwuQCxYllNvCO5ZleTK0BeR8H7
vSOeIpcWu4ASW3VlLLHQMqy14+jCuGxWVAya3DzuIf9RCH6MjYzz4fB6IhnnVGbq
xys66d5nH5LWNktSZW25rNOy6FdWfky0oQR2rw8+E4BrZNmbQhB+a640sDpSrcs6
t86dXuyxx3FCGG05Bli3K3tMRHZq2tq5EkKVHVmj0nIaHFXYQzXomFUcgLooAdzi
lbi8jbL92xxQb+Fewub0kwpoN5uXKhYEN+vbJK85/kT4ClMdw5r7xvIevW51bfDt
lTf+lafoY42XJc+FvYdPqq4wsSTlA9nx/I+no97+FkJ8GQMU7WA48j1vdd7UKeFY
jbWIrSDiY5OEAahhQZUCKCeJZcehd3OAwEYUdtiVAFqURGiaHPc5jFycvcSP2N1A
96ScNopiu10zsZvQ538n+2bhnXO8hNtUt0jyHPwPoFJZwBOolH3vdvze9rGngine
Vg1ExGSiYrtwd3Zzf2BTqUb/end8ee10zbM3upwUkhI7Srlvicf+75S6UHpSciaB
3OUEV2QpzOUJ116joI9qmTVz6OPZpAHJAewGwGUj6XW4V1qzQdiBadO+0597YOss
x3pe37pLhbA2npr0zHhaO3gYSeg9vKij4+tk1B/LMphcemnexpxnVRckH4KnUShf
AYNGIIMBxFWrgc6iNhtoZbZu7bHpAfHg1A0AAdad6ZPpyl6/ZO6dIT55Ro1Kdo8G
QDNBQehxpVo6zBk+bfsY+eZ1lyutyOWgwTVkBVgPefAp8r+fw+xysQBqI+Jo8seP
/WyOBXaIpJ/Catvu5D2CxnNfqRyCsCU1aZ4asHjSBScFIA1KRNzWscRZNMalLkEF
sd0mZkRI2rrnspQnJV746I/VL9XP8ttuB58XHCvvHVzXiEHeM8P4Egsfrb/pP7j1
RSLTAXnpC4ZhnNg4X07LAHEZGyHBD7IjyCE8iuMJRUoQUX2ngasWWOwaFUyw5jgb
4M7mhPKacF5NBn9pmp95MpOtl8hc+LPOzwDmIS0tht7BpxQ3qmF+Fj9wq5EJHlIu
L937+rfnjaO+JWMLxbEgHyu5RV9JE2a1gkTqEl093WNnkFH/gZyAJwPGNAxgDqMZ
GvbP/KMkACe/kF3HVshRCC6uUuSPqSykPL4axMm/9HlzLuxCdJ229fwZoU0JnHEf
LUupf82/FzImutOYssZAE6gcfSqUgsH7uzf3bXVJAS0BHf8eQG3lnZlHQke2VFsD
iHvhHcyUrQSc7V34dd8SwY3KbC/RSUh1Zg8kzzg2x+xzdFC3Sj68ggOmxRE3P9Di
GHfIMZig5Bhaqzb0il8aGE9gvkFp5HpsGyBUD5Le0Z2q/XJI16G60Y9ZOkgdOtKp
ac7ZcmpD+ktFq0fvgOdLOVCIpPr6j4Ws5GIeffm30cefBSRdwrT9c4R6pr7Qb8Qa
aa1KYcZqOoRXfJ10dhc7nBtjSqTBOd2jK1sZsvSbeklhHrCm3pBZscqs6T5KJf0K
YIi5WzL6VqJ/s4Uweu4hqMKUzNDWyIxzGt4nTTCP6drThQqq7/2mdis1l8iUSJ0Z
v4u257IlGOAsxoIdqKJWioK1mFOXV38NCIJY3/KZK0xnu+6IWnmnYApQvDSdyVAl
OBJxG2skZscG082j5GKCCq3Zi//3r6KNQW986KUQUI7mE4mLIPwC848wjcsFg/FR
0gFcbLBeGtFV8n+tElt90bpcLlJM12ECwHsvlF9M1lpo1aW/49QU4UlyJilyQW12
XLPWLIz4OXUi2M5K/Ek9I07JHcgKu9N4YGtZE0r8EcVwztpzpNBHp6zuMrq0sUCf
xad7jhA/9wOxQ5QO2h+/VhSxXvr66xgLbQXqmm4qiUseNEWbNQmde2C4s61gNSer
4+y77+ssyHZqwin4OzBHj5Jk9FVcW6byewPCktRxUuwwITVE3sXNEKmKEe/YNXR+
++SRiTdUTAWlPdwYdfmOvTbNuhk8n4WdG9WiNWzirawOwem6/uxdXCWIUiEXVhpR
7ietdhBQx7IaCOELZuBaAraG5Sqc0+4AG9gfWtSoV5c/AypsrfTHFy3AOC1WwgmJ
OCsu6SzE/uMz8f40NJ1io5kqT2+EUFhQB/cOQxqu0Jw2f8LGfbqg74QyRXiU6NS8
We+ddUx7YXUiGcLO2dCXVGv3u06dhQPGg/JGGTfT5qh+jh7drS2KYixve9T/AJf4
t9ADalCVs+S8bm3l+w5WAzh0nhpH563HfxMqK5PzpXGf08DzoVKil9KQ3HDOYqO+
kYyohTYEkqBcq8bqgggkAHg4zAayckvFDBGq5R+9pFp7Pq0lfnopxAi+7THRdCOs
sjZdscza0hrnNhvsNa89jgieXiCOqj6oPWdmCYQsdBaKkWBjCGlO0u3Q2KHp1L49
ep8iA9rhwUkVU5i+Z8YfCFPHEmfGGax6R2QtlD/F1XR/E6hTjbu2Du6/nw/1NxM3
tARN1AUX5LMySf8cCbYuXnV1inM6Z5jq1wyBUN1GbyiBTafyAVBo48OVgFMXKVl2
2khqq7bGpW/x2J1AMsgrMtjZcweduJdvbfrOHwHaO98pzjYswkxoFjy1e5Sp9nRS
p5dyU+bjigkP+QC+ikhCPQ==
`protect END_PROTECTED
