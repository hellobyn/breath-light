`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GPcg4KJ9vOaHioJxMiH7huevTZZ2uE60oxIFi3J5ZkprfcQxZOvBAQR9EuyRGKPs
sBW3Mb+PZNTJbY4uxIYyRf3SbDm/UyTcoW18jgs6f49LBxZEcJ5adzPO5a9+V23b
84o6nZZ9z/K+4MV/WBmiRvfJAF+MB3VbtoFonI4F/2wwaBtkqV0SzTaJ8nduxFEl
/5HHrIVlSPLRG2jcawPXEhhR6CSfALSyn0RPTbxhpkv6u4IYUF+1TyU6iS6YTY1L
TfHUvcgaCKXNuuQgWtdvfHAjt0NBWl6t+r1mflRkmnyoxf3O2uCmElGM7bF/A+mu
mwc74Usz9A0gVY2jcNcZ/ZRv9KUlf14fGqUQf+3PVeipa+zHpEBvExhuIQ7uRw7w
x/xn2Bbh570U+NG9tfSLlMcCk5iA6PC8H8ESc5+P/ZPezwiaCXJbL6p9eqp/sxTz
0+QfWRe5FF78Elp7AbDGsAHQWeZD4ZOcRHqic6p03BecHwCgDMQh6maeohs/JhIR
TxX0Pa1GejaL7Ig0e9l82aj3rz+vN3LDjV5siOQHQ+GDZizaOKAqBDkWKJV7heeq
Yl8zzmebEEsTplQizmJsilkaSU4fVe35uts/CMrY5ZFnefH+lcpujDKv+UEPKSey
ZbL8KzFDIw1COGt0rMi0ojo9YyC4a7tX++nf6KqP9hB3yK5mFhV6rpfsjoYu9L57
IFgyb+2G5F/PEpHecizi7zNtTOxwV2E2zGBtE1oDL8jldj1tWfz/R0q7hLkpsH/N
HQb7NSBkHYW4jbbHNqiRa8gH4UZl6nENV7GJIrLmr1FmyBbXhX10RoQIl+Gk4e+c
YvfUHWskF1sGCv2DfMDtsMP7ln6fKo4Yndhf7ma0TSKRnGBhoosHVGXDTmLJtGB3
GZkKB/jr8akqEO5Yp/LEpZjxWI6D6tPzvM/+NLqhdRwxoCTjYkIpUqA6iovmUQB8
S7WXDjmjvM+zlqsG3E3LY7zx+EbhaY5SgMXnh3Q+HKOnFxf7/Cu/J1aGxOCTUQpk
duEGiYUtSsI9/xBhvX11B9TU3tAtv5QnR8ifgvnS9CIjViw3DYFnn0v4fp4P8T+u
zCy9ZIGpA2m8JXGYGftYfJ2d9qDVaH+JdmGrfZUKDYAB9fEhcW5vdF+px7ROhhnP
K0SnsiuPcMFD2/XdrBrV+lhP4VHaTbOw4oX6/OWX6AqgjE0aWiqoteVM4QdOjbCt
inY1ZISam6y1bkHZsW6HnCgIcTV+lfTtzReUz+kmNpFuwajvop0i5aL82nEK5bMW
5VUHvnrNBF570zCqRots9lbV9VCXn4Ti51txOdvcU41wBweBaBWewqftDUBHHHts
sbYUy9ReOc2O0plHL63lZ52UJVTNtdGpdkj0G8KS2YzGRApEanrND2xBd9OnTyVW
6cyYuCsQq+mNSZ14TLR/ji8CCsdZn3GbBQ+NwjqCA4h2wnn1hcpD+eQtuSbwXVZM
x+3kvv0EhMjFFtTZV33UkKKOjUk5NVZ9xBYlnCGaVKl7c/jKKQMtvBGt8NIJPxnw
yqehuYOwTty/lKfQEsk+3NgagaqUxG1/j7t6JaYl23mqT29yntOx0FBmkr0+HSdD
7QVsE7AlccABo3NEJczGH4tCbGrZot2DJZpV/Azg9zAytFwSu6TrcwHVmxgl6V9k
qc2wwc0khWXUWL1UJlDoEao2M0c5yovzqISz6XS2Sp/UGP6ow7/uqzvuu0EV0Yh4
owsBIcHfz7PeCRWBjmI04TRXOGlIZjeC9ELSx3KhpEv7iuf7l5oB4liArTsTMvnx
7yvetQ2XXhxwc2ETaNtB10OzTZsalB76c17fZjALt00461ygabDy8ieqAHNXjJjO
lj4BeQMkoSlIasN1dPHQ4HUpiv9hOnGRI7kaf7UusT8m0rK4NIsqGyZcoudBiL7N
3nTYfA2WWdbugxJmojNoh1yuLJ+Tb2WAEmXK4hXygy8QO+HH6ZT3g7SpjkIsb8Fk
ZmgSmlGDbZZwIupA75gXYRUxk554BIb3Knfs/2YjJWlzSeAbo3W/l41o+1YV5WmV
39VcmwqHpNO5/CrFUKC4YWYgmqG40zKlvO/tdmRMLjyRC6GRKY4Hvp5cy+doZsRI
4EoxXPIyFXRTpEYrv9whVg8ich6YsFQQB3zGGHfRCQlHlhtv6HLHB27J5DtxKUkQ
ZT0FrBOCqzIaeFESHZDmgV8oNABLPUU8r/teZrYqKT8sLlBy9jj3JMYOXgPXXaMs
MM+JnMVUCc0efMol/+lum91Kh0pp4htjvP7EOBRAJ10MCOO8e2ZaxHWstFJNwtS2
KLhKGoB/vGalMS7SUZUUVGTh+PY9HMew/EFXr7ca1EaZp90i0xsa8kP9N7pVKdlo
6rXNS5mzq8PMFEpOY2nCf+++70GkPk/Yk6sR7XxTH4HhJXzoG5an4EI/D7c/LxMp
ljXSWcvJXx/P0WmToxMiXB+rxKdszsPTHWb0paqUDYzGgz+jp24YkXPIcnxUODHI
E/wTadRf81oilpvfwCWyimIgSR6CBSw/ceP3MrIdZEQmsgIKyZiWzoXOwzLnjtuR
/Hlm4/sztgAIfi3HQsUx+Ir8YHHI17EnGVeuftPrjCPFqPFH56TgPpE3aSOPgpYy
DqWNjN5mtEiwkhCLVs3XW5z42yzqkYW1og0MNyQSGCEjpO/q0pL7kayY+0h0M8yG
nk+CFY29OP6oK3nxb7XyvkQmFNeBEKr/xEAC1cpGFqOrTRzcWB0QFv7YwvipTXet
10X4y67seDjL8fm7cNAbQy9hMqDQIGKmGoEgK9rrBvY0oQKLEjYuNIu1cmLuwKK8
phVzdmVWkQqAzVGNoHDWDDU4bYbcvzYI2DMZdIzkvK+eAJ8h1Ge9BmRs2QeJsZ+s
yhdzkElPMfhpTCdbRzo1n/mUw4H6HgzV2KGtNWBeEDQe21TkwFyGGwjveOjUc6hI
FpnQ/KQewiCYKCwWC5wRH5TWQJu7zSaDKSUgHC9pFu45+OrN/9F/CTceBFe0LLld
wNhHE1eTXrkVuBdjQK7CEb4uljjC42xinzGNlSYUG0AL3ZeWNGSDWzD34djBeThT
jnJw8SPKxezISYME3qHQEHkfbL7hp0OeejHAjCubP5R0S7nGQWGlGUwhcb6KgnSb
5UZDHUk7MsaXsObC26joICD0MAnNamkwzJ3qk0ta1pbkd19gGQxExy+G00WBKaDQ
CU9N85gcDdzgH/+rcr0LLlNJ2FYeord42j2o5OANHf1GOks9aLNMCLTrE+s/yxgv
8Tb4GjsQNJCEZLbuEYDsAfBYazsxI0Egdel+GjsxNPxnHYewTPdjB3SJaxpYcbd5
rvHPL6/tFUfhwGvWFa5tY7GChp2X1xxqVrNYxykLz3WFVIJM3SAX8inj4k9CLr4r
zXjNHjvcf11GOdo60ChelU4spTdbZLJSZ9xjt+t7VYWNecw4ONsvk+Z/EAfSOhSD
1Q9qIGkRz6c8hSV/LlHhnGjiQZQA6xkONuyHzhO9TGEirkIxBCkdswoCInrNaA5U
Cix/S/ga5IY2ALiQuAcbyV0atxtGNMHLrLNWMI9h8NkEsYYMUX11WFR9gcEIYrOI
0bRWbQsYwxVID/XXzBVc40dh59cJkA9c0WuUavbOGgkaZDPvoXy+KDLG0nr4KrBw
cma33lof3m69tzVXnJ2GUZFo3T+EA75if9NpxNp/ouzCO9cHqBVOcMQPeKpwOeCx
7+35OJgh/jXSX37lJmy/qzGB0JdC5QDrKh9jNwdnKx9CuHurVKmE9lyRxEpfUiyT
5nut5kqpzqeHK+f1LM4H20Nww6j26Bk3EDPbIgavFQLqVwzT3uoEW4VFk0wS5v2/
FxzWEJNhLpukx6XPpm7Bvhgq46hRoefRgDfkUvHoseKVIBtorJkRoyS7q6H+w7bO
n6jhMOiQ1eod/3Qo4i9G9eCfkapJFWYwJKf4F3riiEb0F+Pm4y37E0ouH/Iulxyt
UpZUDUCn6Qs/JOqALYGDiBoFj9dU417jC4LLM0JID3PDXtDQK8o2kAxQs6oLT0Sb
J4Tib7QVb69dOupf6XwKpApYZdxf3sUBAJbQBEkubXzJOGNfM47Ob9DpXOCRaUva
WJBQkcocxHDgDBroYNDOFqNLvpdWqu3qTzrX0OIsauOV6YqXeGr4uC0JjJz8R4ZC
+k1BXFy9Dg0SvX5GGKM/5rxD0u8u4DZlDaYhAQzGbiS+UfxVwIWAnBrOrTUbbv+4
OJBMqy9pOUy7qeV+vzW8pDuu5DdzqNgtvXS5x55y82uekz8UTyo+EsJXIpqpQOyS
NOkncc94UDocMAcVW67sIGyUc7kttH9jQEGjgJDAWSXizSrG0fhyBFQPXowFqfiI
pBfd6hy7frxgVlfMRQF+zJvSm/oYC3VHMYk2ETi2uu/nhdcwvdV2l4ekWDf8i2AG
7sqopGhVyThKbucLWszSjUi9nTJfHaOiOZss+bH9Ga3lZb8f1G0HcOlm8uO9mYqu
RxGkKKdPNBqdgrV0KfgrHarMdG3wlsbWUH2UpymNVIH2gqVtZJ0yPC4xgNoBDoxR
5pgZojVmq2qYmFd2hCeEWhKQ2w0uV/0bdOzARKWHNMwG80JlOU1mmvsuQTXnKAQI
UZFRaBq65aKn8azEqAj1Lj1DC1BxNwCQ8tZHUTMKSdt5fUXeLaS8eXyUgFzHgT88
QnkDiWLOXA6NeZTohjOhNSEQLv3oOHEjLXd7Ls57waQOCTrCdrzS6Q/pHjo5YPrk
MW+rfKkZP0uhSjY47kIVjAUOApYX6m6ZOqejxj66J+YhkI9PtNU9rK7TV2aFNHm1
xHjUE+PN3DzSz1oBtTIjhbjfOa0hWTjCev+TBXqo0wkxOw0ECPP79lWabpWRhzsd
qzXmQZwG3OrG/4/1q5Y+ZJrpEpcRRZy4iAMNb+uja9qhzkwZ6WwOB4rtuPp8u8DM
c25YtQwZ/FJOWt8iRD1AGrM+/7uibjwtUqp8DgJit8g=
`protect END_PROTECTED
