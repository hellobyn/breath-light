`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwFuQ5IzoAZebAZ94D3H5DibW43F2IPtG6gATK7+wLxURQhoBnyNCcjyIwmwi0F2
Mcewqum++oYrrOuj2G9cuSpARpVFYmXEdKwZCynXTov6uDEap0rJ5MU1GlKCUKXl
KAHhgv0bxCoMCB2ibOtNG2Fghn4e+uKESESFhOj02x2x0DS6Pv4idM6kBDBqnGxY
QzK8EXa/9TIlZ6V+onZlijAcKncSo9MUDBp73Sd3Ml6/Akn6V7kCZ5JkYTmWhVCs
GyEhtLic9EjP500gPK3Qfw2cED0ReU2IER65Cpx21KW8TSRtBNb+gQz//Bu4vjRC
WdSEDPl+FJPqzfVFQkzP26NzMsnEk6y+wmGddugAhBhusTF04su2XH7miI0/DLWB
3jrzUw6Msrren0/mKl5L0vqvVX93uOIw9u6UK8KYmK0D9lKs8jwRhHE05bYgzmq8
IUsb3cCgro+5SPq0awse74HYlQ0L/+zRXcoLxzL5VSwJGuULcVzn52mSjOZF1ka/
UAyTnY7UZNBTB4OFl03vpwG5MVtIKk5ABedFxlHWhIaue5FTNMy71soqwsxPVRkr
IS/WBX37mmqXp7FBoIDmIq/QXAQebpDqw0G9ZWBDukdGSo0n2sQ5s2I6lcDQIp29
H9Fdu8OOisszzCZHmwNBioR6V6ATTH21+sU3LNqhsGWk7t9j9ZETh8pfY5Iw8uwu
J4gePJjNpvfe2eWqCe8Rkko2HQS+CupTnBfmymIXYVFbBcuQKnZGFsFVcmrA/Rn4
2lzM0mzCjPh77eLLblLxKQfPYHFYf48L48A/O+fqkkW9B2JGhYgMITjpiDiCBOPs
RSzjrtpFHh008cjl5OZ1tbK3J4y/KkeyjzWlBbfo4MZ/M+TaQCQIEiRgC3VFKXec
1JK2SOEh49ii3RmaLbGjhqaP/9U/KJgbXU1tQWW//QdxR3vFyRV44vnHKtlpoC0h
EXOJOb/iUvlwLJapEMZqLQl5P9p3CDoOi3acvTPq1D7Y2KyCqMyDfeKjYS+hOu5f
GPtedE6zWCfDcRgmyzQwJBOi/glB7arWj0UHnKfBoZm7dTdeewf5d8ZINzBvODAl
I2DPRnpo2wC8q2bKr/NQhRy7bKUahc7+Hkq6XwTHttmn3I6amAsN51CFr0VkEkqp
fRQ1b1rGD+nYwlMOwHizsH9VtW8UPEyaePMgZCsz2nLbZUu+MaU6Bavg2merK/jJ
WzaPShORH/ssXYD8nnC0Lg5HibL5n5VaYoe+E6wmiqLgNSYFQkbgKPFEjaEqYgi2
UYU0Kjuanu3OEW0XZoDpEzn/hOLBckYy7j9tm2L5l7UmBFrelXWSxIcl5J+xTd3J
q555A/G9KGyy9wOtU0V35htOGStMEkSeGk6WCM2CVSQK5rb73/m7ksEFrLMsleXJ
pQWo3b1Sqa5mq5NZn4++q27ycUfN5x9xo2gaW9l+3nNpKOelaS6x13jyp8ZBVYcg
yV8W7EpO/28d0w6bIwVF7MNAcg438NZuYvbMz1hWNTUnLqxEAKDKpeIe+ewyCkCb
A4s2oEriC3SXXORi7hNIl5KAfIK5xwJLY6cgRes0OsnwlkiEr95RDLg58GOb033u
dh3YUsNIvh6SAFPsNSCItYTwgjaWif7yPrhF3ClJP9BujpwpvmpDyuo/+cekbPnH
HFZnlQImCjw5/BE+eTkdxwrq/JqyRXRFLMMEtZeeOu7rT9dX9LoaJZzKRoRRCckd
ZF/l1K7lgYG7ISgeawdKGbDzo7o2cIQLgs+33wEo7+JSrFTPPCu/54+exoXcvbbM
WpTVZfJtIngaZ3LgCx5CCH8L448HhtjRK8QPB6Xh7PZEob2BQz5bum9VUtmNrYoH
7RHYfH/r8LCQzZBVxpSPWXBE9m2i2OFRi2rauZ8UA3GPXnmDiyohuYSl+tMpFdr7
xtIPgPHsdv4el3bKW4lvwXVnuR+g6B9P2Z7zz058VNNPZkA8Q7ZM6XAgFQJ7E8OB
12Js3TuDlbEj44kDzHpfRPe5aPeD8Q//qdOPZaBig4MeNqAQWrbGlnA6DC+w9e2u
p6pQgL6rwm8rYoe5yJK+Sdyc/EF+OWDi9Fxw84b4xl6qPmN0WdEvFcM/1lMe8xDj
r21vCubEPIXzFKFdp8RGm0W8B9ZPH+e5GQ2jU67bQyyV3vAxjJ/kJQh6W09Cwngb
ln4jQ3mn7PBFvzF3pqt9QC440csxiEpD1ymRopWxEuFHqlPktNqZrEvu2xbCmD6f
7yZoQ+BFwXXbHtPwlxuBEFfWd+BLi6LIV+yxDhF9VUSlmWGHi/ZAWwhIWjc+fxI6
s1a2RF66CPF3tSunuNjgwVym6iaOmgTmbcWP0s+L+RxrFbrZUYppnUNVNbRc0+2V
KKOljmEa4Yq/ImsglJKktIlzmbfRdj4USxKZ3Y7OLeWfWK4VznZY3OetjMcxkJ3i
T8U7BzCwPglb6dMCq8BLEy+X/4E71SELwQRRIqmAC1ltqe60HYbOrbDdpOde+x09
Y4dIwmCoVMpcTMSYz/rDlK5JtFi5D+RcrQ6kZbFUn/u2fhK9mZqqTy8EecD6F7DA
sSiiigVAynTID89nE4vac1s0m8XdboTs08AgeADS6yKp3cZ0msimS2AbywW6aX2C
XjgNR+XhPao0iGU7KY85JiLvimfWCM+RfHPdmhM2qDGnx1KlHAmtnP1w0aGZo5F/
mr2mO5YaQEIeGJVuTn9i57ugYAiFCTIWI894Pjeb/5Xo4Foi8/L2mTs2rZtQkehN
WQpz8qwVrglvrUKfYw68uoqo6sJDnSIzD5bTc5Rxp2RcHISXttt6DLpP9sMQBCbX
ZvYmiOJUyfTcINpUHNdHeA9xjfmgp74O0hs9HFf17SCwRgX8dOkjP0aBecTLHQsO
Y8dIXflp8PQ3PJHgbu59QpOTXuxuKjWes0tPVsQadiNeGJjNyp6SeVwnuLxR9hTF
P4c9cclagVtuf4RXJP7CW7wMxlsIlZxp9uwyeh+mWECISbBsEobLl1XF/viZq2ER
A6CVh7YNk0UYFsQfzN7bKBGGx9gsEY41nHOyy50ygAFTWL4nPv1+DoPJ9ZB1XZ5q
/3Zp2S1DypzH21eg7OTc20bzd7kMQhorwWUm1Y0gMY1RtqErNz6TBQtcRGWE4y4D
vHVVEJMERiT6NW3LO5dWDYPkC2BGgfgyxKbZq1Kel4TOT/dflPTMCzK1Ep5hnCRU
eGpGu7UAndfMT2ESVNdB2zD4sQ8aiDyKWv0ViyEH0siGH7wcGHW6BUjdFJo/07A9
rXJAVEQ1R71LFtVJDtxtqAiLAxy3jv1hoYshnuzpA5aQCbbo1/yZXkfWKiSwXJZ5
lAxmjBUEtC++TE2DPVaxee4VQi60mWywOZ4wxa96m6b8OpQit57RZ1gm/LxN/cWJ
/2KYTGtw6bSttOpylH0ycSR6aTU9w5XcmBBXOedGEi7pdYGTT0ftt3Y8Jr3ABGhQ
vPIy/es84hlMYWvr/kW/tilzbwkzaUmBQg8NZoE51NgKe5bogt+Dq8rN8nHVaIcO
PIH+9C6ZKwoBfRP1v37YtH1aw7PIiEEpci7nZ4VgQStojPsgHJa5DrnyDKjihGq7
Dg2jeCQ+nhfrBT0wwiEUYr7Xe4PAF79qRbQt2RyAyMzNHtlfJKAGyYLPYVKD87Z+
S+Fiwg0B3u6p3U5rtLLdE6+oJg2Y2ugrTuT8tEIc+kGbMvYYsJOoLiKi5t4u7zFL
+LfvtxyfDY6kVSebFWl6557UFLrVTD9sgghsTNw6oJF9cW0nGwpi4lh4mYyUsaUM
YXIm83sN3iOxMpPsJhuJWEtosiJVmXls5t0D7Z9Cl24Rb+LTQqh7d2MQfnJXl16f
85nT9zErZFJbZI/Cu/b9qxRkSC3buKn14sBjwBNwMauNuavBt0hS5SgNz73M5kDV
juWJ0Ee0gd9BaRgXvLxrpLAt/YNMB6WSrWr6ZwSyVd7bVrXefx1F9pRROdB2CG0j
nbgjI8OT3AMfSnflIMyRUab0YNmGzta0eWTKKheEQnYJn8+Qpb4dAXeLa3QQqYVp
xh6SWx+pHxvRW/skWlIb+OXIX2u+OGe/W2FmorGqkbkld3cvUZ4c+EiOSfHr4Jnu
rRaas0BDCntbJxfX0MEWRrFaM8XrZmdz526namd/EMXcXyJeTRtH+w0XUNm10lIc
/BzhCUlq+BOupzKNvRfYtMFJZDGKmAPTwl97L5YAG7E4I3j2zK/GtAv88atApNik
jStJo0jDmVb3vtFATC21hagRa6u2Zh0Ipz/ijbDdu1aZL8kxBAJMHLLnTpKTC9Vh
RwmmH1ZkFEGwAXGCSghPALj+ddYtc0XNW9pidhagqgjmqMcrOMWa3dv1KDvxu0bG
gSASvxrhmyQ1edWS6LCQDDzEQDGt7d34W0Fze8NgxbKgZdYekwUz4f76olvbdCkp
feWwjqGOAoapalDBeqqQ64XdUQcujLeaAt8wt9pIhJ7296NgxOiLBRIUZG1I3JTK
WoL/aqWypMokI3RB5N84yIb+/4GR0tXjF0tFAutgcJxqATaRvHI9KnVjtumh+Ce8
YTCFar4NLM+Vu4y86dTNdqYop90ehVBu6g26e55j+kwq0U8WpwN4QuWeVqzY++pF
sq219z8C0O0/5j9XjXXPjCPOOecGltvu7KTXVrxRYueEwnHs3hE2JxC5hznuyGxe
UWBtiXTfAbfa1sAVzwoqiyLv+SHXm8rUaydgVHHPy/aElFnfzRIbrVf+JhMZlU6V
gTBTUu8STjnOY+oLl4vWGT+Jdb2p9xLF2VVISqGclJT1dKGZttWh7lRoC9rLxKpI
ute7q93TLnYV45DGWfC5u1LmhQWrfLexlgvu6plyijhwM36Ls6gJrACsnngYYH8/
YCaalVmqAfEfshEqgT+XfQvHXYsUxaDC3P8mcZUOWp8CjviyW5Y5yKrcIHQi+55q
86ChzNaIerMcAZHyXc1nwgUSb9fhcDicNAsqoD8jObInbLym06Enw6BgkJQm9dZ1
/IAhZRUh6QcAEa5N0iozJhpM05Aj1JjiQbDplWXgVsqDJpjgEOSi3fTrr3Wed8QQ
O+jQv6nk8xTvGGdClmRDT2P8RAMSBUbgyLsgyc9CcXS7dDrUInqBFNNrD5XrVj3X
UnlF+p1se75frc/FC8JgEIf9AuW33Pe504dHDQ5ZUhxEI75KBTGJJ5+H4DDN/nPt
DfKcLnTihDEvqcTOBPjDQQDkrj0hOPi4QyumWG/5H57dUISwi+Fl3uAziOwIUtiX
AxFMCyMfi4uLuAg/iZRPSq345FJ3eyJXYPgSYj3FAox2pCStPbKmW3e8l1ZYAehU
i/pWGd9CYqlLpbzPLTuFKc5ypxp3Zz+H9rnqoIAeIH3rbkSJYVjQPAvNXfE5Ad/4
zVTL2p+f0AsjKuTRkHbrr/0j+0gISdL4gLeflZ4ZRVjB4vFUE9bEr91M6aYDvHWl
76WjewdSuKTTUy7E1+yFAY8Ya5fS0eER1ydlcyfFB/Gs3Nd6dQVCzxSqg6iGGXep
AQlB9yBdIqGCSsH1pHTgZSdortt1buu7yTWbpGduMLtibYxZtv07h7xddhqrKwX7
0pK+TOATzighwIo0D1azpWSTLjAAp8fiIr34SqxqmAX8ECfigq4CYm58zpPbNRIT
J+/Dq7UGsR1u3++oxRnkmSmnfjMWmQalusMU5XE7OJz0zhRl14Zzpz46Z8yKmi1c
BTpGQyp+64JaYDsHfqhOUvrUbJqmXpSIA6zoFkdo5K6SS9NJ+M5XvkDRGHfsYad+
sDIl0R2YE8r7UklkBPopvseH9wQynfSAVGJ+9ik0Car3bX6n56iP/A8UmKn1sHFd
73g/MxZuhnLBUeMDCSKeFxJiOil7pzkto1vdd80O6EMnnabTWo6vuXwD4X/AXqyw
te5wqPw0XRCO8GjDopC4drlXSF1TXcS3JPJ8KdyzIE5YEDqMnzPFk0w6WnIm52Jl
n7alXpXR/l7dH1nJqRf4JlZ2UCkWaPj9JOmvFeyxVAFb3RotS/1tQIeWiKmGwuJM
Eayc8ljk9lvBE2waWLJqjMwdBvli301+2z4RJpnbJw27LKo628C51Q8RUevE/4pf
eizTGNLSUxJ4WRTznc2PFtKJWSbSG7LUk6JmtgenEPMamnOJ3Q6+mdsIrHJltFDK
ViF6BvSUHqYmCIi78VgR++BfEI6J2oEFlsPycYGhcvk/00FFjt+4wBnbvaKz2osu
pwYJ/etFeF86wYo1CJ8i0pl5CVFEANTRdK0Ur3N8RzLgtY24fJSg4FOCMxUJf8pa
/Yc2rHLIQwCG9tAG1L8we4TK6ZYRWD6rYyyvHiLgSbTvFO32AKIdRN3RCS/j+6D7
KnULp7knZ8bxmCZRsW4F7Af5D9S6OwjWcSpYUNqnDxHlD2QUYjN8hH6Ed4iIBHqb
3X5QyTj/bRSyFXg9dn+5L5qsdWxJ+9Zys+BaI7OFn4Q4uhZO5Z7KOxxBbLdYMsgb
HZBMA7I0BbibcB29cJXU7CVo9VOn73Dxp9iwBxWQX9pnip8Vo2kd13YdKWlG7HR3
0M444OllhjwJKHBiB5wSolGSN2RK6mjufHrVIYgrFUSbEOQJnLP4vOFpddpBFGqN
K0aaoYcZY1iK6QMo5hZ9tM2T/YKvr4Il7zu3lhtulmeW7p2gXnfwQN6ufz9v+5V3
R3N02yOOM6IdaJqY4dWt9pZufrYxRIt2uQyMH+2DddQ5mtj8Myy5MkrQ6Bfb+G+V
FYeMwA5/x0RvA0Sj7u8qFLR3v7utsw9wI8+olbYR1J94IRVbWPzU5XDCWxRf0JLb
9ut5agKEHMmj+w19M2EXcPFnqJqZM8rnyDNv7MZCGx0gB+7wjr2W4hlF8p6qNkKU
yfuNb6DC7euYUFj8696pY7xcS4pFC9mOf13TWa04krVIehPWxF++e6cGtR2Rg17F
lRgVqddNutX0WngwhD+MlW0ORU4HiZ9F4/4X952ztByDESPlGxY0CUC+TiCyHjWf
GU127s8HtSA3ExwPjPKrT3AF7Ms9mKnyzns8uRFAryIDh6GQKf6hIyY6MZ1AEWCe
ESc758uIAGrA1L/AAlGh/ryUuUN3csnu2+vUxaSoooVR/fSrQNZqF0yDQodTwzrk
PKpkcE/KBmaUQANztI2h11GrAYI9hetKc/wVh9jgewn97Pef9F4pMw6M84mXxjjk
ZIDJAzRgV0HSNpbNzkOjlYg7L9EI5XuoE5mOgmgajCvyu3rDaf0x9l/J8mspLwm0
nFw+l1CwnPh+gN1zfc7PPSxAIR88/Pi6tGyLBnzYGCIgO1wQHkjbOv7vL091YZY9
sJA5dRK+a2kHzvC4uS/RGfeC50flXrBVrA1e1gKVGu3BKqKcd+pYLXJ0/r+aBZ5D
DJgDFJ9KIuXecXYlgK3TwmZ4rnc9OyDUEcIrL/LE3MRvI6rIvPyXWmzOri5aHMdv
zvUgM0Y71aEfik9ACD4Ww3+US6wL9iG0wZs1shoMgWDR1gK0EbK/RsE9nENj+20w
lUJy7x/tt/+Vo9PdbPk2r7ICVnx0YM+96imWwXCN8ttGpL9zKgdJ6zKbTjG9Gaa6
shyXWNYmNCaaENwnzTNLoA==
`protect END_PROTECTED
