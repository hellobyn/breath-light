`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiU4buhXB/FzCRcbiYgiWRjXcYii1CqydBgLBlLE3fLs5PICktkimtIBJnbVyRRg
HFp4Jr0gunwDUBUGNSjWmoEv6965n2kX5qyUc3rvZ5JL4Ygm0gjEFPKm3KvTTl47
kc0VdNkXjB4DrpvGMnAujEwPuJS8osLZsiCHN/X2rYVzyqd6xjPYwBp0E/p/5Jsn
mwirRmy6Chuy9940tRshnHQV13YYNKrfCOuw6Fn3BTPAMAiQfeQjM/OGjAjziyc1
wHf7g2rdNbPbKH1/2BXK4mI3xvLIkJXFF95xcrJQLSqfgMWIuY4LpH293drCr5qY
OGOi1DVIFOmUpU+iXiYJu2w58kIW9tOBL57rUxDzXzi15BSRc9irRNTSp6g0z5u0
IQJ99WWs1H2X0hojrLFTTUIPZ5E/8n/NVddumx3LN6C7FlQ4133N/DazwFZLBnQV
vaIyp77k+wcxwXSe/5bs9JqwQnSbaJWZClImEH19lwu6eLWjRIYoOieBaRgxKt4l
lGfiaBqRccT+BjbuyipGYFMLmuTLNoPiBSXm4ym3y+Z5iZ9RxWMEDGu+BoQtNu8K
TxaU0cBZLRYCR664WhIFRUeWpgnqlzeFW5lmowSDTKEHGJJZFo3wHDBwclOVTh/O
BzMXbMC/y19PN2/UfsIcJtvYnUgt+QAbj6zC04+5KMeys9K0d9An4g1oPi6D2CyX
`protect END_PROTECTED
