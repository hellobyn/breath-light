`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VP74219SgmR4oR5HY2Y262pusZNgNdFAWHXuFf62DHbjEiz6o2Ni6aIAvSVTVeX8
HLzZO2JPBT7Drnh8KyHueaxcEyneTQ1ohm4beMhrN12lLk7qqDxiebNKmOh4S/NZ
Br/eNRiBuAk2wzV4DzXAKQSS6weRRmdnclogEuk7GMwq67ZDYoxG58QLT6pYhdKn
CpaclmZww7+A7NWIsf2AOmzjoDQOtv6T5wXnJIQLH5+KorJCCIdJ6AuD0crKIou9
7rahs6k9GQSQv/AZwzW1GcocH3KwrwWY+jSkWP8834mDLxPu1MqXPtlpf25nDv6g
wYnZaZJetstMKXkkC+OhQWPlYMEgM/N1QxaaVxg8yQEm55Y+SR+e0niVr0bwTgLm
6YdSt/tBmykYTpEsOyHdD2dNXq2iRWeQPH/B95PQiZ0SiNuh0c11019M/c0kRLkz
Q6utWa09bDMeDLcRi1tvBU/trHYTn3YkiWoKOgaGKE3BIAH6JzQL5CGH228L4d1R
YZG/RofXdgZI3jt6TaGqZFDmaK1zeWMVtZ8E0jkA1CAlCs8nDwgTRrSG8BgJxLvz
JlKCliOs31wqxg1/XDBlnb+wp2DKvLoXDIpcfNpAbEO3y6bK61L3ZHWEX2GhJnL+
hzpiQ+8g5oSR1VOB/cOISb8GWwCUah81J66S1mfVvZNZgso5PfLSlkf3yNMmrdkt
nTrId4UxEDK2u1361cd1bH9reFHeEgmcnPwURHThobWhehxjS7WoJj9SxMPkMRwB
GWTaCCUC2AQyCSDRy5pO32aOID5gxToVrlfpJVK8UQYVtYSkGd8bNkiBBg7jgqGw
EaauLB1fM2Wh8ZReefcQqjT8BKmxSYMpmJbazr1F1rvXJk3i1ptLeHrZzBvG29a1
7WjsLWbJHU3WkGaNB9DBk1kc19paQCi5P/DjozPfe5VIVChiuTKm1cGCgew9uAuo
qIfyIkPbTMcCPsxeYIjpMP6l3Ju42mcLn22RmkoeGKtl34sKtCLQRPtUExOQmE7U
tLP4ois9kyw0tPLUtMcM1LF8XLQSjeMB+SbQzy2hL9Ui+icJxO1vEbnwybck3k9u
d897qB4BdYmDlRc2NlZyUw889ckDuMOctT+uiSl6b9el5MGKJ6ha+nAhVI4nfK5b
hZqjS9CE5841vZM/GVuKB5zeS6X0PWNHuiga8DiGUEvxGPqaGcBXgEfRODY2yw7/
piIN7EKl2pnir47HsRXLBqqESHNZto4cRoHjSGTVHeg=
`protect END_PROTECTED
