`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHDHrocXDZ0DgXcOy3gK0dhEw7raLNyv/ZJmZ8I4tzK5nQ9RJdWqpzsGrQzMxSaJ
QNHZNs49S2szzIIzfPLaSVvPQhRVXRbrflNTDg2PCIDYNw+Ri93OrzUCwCyBkP90
TPquBx0v6Ngrn03ecaeNbliTOiZ6rtZZbAXKIqmqXYaTqg5IvRVACr+dbReT8D0C
v7VrUdRIy1+BISpfQ+duYBrIV35xKHgyO0ueywaBOG2cXMojnayoQxASAx7v+6Zu
SEvXikKCNGi6jTcE2iAj0PyjPhfWUdbdi7ggx3Xg/cV6ybEPtxYK9OCTnFcT0+0s
u6rJ/6OGBnqPwCHmZxtYmk3UJG1KVJkbLWk0E5JDy5XKp1O6k+0MudQfhCyk24KJ
H1+vOK8PljcdUFdQvi+Y1Vz8XgK+LSzaD3TsmMrxt0g3olTH/dvSj6vWYeYmXDy7
+8ecxBIfKtXObdYNjwuk84F3dcqDgqr5lUNfkf2lu7hEdB6xS3o+MMuAXkj5Iz+h
TyoyD4Kr/tPz1wM0IHzHz+gu2FlzrsHsgKZWsgauluKzOJBgzkdFHJv7h5uykOlV
o7qos0hJs/syGdw3HdAAkFsGsCgGeOldWbL3KJtEZn0YjfgEHnjq1HpN4zmdm5uF
JboJUJqsgO3xUaybrz+6uemzQkWXm7ZcIqAQbHjge+k49OxXsXUD8a8vf11RbkZZ
MGSRkLcQFsiDp9rF+PQhL18ihJVipA+kSquBEuelOL1hSNEVe4m3xcHBqKlDS1e2
4Gdng2RHJrrs1NLFpr5CkjSD46kfCPG004kBnt0VNd39L/Qn1oqwkB6asqcZyjRl
Skv5dC1QtkbwBSpQvP1O6QBhvcAXfZz1fJ8TLepdcV4/4SC+8P8XU5VXHrX41klk
pRAlWGrDmj9EFueMZ6yVtw==
`protect END_PROTECTED
