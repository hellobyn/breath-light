`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYqRGMMKUMeQoaNrl6+jAw5865a+pz+08xpu25NxMqt9lHdfKEu8OQakW7ocEOjS
9RIDxppWH5oZpm8gq0noOY9wS3eTP4pj+BiPX8pI/LHQQ3vBPK0mFleWaP9+4ixP
PMdamQnD2zRSHmbcjTvNbH+ULCNmGNzWOF/mzCqUKDLgSE9QVr3vltmH6in05UjD
gTr02uAc64/xcyEvsPH/kmo2ZzH56nFUD2MQxNPihu3f8v2upco1hgPze6EKgU7r
M1d6nZlzcbDfAQ4lwmBhqxmGTOfVbN3rofjDwXY3Xy0rzr99PVraKofjcqaAADTZ
MZNlpBCgIXFFuryQrrsNhw4Kh++o4d2Pk+jbzVrvhagPBkGWSpU+O/AxsPiDkx8N
21Qb6lCNVbtZjhoIUhTG/ymcPf8seoMfcEr+NEo9Xnlgfi7akbeza1gATnGjU5A/
yTwzJP1jgCjW0917qkRhHfHP27lhd4/NBO3o32vCLcaXJi0Sj1PRWmtzTly5mW5V
vNkORguxeQiAH/MqqhsN5IcCdQUKzNIw6PEQLuTxXn9SEwSRP3q3lTowfJIBKuMZ
z1OpaD/g9qcwWvDLbBrA1d3gyM3NcMf74K3P87Y/QI8K6D9iZaYvbpADH+VoZRoT
2dsHPP8J/inEbFK4jQQ+jtCwo+fHUj4dVJeSavoUfHqRpJeYiNE0exjocUgnCaBS
rQlpXRtF8xmJbe/aHrpg24BIB6ofSzkGmI8CZp5/Hx3cjSb6EneCQ7g/NS9xQmkF
J2ywiBFH9NLR0QArUkVYQb49uOU5Ab++ONF7yUZrzr2XskzIgj0ZnHkjjfQgRzSK
LVrbVxqbFV/jeQcSCfG9IVQ5l+P9+uuMQ8979RV0boBeZgSsqddnaBgwnjpxHrq8
WrN5naD/tucmWS46WQHaEw6wjHYHjCNziRXjvqKKuCR1vDci3S7zZc0O1BgNp9Pc
X+6aP58qLbn/zWcpJ1chWh+MjHasfbdVQ39/DCUjrwed9y5yg+DEEubDzbTBm+n7
X8uovtqHRC4GOotWhWFUqxnKJ8+Hz1BtyUEenvlswEmfw1dD7aZWwxAb6NE31O9S
nnKUgKFmGrqDAngQkIFH5nVKyhAHl0ct+8bYrAsodRt3ek1+1BVbk0+55RuP7KLf
/HgUrXy4cw3EH+Fa86bKs3t8G5mS0ZI/oSv7VErsGpx9F2B61Cb2m/E4P9RU/Vpa
tUXonCrfmYvWKOMM+TRH/uTqvTJneSxwnG3G2FrO/Wg7zliM58JbDRCvlpfivwE1
LqYTd4T1b1jz0/qXj3bJqUlF4KpwK2ikKBRIh4mCa8Wbnkww2zgSlTaubM2wsUXb
rIkqh2gVml8kFLT4D3yGlw7twtyjN2aY9ELvYW26AwRNiJdbxGtZIgVwB2tmUpL5
px07bUL1oXRJPippczvx6Dn10XEMxeG5zvahCwnzGGTDtKDvx+XgjYntWVPTBLkA
Pf4EvY4yv6iakbiMmuJdKaOdMtpOLDKUkh5mzNG5QJRuz2sgY/nehfI+yLu4g4XO
xYffHTNNw+Hyyr9ORZoIxrmlTmY0miaQF6pKAgctOdZsGLGtYvmEYuPzPnJr7c4n
xDhtssxO6UHW22p/XrFqLFXi2UhMx73cA9KVGEUczXmZDq1Vd5+/GfPpDrWvGa62
uMp8PEe6LlihaDXBJPZS/azzM8sLkNN3a/W9sf3THSMlznlkZcs0/ruwMvV2c8JI
lYl8/3holsdNHN2dLeVZjJywYg1Y0f1CE/HIj0pnKNhjc5KOxPHLgsAdOdG3o7or
VIHnn39AnaJ2bjgo04qHfU1AlmmsRg1GqI11WIldvw/dadtcueSOcEVHolLtUpoA
ikxZENkAOgctEoHwRNXQ7yFD+ZiKIPqWBm8bwoyQ/S2fHSE7EqUEwnWja6f/88qi
hCM4b4q4godxkPLUGPdrWQs+UdFGxxYKjK1f69YX7Km5HIwswv7j3Y4DvyPcpb0l
8KO5vBti08w1w1fyWKMZL73MuPMsA78Mc2jEdhpyNcdjR5/ZXjyGs72p127/YLI+
/1/QX8jap8bmyi7CaUTPbbEa10gCPH4xoJEPqV62gX9gfLHhPW6vhoS6kkuiFNdN
2wp4P4zHx9Yer33OkzG+AU+aTUzkHM/GO3FkhDkQS2cweR6sYN8dS4aY9rMgNPn3
e0ztwmyULlu4vrkuB/DA1IdqkYQ2RUNli7QXYxTlWph5R0L3zepUQnxvuUyN5s8L
rwL5QE5UKUP5ghE4Pt+I50r5RcaTPyWtZVPhcPGIXeA4OXizkTWgyONaWxXgUXPX
DoEhckY4/h+zy7SMENRAOrpSlCKiLtpULX/JRaDVK0F0TaOir0K5gt8lAtsRhM6M
Wyb5oeCFRFUn0ARrlu/O+5KJ3FqVlqnYffxJuUdUZ9RULoi1a6yngKvDGvNdghJl
i/BkTjoUaQZlowVX5OTI4JkMOtN4wfXAxLLVhrNgkQChbmtZoqiyMnjH16l+a3/D
98RZKeRR3wGTPykcm9Ht472oqZZEA/33MQ98Kj5Vnk623KQvJZ6mFQcbGHuz8V27
fo8o7BChoyv4aIxeBEOjX4VP0fMvHW0KSkcz+4nGfUhZs08gj+OmjKVxFYLaKDNf
aOe1Lh8M5B9uICC2Q1RAzWiQasdlo6lXFGWKIAtq7QbboZDuhFm9QDosTVvRd5fG
KFsEx58fmu7ivo/jJgh8Rd6f3yYaQHZ1djSSi3407aBWACYKj5GfKpV3WwHuRZGv
tyQFCJJE/Bt0iLQlMXMtjA7ayGX34C7qI+igYEQESqlNkrsCY4+Eq2xY1zZzNeWr
YvQhoV/XKC3WhkqA4BZtGvoNoykfMH2sGoQHDeIBkBlFy4M7SVote0VOQguEkF4S
nC66fMeQ7+SWZjsOtHJ/jBKw3zp+n9uXMKCAQ43gwuqm9IXEdtfWc0q9t0H2BINj
2kcm3kF1HauIB0qkFpoA0OI1zBXYQ55uM6sowuQ+hhSKdO8yrYQ9DMNU8DlAlAiF
33xjO+3e7RqdLBfZ65fvdRFrTLqjwp9bjHk85k/D3LaB9eg2p6XkFGVNZe4LiyGC
VUx054s6d3ODIjgYW4mj4ukZ4vvobE0HY3bmH7BQWr1Gt2YR32UOHhn6CNZL2Xt6
J/4EzEmozU/JNvOQxoWoBBAwcr2o+gYiRUat3PuJ8/J4LtkHwk/V4OKR+Mpg204N
7ic9GDXsNaw5LGNhIckZ2bqRkg+Z9HONhjvEI1D5V9DdI3eA30dk7nk70jZUjlGR
ieohtqYKd+R0MKcmT8wqol8qShahth1tENfmKB1a1QvZJVw2dwdOIBfvBRWOBZd0
y9bkGK+f5eT7u6NLgPtYcUMZZ7t6U0R2M84kzElQL3pCmF98kxbOaSz73pxTcGhb
o75wi2uy7yh/SXYfx+zn+MiOESB/EcSSWUw+7lLHKf2NQXuanwjaSJduwc/t6Uyy
La+Tewh9ttWQJV/th1roIwI4fAsuBi5dnbJFZ5udAIb8FEmZ+SczR6Bs2xYgcUp6
KLzFXGInlw2ByhuNDivGP9La/KynrRJzXP7OqjYFm8gTGkhdyMLdS95bbhM7dTNX
PYFDQDjn9In+xVFcVKe2M/oFKljCjAtsNS3CdV7nJZjwfIoYb3kv4GpCioyZyc5c
dHg9PGJveBXryyE2lVrubpGggQjX9KwRyS3wFXpC0SfBCikdje523wPoLfe+nGpQ
UXBmZYWnxcUCDUwGOQmasJXyryCjsqdTFallu+AXybMSFWVnFcseMrT+YnKDEC7b
VzJivKM6IRiJuZ3bZUNILKfbCoFkrkdMqKFietQDNCMNf0AnPzVui/XoUsVZp2+u
Eej0Tk+XZIybrzpWAm53haqqpQHcL4tLtrDTsAgoBCzPgIk1jjvT79/qs5YZaOg9
9cDm/ltrl2qr33IqLC/yd1OKPz4ouLFmiCdP6NRM59O4LJ8+TYxSxxa1n+5TGdH3
6nIIdC/PyzRnf4knJIWaBK1OuafCMSlvWa2C7gM/e2IMeJTPsqIbkVgIneEFvByn
4JlrivcUFKMrQRklPYGjPEnqW5bdAvYQto5Unnm5+NHjqcmpATltadxnGUBNWZz6
VvOGTUTQ3rh7o1s30zNnB/Bh/3ofaP1Bq2cl+1h9qO5S9OAVIYrljD4h+SV3FoyQ
/4xqKnthfsfSWZIlbycx0A2uPBilP9qxLDWgWA9VSwUrYJwGPAwyteynaTn6zcDc
tHhqzsuaXRjXi5V6fRKGSCZ2eI/s1nDnp3naXeFCZ94lrKXHfAQhch0HnIy+RB+C
XHPtCkiJgW40UeQgShDBviKxxeLfB5Li9LgFFyccSA47/tvC7/ZYxaX/2yNs98HP
7HZYISy61vRgR78Q7wa6nxk/5Zd9W8Gw6dFqfdv4b5WztW/ZEOLQuJA6GWa3YwWY
y5yd39GbUN3SCGgAKdlaxrxE4BWnh9/7Vm3R3+zfJu/O4MEaSqReYv8zpLk3NMGe
6qhbD81UdwM34fnuof8xHOJxf+D16kkyeVrSRrUt2GnlVAaUFy7oAH1v2kRBi6Hd
y4AUKkGyKwwBngtpy1jrgmzSHKPVLDcE2eyCA1Agbb0NmJO/l4xUl2prymhJUh2D
HD7aLGekddyBdW6OY02vQ1TOpVj5TkLiHMSpqhUR3Oly/I6AthOaDfDurDFjHiY/
53+FzOziTct7Xs/RiTLAquy/parE2drQoFBgzLJbb7XZDHfbp2AZjYIwNv4N7QZn
kCUO5LtL60vmtCx/Sc9AXJFKY51rliooJ3Qfhanj5lL4piWJUJ/k1AHQTh0Ed/q5
`protect END_PROTECTED
