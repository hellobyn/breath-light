`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUNRAy3kIcMf3cxWzRxt0iUHS/Y0ces5la2tdKPTYwVbVL9BtrA6Awg9Vc+Dqg+r
dLtxcbPeZRJz6J8G6Lm8Mse2mwUMPi948Z2oBLSXzdmh8g296qCGn6CxCBs/QD+n
AUgjY5ZxZsNwvuhjOSZsi+cnH1LCH/3oWwXztbpayZZ+JKbEXtaHmkQ/SHewUSQX
7bfpY+Y09dhm+2j2fp8AuITDgxLHiUsCLpTc72PjPfSll6HIr/A0G72EMGlajoQP
psXxUoIPXOYcAcbvODVmu7H1ALf5CWdJ3eXYzHa8892Rb/pBxkPMcQTNZbw9b5lx
aJgbeLj8t3HUSeTtoKfM+g2F9e1Ywj4IzsgR1UkegYkJJm9O05A93qhjt4CKa7RY
x952Cq2Sw28SRQHx28/NSvCx5X/Z25936SzsfGl6me9gJSaxEcjoVGnYAhvpwyG0
cXfZg6bLX2oCG98IZ5JmV39BHnrTurS3J/T5+VDC2ZOU1VMql6MVTYZyr+xnSUO1
ASk1NBnjv/rCxAfU2SbPMw==
`protect END_PROTECTED
