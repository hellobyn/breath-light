`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jufyS3BTqJocCqKFx/esFTuoEUAYcVk5xQl5DYBeCg1yMJDG5/MoxsaK63YFJZ4P
XBxQPoGqS0goF6YeCuJhiwVo+Nxw35qDlZKJjfjSQAwHUdjTVN4lVznR1hFmWmCk
jMbIjbyKzvjiqH1N4BGDi26eQTCd+kVPGcmFBeFbXBxOxa4YmFka+qbFXd8o8+Ap
n4A4I+Qi9GtBkRuSicvG8U53sXGRHXmqAt3BuQVZjo532zH0mrrwdZ93jZi+Ri6e
A6wXWqihSb5VckIHQTNJcFV6BvV1vE5LpMPBhdME5uDn9KPga43jGQCx3zyyr7jd
7/RgODCXqP9t0DZciTSVFzLCISN8ShAGN6IEsEpeI4E1SwHQLBeLorjA9sUyU0s4
WmQztsyIwLd6GL8oA4wfEgjNJwjtpcyskVZUiPFPGICW7TSP15PAApJDAqRTA04J
rXZP8Hw1niOUG9UgicCCNr/enK3d/GmJISvHqzjUEMe62ddKT0IRJ2DZFJdzQiyc
EXHbjDpa83gBBLdxskg/P2F1HlmsgozLyBowFgoTPnywfEmNBtivVq3c0igFCyYb
h+CVnWl5d4dX0XPbkywBfUEE1kJdGP03gTolzU4fDdeKjbJPDCZyQAjiyYL42dRD
dSTBbrRrRTLa8VTJomBg80ToY3FWtIdQUvkt7NqlUaHG22uDxae+d/oun+rA+JL6
0q1X4fAilvL2TtfFhjMSAAvGFbHuyn6LyMQ/JAK1Am013/vhTmIizVpD2TefhQvn
+7zWcxZsr1XDy9x/vNtjhQgHXlHa0cDQ5T3aoufHuA5Ie1m0gS1QS4T9QNfxq4Fq
S9k5UlKRmYJDqRWg3WxbVT1RVl8ohl+jEEpuagnJ03+lRYaACYxDbNOIW6KfGsTo
mx1HADTzTCO0l4fnR8LOvPPlCaZBp7kaGF4yWmb1x8ojNAgICAdvKpl4sVrcHN3B
soeyqtj/BhWF14KRS2wRycONv6cdgrEygWaR/a63/BI+1ZpCRldhrJ/4EcVJZFuR
x7EaLfQAP41vRFCr1JML5NMWmKIJspHVoFZnM5M1Eiweh6ARsnxaxIbWVqVQGToy
oGYpc5xX07I3Jxr2mAzX7Z24DzPtHHwb3Jr9VGbEjWkIwQNhOnb7l0omAx6J/r3c
QALDfrhUv8IOqvww4Vs/0HOR55s7B1xm3+44xsDt1gfyiwrn8lPXkwd2QPrRzw8U
UpTIdhratrU/0XoDnfITnhewcJ4Vaf9/s+tZWZTttebpOpXQhv4g/JWrc3GEemXM
xfTmwyLHjwWg1hrL641tVTq+8cMUUqZiHo8VzG6a7oEbOsDuwYLcDZWc3NAftKSl
keuC7JgaX6itJC1yinqAeAvF2aVrpFsW3AWN6juO03KDYxBLcq3A54cdxuSfHQwO
h3qTFh6fCoe2FY1kWNd+vT55v2JPV4uWa4HQbj4CQTKhcbPyojdzh6ZOxLDrM9jG
Zwq8e3vy0ga9NWvBAorOVUPKGOxDY2d7rvpOsnf55twyvIKObSkv1ig//iXy92f5
gIKttitba2TGUPHvxOVgKtD8v+8vUDOHnHbo92CpIs5PIoNiQeoJaDEeUGL4yL+7
FKoZ6SSR613bwp9lbk0e29c/+J4VWdWa5949+tALz1VdJkB/W1XqWM7yUe6yWrOL
94f/X0rX+QfRPVVcf6yD3QdQLRgWrNA6W8tiURVs50lx08W+ivqyOlamhWSeXF9p
xDdjVd7xi+B+6dA3gJSHYnihuY7emlj3B3qMtDtfJYIkFPlRvn4PGES6qit+WouF
0PZj7I8VHhn3yg7DukiaVrSvhj/rQf7uSYFGn5qF8ODCsdaPBdNrN/Co2htbcAf3
UduF/QF8ov5msLLST0aI6SK2nbN2pFDl5LRR6QgkAbV0d+2LbwmiUl0OPCfv/O5H
k3aFWfgim5JCY3w+W4PRP/ULfnJLKl0+Ox4l/bUUeWx1chePGo9DptmdUwj5H7YS
7IVUKGmdcjn3jPoZ2Dr9YhxtjimPGXJ67N4t/9aL151pW8Dlmas/B2s29RUZfHp3
P9rijs9e4gNCT+Ir5kE59WaEChjJUv5I3lVLO6c0hsLKKgfBIxtCs8HdaIQfAx+7
XQp4udvSpLtJHS8Ui0wiB5r1MFA0KfnMny26lTn3dDr9HzhUN0ZkS9WbNehOET14
3jGy6qHpZXqHS+I5hlohW/ayO/6JGrnmWkdC7WJGTbxats5EZ5fvkhenpXnUwNUg
XHivJlDvX1Emo54ywvhC8Prwfq6KJQ6Dv2nnJn5F9LOataP3q4XcgFlWtKnzihWx
6bJhgCRED4xf4t0wcrBax5wdzBgyZQGXcjeeh1bDg1evmzZy6Bx5jUd9+9L1bP8y
/LxlQD+Kjxm4+6Jjz/A4unn/HoIpI201l0tNLv1F/Lii7BOXFjN2wFcKkkdn8h4Y
VvE79uU+p0eiJCUDAnEDfIz5T6PxmXhOYzHRnrFayV8rXe8mrORf+Kr1dzST/6Z5
cwE1Cby7pLHokdbj8nJV7xRqmNhefMsHT1+12Jj0Q3tzzlYSleE/OydWs/WxABKU
OIoKgdbcgTyqSeLi5pitPkv2tYYD+UO5RzRs8H7UNyancHkplBT70bgijZTXoCdg
DCV8DzFqHwkEGWk83vFLgTkclHMfdHd/4KZGn19Rg68wnhhvreh4WtKljFPqltuR
APuzJ34YB9dq3GXDunk8Ex0HTcuftnS4sGprr7zpd6nqCzdbRCsZrBYV21AHsKrh
2jFGKWdUR1hEMmMsGVvG3JC2ckA4V1rwtBDeBc3yi9ZaqpJpDjTvdDIeWkfJHuiu
JNp1QFSoXorImR4bmxdtvAgAXPkU0MROHNqt1/UIukARZW8pb4A02lYtDF2HZlMz
BHtKyOBHNxWnzVJ5uBXSf3RKSMKWpQn1RwAaUChh7hs9GxDCGmkub/TChtmBvtm4
8ms3Hwgp7RBKAbv35v4rIWDNMQkW2JlPvNulLwEnsufbIPm/XuhCjXVV/+uenFVf
i9ao3fNcSc2qAL4xskk1pLVxMt5CtbsurvuKHLT1EPkJKq2W3qGV+aumjplvLwxA
N3ovyRYKJ6/jbVYj3/NoX96VRKWVBwHp/27sggiQjVWbkfTb3NHB0l6WX1bVfO8U
Q1xmXW7Km20WI90q21TqvQE0eKCUCHBqINoNsLikaXzp4JxCvuEIK1RZnbcIv6rH
U5eqdjxJg11Ryt6Bb+mMRKBnqE2J2m0uP3boO+PHoSHf1+1WqDjXN0E6OrJj7P7l
ZyNln+ezBpzJIxAUMnlH2zTRmnZnoC69cDAiWxGrYdIsmGawa9VDRs++zKqGyxq2
kNXs99RDJWAV/GoX4OOjAhnRgvN4CjN2k7QEXo9kcOJP82kjGIJsa6yJhPro5rEU
z2Rmik80QLpzQAiHJcoSKUOEED14riVi5yZ+DABBt+0pDgXn5G6RTFF/EL4qPjEZ
eqgFU5dSzxfoPduDmMqxMZoAQp8XNCJlRtwyWKhA9PELf+9fmH7Q/3b28n3Q4WIZ
YGMf1e6OruBhI8UK0vhS4WXPVIFcoisZ1maUf0q/rU8NkkKeNrzUawExL1YEePdg
MdRR6vsK2l+vMuzRf15alQHOVb/fgWoEDHrnyq1zOMAIYEt+X9UKBwwQKoJUdspv
ssTSNvYcjGh6kfVGxz7AJ7zgBb1UQ7MmCl7Ab917TTCkA5Ve2OMdfmjdkgMCzWhu
dbaIeWY72ZU3+3MlIogKBPYgIHP0hazv1C1qr9vgShij6syvOzbmRaWWw2hPWr7X
ywe/vQp6H1i5O/x+H2JW6EDToAIEx/knAIuO2pJHvVABUq+vQKtCFyh9mtNbs2lJ
3bVfWuCH2vpo+TwIHv7jyLSMn8pqVgOwZlrQSm9pOSkMiVOzM0ovGd5RqB0R8A0g
5+nLsRSDOmEx7iFhhewIrvoflEUZglFaxFNBlcipfjJQnEo1Ww5TMX7xPjgC+15m
R8gcO7NlAQJ0zzAnoZVrwj0v9afil9LonI2AK8/9vIAhmOYK9QQx9xDyodfryPTM
96Znwo2e8h7PXAjUNRweqjXomy2J4soukMitwnW5ZcTY/NAfEcDXaqMvzcqrMKl+
tdnGAywwYZrE88rw57HT6iHvn7LFm5fVFK28L2mcUTMA6emjQlTBUQHGaH6geVcG
fW/4TEaQCwxsEi5R3XbGwEXwyvfsII/5ydFcPYJ6egNvEkiuCAgteGG1zbhgEwmt
jnVXeYjrPBi7R4NNFx/5VutrhBptFNq8c32GF1tM/HWvmTdS3mGRvWbTwRYz2jpy
fxocWfte0ZUyw5AR5tDNqc9fvNU2A0AhTSpahhz5rB9S0BYSswnalgBGvmWBX1Dd
Yj4aRw4256CcvPflXBCGLRp1LNzqXnbjl8n/PLxVBKIclrWht/kAIc0ZHHHfAESJ
O5ymCOyswG7xZ05PQGQ/jf0MG42fpOcru7g82kOUEmXSLpPSbJjeVseGo2o+HxCm
QMnuAwZ88EB7rSVMZOZfDBTnHZDNilsMB0Zq4M1bu3M2h/+Q+opXBcz4tVs2AA6h
lQjZ+ntVHWZMw+mS1tDBnQ==
`protect END_PROTECTED
