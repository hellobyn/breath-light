`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dXzGj8lAVUW+m6D8y/XWQfplyVj1eon16x/pEq3EeeqLPGXskrzXc7AlSMDi3CN
9KJOBwMhI4oNikwAGVxlLPF2+G2flw33Zun5VDIt/4EPzJ94YZS24f8+ABVN4r4U
qMjVfuw2robjoYm66nPydmhCl8r0R3c7duV4GvfbfyukpT3WvnxGuAY0nUHMZtxJ
4Ew+u58b5mpcQcPGewKIDjWjcSShnsQZ2ezbf97dG9jE9ehNCPoYsUQxnNAwg+a+
RW3Kw0tt4XzncImOMsEKZepUrteVCXF7HLT6Hcga7cHnFyiwQU/zffOBJ9BMJXmY
7Bg0LjqE5Vuha98qSa7tAhqHbCZsm+SKzUpDtZfyTqRckbP+rj7WEEzkXKUISymG
+WNbJzmdcGEje5lc2aokCkd1MIXn7xYFKWATObSOwqknrWeAIvZ8rbLlp8fTOr1U
218ZlDHTJNnLeWTtCkRBY13kiME2hOC++k6IVHc3ChGLT6Nmua27dMKRKFkHWt1S
/RVJgcHFdrCb94rZPlho2vWW1n1PHR4GPZxGs62BBN6PmZTP7kb9/imMqIZxfyun
yPCPnW+NhOdw3f6DcY6svUVnruhbEk4MdUdbch4+CmgNJiC86/CR1/3Nk3P4Q+22
08F1WQSThkoQ5Wx3dcfvFwL60I3WQDK5dxdJcpburKesgfWMekXqC5i1VZuc5R4D
ibFNIpK3HWOJVp02E1STr/pk4B/UBabebxTUPX9cOUDz/6DqzlNZOIu7aqYzGc+v
SnekFAXlJLbIpzh9nlon3KHyj2oVfpGVgfit7JzFo3jJJr5+MGuU5ahFuKLxwNNO
1j6QriBM8q9WYSUGmdxVcnUAp6gpg7M8tOBDZtluOSvkc9qk6kX/yu8osoXi8PaK
IfKQfajCyJswQxIujvdXaRlpDKcVAxc35SbJy0VU5FV1vZ9g0EaLzID5B14ePTcH
QE5kMRqgTDRNundiCG32TpiNp0h9QD11kbUex9ta0dL28WoDsiPVXOOqQvOMpSxh
jpN4hzELItOcNM9pD+gE9g==
`protect END_PROTECTED
