`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHlUH3PfksaxvqXuAhGk5b4QIuONkMqd5jxNObaOwyT9IaKZEMoLORlZpa99iR+t
CPdxcW1KQeWxttpENejj5vK/06cRcVQWVZEA7R2V8nqVOTDm+CD1D9d5/uB6cHRF
A5sL4+JURORCWZl85yAyJgLlTbEimnoR369jTuqq1lvleYbn7xrD5/jHFt0PNZpB
6cyNLNIh9XWs+fuZH+7Z8jS+C58GTH66eeSCJ70sZBiFFDA3ujpCwp4r3S5BLLou
GWPoEAZmyaXAW6LibYotJQSJrjmAlz5bHlvMPSPV11rIRBjDQ44PFrcTPe2mPu1q
oYlW3td3U8iXsDUptwPMBRf4fgu9NQ4Wd5ByBcQ2NvfXoeYddzGbXCGH709PIk7p
GJQ7yORjcV2VdpTor26N1AceV7Tjz1TMFoezF789/8vuuA8SIFz+jiD4URwaaKjL
ELOszF1yYZ1fkywTD2F3NkiGyyem7428/IUNDWv12He287Rk//hsonOoUfTTTo3W
5/U21V6x9NXerj8THpU526i4+HxBXusLJebb2KOF1UNvoG8rDq4iz2JG1JMFFP/j
ZDXea57KI9OYUSsGCOwWKV4EC6FrIYbSRvW8kHgMItS6KKimwF9UoRnMnhRTif70
9WHVCGvvNOAiHoHjsCsI0+wzFd4zikWjPjMHE195Esc0Y3IbZIoMy2rngZ98VosF
kDrkiKF9Of8ZORWi0+Qv2HLuvB0QmjHoGceQwJCboPr4ehKjmoFvVQH4DojY5krE
vV2EKF3WF9A+fEOVeMD6EWlNHLAOfJd6iiZMbVD0OI0KD0gru5WZfptRts4SJdLx
78AMREpS2qBdpSp0l4Z4+1ySVuWGP1t1aE/hT9HgbSAwEqpvbOl75MCPnE3AUBdV
tqF70OTHdfz6jOmeiJ907VZnrQNqAW6Q/At2WBkIt2+OEqNejTT88osRlWKKZ5lt
c+y6+xPC7N0pXVUUSV1kxOy0gK0qZSA9bB3uW9rfloM3P9ylrfaaJS3SQyW82HFH
0Uvgu8dpgZ9B4557LqtWE7IfEzVkg2BKSsQ9IE4nkpWq2+a5MxbWur9DEgqrwEVc
E6D7NPclLUbu4y4chw7BkXBBzjRQ8noyvQFuzRyeerNwL9ybo6TNSgWYzjRbdD1w
CTbvA9AXYOGU8ZOqMwZTUSRBflIXLSmtJpETOgoJxdBFQwZtW6AohAyCjG9vBecV
UdwulMMgu22ABSli9gmzVlL0qYopx0AazmeqzqHUaXBJtssv24bNGKighxrqcdtD
7kv1O1t2n/21arFLup4q8wYe2r5YG+21jjE1l53VvWxjR+WcCLnOC+KIEnbOC2X0
uAE5uvoTVqkb7d9mecsOTFpX/gn1mTzj6jOVt7WKH69dbT/TBA42mY6XQdeh7NW/
GRGISusCUAHIbC/UChpfNTKWL/9Ddmgk1pOws3VAu7ms2HvaaLBQJo8TmdnR5zw/
w1B3uYRcWa+rFH0adIrduVil5NN3zxUnHgwbPGA/zOifabUto2dyAKRVXTrVSfx8
KK0n7X4DcA+EpnCof56Yz1sl1e8aQhDcsyep303sg6Rvo7iOB6ws3+/YmTqpedpw
rlZFWmbY0bGhKv6cCqZD49ZLBFDH4awI1xCqPAV5oM4FFZZYVerDA3vwAdZ4PnhQ
`protect END_PROTECTED
