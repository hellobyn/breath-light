`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cktUjRqoMgaFR+TAo+jNYYbivIFbvwmRh1+0jsrno33Hi4xOaKO5FNkR+lDvzpVs
R/6M6sREKdWpYMOkna31oAZnA+3LQvi3ZbhEwyAVhJg5g6R3Kzppv22jVGlGK3m8
YaFb/7wggP08+ohgH2e7Dco/kU9nlM//rll2dsJuTKYXsZRdE1Eqb6mJ5izcV5Qi
T3XUH9O2GQ6pumgf/8GH8XcnzAG2VVo+WfAUenmcVL8DDl/juLCc7Y/dehRixpi6
SwjaRJ96hJzUw8+b6RpGv7yKDxO4Ilx8fJCYy8fpl1RtYEkpKaUnv39ghyRXLQp+
jvG7uy0rQgJcNWYveGv5JffIzJX42aU4aaync0U2F/UYaPQo5ReMWORyspoSYXUy
Yu10I1t+rEIOjbZH6Cm+NL/sv70Ui833rpUAHIa/M4jToaKSh+sBH75ZFPEpqIWv
Bia8HX1dsoMxPEAza7r6G6gGLSiwcsfCy/YiMSaKOl5V6fMdM07qqd33RJtHndBA
DaqNNi5KeE+K2rYb9OhZjxbTUKWbCAXFyQVN9/uelWsksWYlXT2t749fnpYffZsc
D9GXP8AwhFGHT/WPgy7NESqD2a6G+zhTUTi8SG+qmRWhdtcug6FPxclag1C6FDIS
2kHfP3FFcx5EMPkkUI1rL2nCsxlWLCNqSsPHFQH2rT44v5JJNLzyfY8xj9jCykQD
rjhXHmRAMxu/ypFJ2sJKoJ0I5Cb3JwI8tPnG24M7h24GcQMPPI/Lwijnjpvrsh6v
55wrkFJ67eR7PbZFFHpRFzFCcaImxzaSAipcnm7YluM5RkCWvBMcDbin4BqNgmi3
6voQveZB7X4jzVOWO+9aVeqgSnMZrFGPxkEBcXStmV2PQ1Zh4e30fcW0IRQCiTxt
gc3FrliTR1w9NQEtGfID7iwRFX7oGXNGoO+iKAQjRksYNCdH4ZUlTIq+EEqDihzK
xizJmtLdjc82+ynpY6xEwQxpWVeGGD5KFUhIzaY/GLx2mOMU5pPyiLsF5mSOWE/0
ABQmI4oIneaM+chGIF5aoh/hge6wHmBUyZyC5Acn/kjK1pVzhL2j6NeNlVJFyDPA
bs6PXhi+ybouwBOYJSG2Td0c9+HhMPpTD5DjaJ+pUaKKsgL1SiEZuiOxbxCWSuUv
ecwkH05uXpDh93F1Pqh5Ye1EL1pb/+84BttegNY8ShLD+t3+MNYkcAwiqHMvZNAA
uoWmibbk6POu/VK4Y0PECOYPrug6hY3vNFwOnSpnaXs5230dkFE0QTWdO4jLDwNQ
WvrGjrpJIAx4y70beuiYuNCvHyX+uePlr0mfPmmDdjsPrpx/FvExN3VboKlYnWV1
CItvYHaP6zyrMUsz5+tsaaADgfyYoI+G9XXoPtWAlNxxtHFDjCzBej4vqgiTOHGv
1CraY16ZxyNbRHnnCwHf5R6m93o2Y8CN0k4+i0uNfl7tuaATN4XTVLeWDCpXjHnj
owlrlzhDUGTNN2vjwDDwmArdCiHW4u96ixuVSFtvVq4AJsL7oGfdOqdK3h+YTnld
O1wWk/RaciPRFfVI6Jld2kuyXv/tYCcyG5YsAJRF688uD72YoMamu48AagsPvhbh
nnjYrRmOU5Yo5W+SbZRYaPMZPY5jFZ43XBe/2+uOCsVXE/ayQ7IdLaA2Y6ihEhiG
CMkvhyQGi6Qd+UT7I7qRaiOxoLw5Wv1wnu+kdA+1CBb6XhFXIw1dIvcgCv40u7bq
dloj77viAhc4byfV9GxqoJCgOb1jf5/rK+bHt1Cv3ByQiGfdIjJ9Yb1UpQQJSzJ8
TQP81PswF9WiMiloEnXeaTxaTNluKwIPFtRKDs5DbpYFG23Z59Eplb88j0mqyptu
wrpaOqkbF6B7uc24+4F1QL3wohIbIJR2/DMR3o/18eMOUaHDOIEhPj8GK1eIEZ2G
qG7CIygphZnCdMFDqLMz5ZPSLlzacbJuYCdGlPoGePI+y80An/FO5AS7ZoouO9d1
4ku6zorknkJ0I2S71AqDnEChtrG5uFs/6LAV/W4r0dOzkZ4Ex3qA7nZYWgXxVcgb
+jfRh5wWrIEOkChXeTumG5Flsxjqz4gsfwnB6EovlYlKsLLuOmtnRC6wqIHXuiUF
HqWfeyoyRz8XtFzTak50LinCY3MhLb57Rzn3HWLlzJSvZmB9IqAGWDj9UBT3kRq/
r+48cXmVSqKHSIrSrw3mbuNkqA0QWrl0uz9Xzs7FkSX0E6P6+26rTRlIJajB24Sx
tI680pkU1a+UqFdSG3fhEt1EL8mf5Z8vsI0yXr7R6eYP9uaJRHLHSLpWFfdCKXSJ
0qXgzJE+y8kuc9dDwBmuCyPCCmju/wiPo5xprA8GWOmHuh88NnKdxaB0L+8WHBO7
mSJnzseWgune3u+PybQjbFxmhi0MrSc5UVI3SHR0sa3+MhPzZsBO6TUUSqLYXEEB
Wr59fVBI6SDwXyEd0xnEu2SM7y6lsnPm/pqA9YagMjS/VYTczn4N3/ldE5uvACsS
newp66gYkZTqibJRiGW+fQMTX6yI8kd2zpscBYTqbUTljbFQW9kUmhUAq2JeLMgv
0nIdpPYdZbGw29O05QYvu7yA73Y7CsmGKE21UeZEzbBByXkXesRNpS5nMKVcBIrj
sHvY4+O4HGRRqzZekEPKrRqOgGxZ4x2XcKhmWve4rkHur8Ls88nVjUHglJ++CKRm
Kn7GbuGs5CdNY7dO+QhAsdHwMQulC+ErrqTKxprqLsJgBJDw7RWcH1xk4Jerv5bs
oPDegDVdxdYp9sFgO7EoFDo0JjFlDb6xOsN5QDOi/7THjzvY8oNrYX1xT/po3YMl
c0OsA+I8LZlwnQ0dGMJR4qOUfOg8BrOcPAxSRBPucJODEuhnMnGLygYk0S7QR5Mp
ZkstAU24wi8n/me2763AOiFm51RV2uqZr95g9kstqh2udRkSCi0pqfniF3qrYkLT
cjvln9d74KOHeStJl4K2FEU5H/LIzOB9K8erMMVr+vPy4X0TJHdOXTWeF/uW35Ln
WtPSUT6j/ryeUJRtnH7NBDxOQlSQfFOlNP6v/XQw/RcThOKllWoeEwlBJ4moHD1R
eC7N60YBSKcO3b2tJB9dBb/YPJBCdOqpaQC9dikY8H7jvdA7iR8KMiTbO3T+cB+Q
DdQVuPE7Xz3o2vWeL+G/InHqi5GhVRZKdAgl29iapwneBFrYiaOr6yiNgoLwZ0k3
jcKtDLpYGC+Ky1KezjINSPGZgW2C+FgOqr+xbA/z92WvR4JtS4LX7p0XGvHCz8CA
ftShN/93bsgaWJHXa0Sg6CjEJxkA0f3Ts2Sv9FcptG472O9GLhiJjn2c19I9/r9E
7L5SANRo1FNecg3iKh2qycdYH1KO0K+DeCjU/UUsj4U=
`protect END_PROTECTED
