`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7/R/CnrYxR/FNBcfmjwx3Tb6yhPN5dnP7ClotAIoVaHaRoTiupNJXHEFzOqhex6
0TR7qQvMeJ/n5aCgP6FfTZEwxpCiiu4p0GDrLbQe3PWOQQtM0PrLJuP2qs9wFwqw
uOk7O3x8Pi0dZu2RJ9QBB7nqcWTo4OYZgB4T5v2UgplQF169td/e220EFKk7blKG
v8CGkVrLyRCQTihbhmdTXiuhtZtbGQzibWuASTJ6Jin1bRv4nhRSNj+CLXCrJh8X
YWUetifalkFJwc823r0eskMfpVDRvxM8zultj3ZJzoBTNg4N9ZTJARKIfUmuUW0R
18thEw8EMxdB5R4z7p8Ff89x3yYj273+Hv4fwRzdYFADgmrWY9ddsd9OV7IjCO+D
iOUALQdMOw6cbpquXFQE6/rE24E2Gr6uVY6GanFX9ZHFhygJFRGsT7jxjxHRpIyd
/Qg6LfLx8uxmoXLwu+qIojW7UZn+QUx/lp9s0W+MYIS9X+VrPbdj0F8DqlsfJRHd
eT8yMvZHKbrBg+KFGXCfGE06PSgz4FexyIdZS0+gytkc/P8+aLoNaPvlZ3xAC0OH
iV0gETBtwHmgBIN1A3rUGMU13cEEeQswl/DLIhuXfcY1nTvM8EvP+KE1KvnQJFOX
R/N9vHN4tKoo3ecbRQh0IOYGdkmXMfJMMIghO/dZ9bSMjksZuEW7rrKbAzkQ84wP
j2nP6uErur+3KQ3Os/EKgm6WWW73TGwaoB20qCmwc8Jbi1dczgfvI4uzqcDdrgLb
ZwkS3biGyTbq8amP8YEQ/mHBnOEDmfKEqmABVRpRf1CpO4D2TLMMuaL/DTdgQmN8
Um74kuoYY4JEW1AOOGCim4GjA41Eb4VPbaIIIduCjPPlYHqFWYht3uh/R8t23tLM
0LD6Mj2nZG7TbtIwwLT1aumgrJmKsFEfz3KTIYLJggJOSMpPWs8Uzn8sy8LzMazY
Yr0fp3ZBlu7WmCnqU3JzfKIhw1EDANiydxSXFv4CXEhxJZnNLWan0bnrFNxwHwJm
eiKkAoHSGhHyPxJB91S14Dcf4zGR0AGpGIXbqtVtSIDc4Y+gIvYVbswQwv8WE9q6
usDRxttmyyHhCwjlQ+GkrHuoDuTrrF/uWUg+m/UR8pTFMpsnaWaNqB07esa30vLq
k2jiTtHGfhFMP4zpkjQfkdjl6ufZJ0qR8jZdd4ZZUbC/17b27YPB3rhxqVMd/r4S
Xf0/feGIVUU5aUR93prErpry/ErXfSQIZ9rGg9wqkfXgTWbowCRknQWl77L08Hp8
rlrZlq42dmrGHEbMHo4gaaBbD5FYgyDKRU9Zg4wOGjPRF00+z5nnulaaIsHHAg1Z
wEABuzUr1uvKHA+tYV7QT1Qs5AWv1Z1w/eYY1HthjI1JkZwU5wtjHJsCYkv6wXUZ
0pFRKvc564vpDbKmHuid+mA6bcgOnZID3dcbPpKdMvG8kRx5oNurRe0Ep6Z16zUu
1oIwQUC/ozPsxti6lF4Zq83SppUdsKHarHZs+iRCJhOrG908Hy+dd/RFXhdyltSr
Osnb9FHflz7qEeKhHfFlIDEFrqlx7pTErwIW3GZM/h+/Kc5fK/TP8puXhtn2ubXe
m4BURuH4KV70Shm3/x5BBhQo+GFq1g+34q64jbX39QJ5G66VDKeUX99Phz/+jzCo
cMoc2ESi/1AiyuEwubGAiCPWcOZrJUIciZzUd5fleEccHVVWeDfFyMm+9J2c3LR3
dFUozGslsiqt0XGv1jKJB2xOSk8oK5buZiIi07W6hUd6gPlHSj2W8vQlgcfMP2yr
qBiYJ+kR5wnq1HUC2zjGTTRKs6sm7d2jLydut2bBplX6uXVZR7oWGeeDnlsgE/Fr
RcZeZO/lFECS5XZGrT6reWStf8JAkQBwiQQCxSyh+WWyDui6dAn8X6ZzhiFj65SZ
yZ9t9s5TPG8QHqNTEUrhzYDAceNiYB2Y2fiC8MsgabIdbX41d596yd0RUi91t4Ij
JNozETWFZVf/8kgif/iQGWST8ofrTb3OZoN9DMWduDwwQcgA55rE3fJIPXagWpaA
EfCNjPXamEvO2RFrLltN7LidNdc9NP+/rwcKmzpx/R9rmOe+18upBi33l00ckQjF
Gu1agyKntUaRcMPynw2H1i9Pz6Ac81ycKgGbygNOXHbOeMKImAUWotXnZ/+t0g4w
lmXuwiSf4CzW6XAoJjEPU5VodvXJLmCk+axxo+hEoFkRRHv+VThrvAin7+tasWae
VdKKphoQUwr8zQTNdP9nBAAYMcZJzZfNoKba728ZG+hON6zbIEtwCbb0gj8o5vj4
YChMsH6fjTRqtipbHHBc26C/nYbRuRbQkhaD0DCY7N81Z+lRpUR03XlYRdM+mjNx
IX4NuZaLN4J64KBqdIhov/yH0hVSumUscSw8Qk9oGBfidr+IO2yA06iyq/Z5dO3Q
G/vMT671AkbxDVq4FD61moB3xTXa3veZNJ2BvVvGxNyW2uIl+T46Eru2AOvqPoix
qBY05p7H3b4B/E4IGC87NQT/XeEdd0I6WuHYyDDTheuiY7VHl/iCLlyVy8SdTyQX
H9nIn1hD8WV7WyEoVV3qdg==
`protect END_PROTECTED
