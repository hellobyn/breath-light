`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEHW5kVLSg6hFSanYll0r7VGzUxHeKWERYERcBtlleysmXprNfAUQkAa1x19qRjS
Yv84M5Yz4FJWMgNvba5KqWCiNB/h6r7Y8/P4LsRxYjFtfkwMrEupFO2N5XIpZUyC
JwQ4DKb4ykE3ygWmzf1bzAs+3WP39XfklSOrCQySXBF0Ji8SkxOUQyUJSG7invSm
VtCEGf0qMb1Vmn1KlddC+AkdhlefvQZdMJ7SCoxW0JnwGNRYFOh9QPv6Kfw8fNh6
xZvqxAZLJLZgVNaOIZ+XUYs8N2HKN+p4d0lGfZN+0ePgIpXW3eOnYcR50QnCN1Xb
EzninA5CBsGY2h9Wd3pVyhJeNoj+Lb0UkSo0l3s13hNr1zaJwNO+odcZ1KEtoqnb
CP9xX1FA+/YSciOl/jYXkG68PU+3ugLbEJkqqmFa3ILX9LjP+Jv6nEm+M/eIgEpH
P8lSY4jw5Nke4jygQsx6RaowvJihTpP8lmn32VNa7cwDQ8pXTVorGev28OJnr6/3
6kVsUU7exevadMFZL7OWtzvc2SNOo6aJMEwFXmc24SMyXflpQKt49ND1MTUJ0AWd
C4WspYKysD7k98+Fj+gKaFMl2YUuENAioOg6q88n4W4GNMVwpkcQuRZDU97EimQY
gnu/SnpeFem9RnwDRs3vCAFnuAlak3hahojRQzfuREhGdr3uYUMU7+okm0qig/S+
Y+0HdHNALO0d8NbT4XOl+3k3ND83at7SxFtmE8DGqRJBxaOCKso2sHRudJZ8LWuI
k1tiylZGgU+e83YJmJ/Oyq/taCFt9LhxBCw8SHUWMN+pTnV6Nd4vWsAGwFGakeUI
AMTIHp8uipETcIaiOBXBsqfXWfsaPdA1oO2CtSMW5Ngce7cDCIRTmDTj9v8DY3Ou
1V5hi5VOIygp9IxEGQQU9YHfwrAf0khoNIOqmyxv3eYUPYyZUv1LiUb30AoVbGB/
pcwo9qHeh2NqTsXeoVFpglXy4rmJaLqMXUy66FUbgoOqDrrNT9WCM5qmUq3nAGhj
gg+hvdUKqpetRHQLDvcPzjyFWmiFEsIOA2TgxABvbfS5ccSHSWqhbXeK65PzSCtg
CWfGVexdOQegJhZamRxCjQ==
`protect END_PROTECTED
