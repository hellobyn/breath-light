`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCfSv6VpYsvNJlCN7IZHr7KkRpwb8xTEO6MmefVDMjCJmnmiymGXiIfxNr0ip6xg
nkgR1AOwLIxX5tNKPdAzw7BYddT3S69Z7zSiCzuPs/EryT4uArndiytBzddFtCfo
22Koif7Hx4E8Zae6peT/YztFh9I+xhxBLMXLZPQY/rLmbLEao+ksh4VnwarJWKHg
J3EgkTd8V9WlyvCbEuhCsDUkf36fZPtT51Eu+6vlmuFhRy04+0vWlgNSVXWUbKHv
7gCZZjqhPFp+MQeZnC3yvz48YVmhx4jb+1wo4tOMCIVRsXLkBYVVVCJJpl5475qu
n7F0e9il7iuznRbcB+OPCeur1O0KbCb3sof5tM1odwCeD/42aIiAFiahgO4VBqry
LU1kIxCMyakDktUbcLhS49Cq4yoGrpR+yG1ySHXN20MIH+nIaXT7//AdsdGZDO8T
frqbGitgYsGAq71M4u/Hds9tqo4FqxZeM6J+lpTmE8qmx/m8ljvrmGgGp0vDap9Y
gcCmW9OAbee14pzDo1+QP0kSnotH4mO/zGZBo8JGkjNehLcTl5m3DAgYzoFHYCXy
O8RrmR7epIaoz1bs79mvdl7sHcz7CXkLIHVcV/0ZuS8VYx0FEa8oINn1pNnpwM30
KFWzzDVkXN7iLNtFvhz7NX5iiz9OK3Toi1ofPVHXwjg/Ohzs57FpwThIvYNT+zft
6erFW1MTqClLpZzf6MvTmuGwgwSciB78ZjwiK4gYPhYrZtbWl9f/+rjZ1ATmZjHv
PSMLfgM2g9aXBGcC+4jaOevdkuZtvRK8j2bBzIZCYWDycdqsuG6L/dl0z3RfBUeX
8lg3IQq2lhVVazs3VxqsygKTuVL7lKik5HTIB6HRDKvlj+1xYJNQg2m1XLaZXjWq
POrKPGgXhUb9G5fWEgZYRitKFX8WAHW5ChvKakj9y/LXEVWCD9poOUvXvs0wd9mW
12czR8Doo0xQAl/onSVs47uoV7FPqExAEK7Ob4Ovz9fJtn7LzhNKE3jVJsA9csB6
HfFKS2rs1I0RK2puRARrUe+FpioRYgkHYjSPUYYyJ202BJ0rUknsF306TwSxCd8s
d2U4lb9gbG0+vLeXSG88MAb2cUnifL+0ilTNFL17JIWpMHXsBgrC/EdVGKD43wcI
LnbVtQTq6aPhT9iWkkgOaDQCm0H3OuaZz96QJRBP2K15S52ghWqGUw8+hhcwC1Ke
hgAMmrOxzNhAyZ2DmVL0ojEQPWtf+bS+Gj6/+TH7Nf5K5oZtSZXixjrukWhWMdgT
OF+TQx8k1sMh+RiHsj8v6fSyU+AvMN8OFLxxNzpoQ+ipABqx9fIQD7wpDCOvUzh3
fZubhsa2VZ9rEooNQv/ChPJ0ZoHfW/ZgH9ML+D/CVDpS8J3nuJCwV0ZmAdzD9AJl
2j248adz9kZp+1fPPDAT5o4ARTWRMvVD0ao2OJpFPysWuj1G0GN3EjQQb54Z5jRi
tyPLqkKdGtzaf/xGTBB/PV9nPX92hjxiOuk+OfAmx0py/8EkodbkpeOh+re5lyQA
UJlFdrLDtUSQssHconzAsxgUPybtXXnTQZ3HR97PWSgUCDZMRB23hw1ujmOkzDaN
4+5QbKS9KQliqmR/W4S1q02M0zbQk/jV+0hEEZxxXeSjBOlrl5HJuSw10CtyG1Oc
FsoHye4ETnh/xrn7dQtVWd5NjUSLLMpK95oXiHOHhKKF84hMOIj8X4HTwWPQ3sXx
8aLE5OSSKhaSgOpBgvkeLCoxFzLE+OenzuMubbEIoJrVB0F78sVLvpEQqM15+pnv
lc5ZeuvPyFNvTHWSQw2xoEqRhUNF+E7PqNJ4RhJFJMNz2RQLExMhD9zdhP9tncNZ
n+redSL8Z9r4gjk5ybF6RocZq5v/Z3jtojPwFO/8nr/xWB+zzh2d+yZrYCMhRRyX
Nn4/UGjIJUPPcO3W51HodFewDLMwF2/j62eU5qe9RhhlMhH5aFmeb2N4/Qxi45fu
WP7tLy8BJynWp/hI4B+xUjl4IBUygNOC08aUJf2SYkOQ6zFqp4sCO8Iyaqx3YvPB
Soc+/sHWtrzm5jBRZVJx1IrTJVD8bYmGv/BwpL4/v9eS0H5hthfzGn24BUtQLX/d
pEzhocVbafet0ar2TKKdCQrZFQmSs8MwCmS/dEwsJgmdn3LgJhY4SHmaz9Dcmw22
FHvjRjBNsREjSeDp5h2u5YbdkWeoGu4fyM4kSAtpa+IoJk8QnvV2oUfFaHPSXHIa
/H38/JUL2QyHvBIWa9p492rENs3E1o7uq5UMJIUyFl/j5Fb6JbzA1Cy3L6sBgwRe
TzwPPcvD5PahC+KAN2V2bUY340zzNPJWg/ZFcWQ1iRZ1Mh77+vGeNepRUYeHMQRQ
mwYLZveJsjzsHI2+DiiT4ySkJE8UqihGq1QE94Jv0ae6F7i9gnFfbQ53Lb8ARAW8
dw5LY+RTGkc/tzOORLBRiINpf/3fkvYzSDYQvq3bfIWOdZS4lwI/qXa0/nMCaI3n
DIxvW7B3yIPSbbqmy7K04GbJnRZeBzt8GRjibhRZeH3/rFHblmJOKL64cr3q6uxG
XQqsna/fohFUjrzOtzszURbz91tkm1+CkTqoqYpBvA8+Zp40tuwUTVs40AjeWSrX
VNNuJWoCMZ28x/UluLkBzDnn8R+8AsCa8m9NuDK+zrpG+CTThgl2vnxU47kNEFrv
qAoTHLceMiZeSOsMHZV0IU+lm839tOKuiER6Ad1WmvE3r0FzkYFt9jgKwGYmxGKC
+pnxM/Y9n3qnwbQAM9yAoty+Ghur/XfwCUvHa7NF8Gb+hnD3LfON/vEIilhNCkO2
BXrMCHiotu1468JilqXDLVeF2+lwvJtLOxRxZWqMIZMQr6XeHkW+QLicgTDPFbDR
HZFU1Um3uYVKAEEdWw2UD4TOMP4V/93XoSgPDFjr+U0vxXRkMDrCzeThfBwKnxhq
Jn1oJp9PeOcti5HoEa4eYa8aDH8Os8GBrV/O8ArpVs36/Puq4oVcqZx5Fe9RETSi
HavXCGzA5TZ/QVTfQYdB5q5TrK+1IAuvu3LnMlxCTwjV2oRKSsF5jaHR5aw8sRAX
zuHoqPNmd4eDQgFQrcPgyVH9yC4JmfsJ401dZtVHmBobV97Cfec6iIXUgycJFBxa
xKo0zr4CZUPmx+U+sENO1nFQC9EDqkN5KkTeq5o+d9OEl1t9Y9W1FtBFIbwPdLxJ
j/qKlGJpfZtwjiHh7ENVO5n0AI7RmIegFMmGns7I5Rev9s6M4gCGKfvLh2a75qfh
BjZaG8NidwOQ/ZjOznc3FGT6op+mqEqaBacCYe28XFJaVfkJGHwQnOhHeSqxyEm/
Cc45Ge/0/ePJcu8RLBorsCUnsjuKQ02Go4ueHlv84xpUCoEP/t8XSuuDYMtrYRgc
ntazNGu6/B3D2CXkI11HVvtIyOJ7sHj35iVKcI7dWPLye24FnXz3szrlSQq6sTaL
gtFJtCh+nHYeRtr0JFUIm6+EgN80eYDuePIVgXo7qSGMwP1IZ2RqrPSwXrrVgwWo
9EiNE1mRv9Erw/Zhqk8lKjb4vzJl6/bMwPSuY7s0Qj7KM3ghXm/M/vogOHKTvgY9
j0/HqNWuTQ1doEBBp2qtPLLb6iXuAFFCNrqG6Zt6YzXSCFYOIsXc6fF5mzPPVuTx
Jd8bhum/yjWGaMbUvsVKRnHJ4cDb0dUhqKNtPkngZKha6pUjKnHz6gDxhCeMdfLT
h+j4uK9kZO0Rc5rW1kLiUy8UmGdj1QnyLKiafgIYMEU/l6UV2y9lIplI4vHM19E6
9YyesiSotVnlrTqFyCCQ3j24h//40HH0+rkxSvRMmlI2O6JdrzLTpsod0f7Z4smV
h4keTTf/0hOdVdsnkjkdbbmCVum3JsRTcL+jPZB7oGhaWVNNOyxQeirAaxePa7nI
aKPPADcdLvxl+fZ8jOvODowC4KPmw83iZZ8UExv07sMW2ATx54cbg79bu0dpFEns
te8gjd/MbpC6dwFPVY+IXa8PmATTpqag05r9ZFmxibFoEHunoPaV/ZrLgEb/Pouq
aRFaTLjvDqwSxi6CbUslWxLGN08gfI0B+H9D+PWtw62FOicHWmYqzNQk0bw6D0bC
K3SNGLRTkD6SOa8bLe2YNhLakZzwBB4U07NR/j98jGFL1F6KMfxUwy2SCMJNgtOT
71AiIWc7t/Ch9EdIKzDrxiRNPf2xqB4OOCscPwuQEJ38z4fzgNLGEkBRZs5qLTmb
16WG3P6wGftN4eSRRqC0nxhG3UgOtvoFoQjS3wqeBncQhyggl0/J3fJr/StUf/j0
5lDNUJQf+/IJhffkEHJw5ZDWtdipBzcUDRUnPwiOVpqsq9h0Mh9Ab6SEa1Qki7vw
n9hG6jZVyTcomFwDqIZh3okLtaMYm9PApkoLsZIdoaTcqyJ5HhiQ5yCVHJssFJEB
IqKSInK7FQDIdhtHBmIQhCYezf/eghYLzxGW8X89f4kUkrxeORHoNNvZ9Pm66xS/
ZfgTWMJn4+AXwxb0XOwc57HkdH6Rilnf+52F7st7X62DwQ+dI2ompDLGiNwrWXou
yYyDqYUsCjdwWNgARohs88Q6rujNHuojMQeh3E0/nzGZ7010mrxvY70jxP1qUyUz
WUjpN9YxP0HJ/fvyYlpk3fEb2y8FU1WPnB2tJnY7ykQRgSXFJfEdRWc/Y8x0vDJ7
Rk6plmZfuIguN4nfSI54dL0b6WbSkOYuczDGXRxbXRK9RP1pS1D7vCpORm57qUNE
Kl1NARytQBYDwkKas3WOtSvyfsSMNgN11+YUTe+WY1ORW4n3CdTWUO5rQr18ef+Z
eY42yPAJ2iCaF+fT6LAGQY3+x37eDG1nbE22d9BgprJpE6jgUHnRJt/WGz2D2Kll
rm2d5BQnrA6hxZJdX10iNfDsbiG5JgcPQcJljTxt5ERxVyk8YJiV69ApwaKx3lde
Jmx6FPKpDUUh4N8qxafQVApQLr2pBQ0crJPHhxZhhOIjJoUZmob/U37u8zT31F4n
4BHjGbEGrzz22Q8Xmi1rsxJzgsw7Rg2MyFWeQ+qy2Q1IBRQv4qVmaAkEblPLI2MX
GKUNOsx5dQDhFdyRbWgU4l0H0gIjMLQRrEb1Kp9a/kc7XfcR5Y6WnP3Z/wpiLg4T
buAGE2lorHWxhjzcBCzn/08ah0oqZogkmTx4z504hGvTjVn6UvNUAuAOJ1IMZyfN
bzCl2/eGLjIkKIB23sMcxrzzYhT708T8v4yaO2PIYMslmILcLhEem5C5IioqfABO
dnbZDq56smj9owrQDm4aCwWk4Rh3xYC2fyfF77I1nKgAkN5zn4VLUAArEyn8dBp+
n06bcE+0eN7SIRlsN5Js+G1q6EfSwSUcv9o5+PlcPIfRail+UNJZIsejTklDj3y/
HzEoawPgt40hd8l19S8nClu1lB7VIToeDEGXTRAhtAaEaFI8xAXtSIRIhY0aR8W+
dDjY8WiodwH09Z1cm0HErR+iNCKQsB2YIS+ZnISY3d4XCCgxsLlE/gCXjh7GaEiv
tGnHWu790mLbHjEeD0hqw+NlPNnSMzUXKJWpbsg39PNLOk7htSU4XgXL0wSIMmxb
nWlYHDnREGtWj6gLrmZxiMa8aKeNaa1HJE5RHN+LJMDocptQuEFMyj9rGlDNHg8k
kfqqPeHvAmsJYKv0p3LYi+ZOvUsC3nOHDndclB/9uG/4LpzcxbvplPoy7ADh3giA
59U+I8EMlRAm6Al4mbaEypkkabsWCznpJeVhstHWcvUmg/ii+reaso2we4WEuItk
CSkr4GVWwYaUgALh3A1KpyXb1jE7r3gysl4bjt2Oj0tLlezH3qHxvryutzkPzszy
aGWQ5Vdu8xZlL3dRk3HgXJMok4n/m/MGM7MlKckpKpAh1iquvaIgZsYQeRMs455f
31TMu1Wh1Up1dxFbnkkKBZrg5UcXc/5PzG3YtqKWJALmXQ3DQ2VNV4uCLetP1Vdt
ah3jQQdkQ1o6v/f8Lsr7ZajO0SoVW4mohvS5pyfiKFM=
`protect END_PROTECTED
