`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNMpkeGsqd0rx6XfHdkGY8+rgqeDGaglM4WVi++oxosL9wJp99GfQvrOgxPFEUBz
/mrQ7yKWsPW38J3QnjC6wgdq6jEP76dNCr2A7kmOZncLVZoMpj6aMj0AKXfPRfY/
mTLRL78icEvh4tSu+nWl3ciqwWMQS5jkc9H5lYEXq5VpsgEZcC7Y24DNJ0PRkqTw
XdDbi3b0cuDH3deJekfmH36JZCQU5Sln7LeKEny2yfH/8CwNTQn1jlbJj1zDweOr
jrltVIE6GA4wehqMZmhhyhqu4QgHvWRvn8lIA2J1AN2cPhpEEHwHzcBdBAUkGyNc
ZAVl9qz4UwuoJoka/xb12OaKTG2Im5nfM5yYMTUTxuUwMkbIflATqm/qLJ24T9uh
MRLbpi7Xewdg2M0E2KW/LH5O1kEKPNHZ0GKEkBI7Rr73uEc1jimfD+T0QBFnZ5zu
+XvYFcGwYsjhBLC09nHPWkSul71+/xa1gLG/wZGDcO1tIzemGW9fen2qe/zEJ9Q6
ZLI6+TMaIC5oj4JUqUjyNrtfM+GMXddHSYaWIVItEtgdt0PBXbhDulwhgwZlyxE9
FTHEfldIjSs3xFlIS7RzY+aBfn68NTmKpneVtxGp1YdJRR/lUkPrwqMyi+pb6MHB
Lkb9ABhH32OPymKXLSsOfnDgLyZW/J064T50wuqwT45ynxjgY9cFiVD+NNXdCJVA
uXdZhZIjnO8I7LQXa6UUi9ku9mXSdRvjYbc59xlRajFpnBjVmjPVycmQRrrf0iDi
3FZSZ6dmsprar32eOVzU0vy6P6Vg/3Ut19KB6DO8vaNcEJVbi33PIFLiLTCS5Qe4
ndrq+o0dYIGQjKX0UXf2b/BHxJX7vdHyLMo/vx9KA/pESL4H9NxG2Yk21XFS3hdW
93JqcpMUfwpfV9S43QshHLWwnmqnV9kxq3kLn9WGnTeomUh/ljiELzsfSOxdS9Mv
gqpQfiFnETl8GRtZAWLGAqyushmWliyMO+Iq59KeZu7aAQ6KoI+3rph+ZO3Vyzst
QRlY+8Hz+wEL4FJFgSZLi9RQRF6oZJ/dnSoyhtixtA4IMIwcJg5+7wA4WLU4Xhop
ChQAw2Uq+Z2m+QLIIWVWX1Neu3ZuK6n8VgBtMeIWjkD6SSWqe19gjhHHR4jbrTdo
sV1i279hjDPWS2N7GwvYp9HqZo8LTtd1my3mrm2jttk2ziU3DFTI24QGLY5UzQBb
UUy3/X5FQeeywRSYr0SlKQ==
`protect END_PROTECTED
