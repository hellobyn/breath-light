`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIXE8v5mRjMSDry6pHKMqRJJ++oxTm7Qzkv8gSzx5RqXBYwoCbl8q/mlR2KdsOnG
Wjkr44xnpDXLCnN1iw5Uh5D5HswS1EWnIIoT5aS8TbzkgYYcFC7n5YCl0lMrlgeZ
qdkdcmrtqsBns1CsSK1bolrIKqgYs9zfpFpZgYhWP1o6x4NdINcuhADcBc/Yuhgp
hl3ri1ML2zFT9tpOJL8eW+Wbyjg3Fl4B9Nc2uJkZyX9XV3XcLhwRTrHQnGoITvbU
4ga8O8b3IdlQUaZ8fCnYjDtonMCNnOUBY4Am1COtzsm50WqTCwHKBn3r2qj1ha1l
DgXibUbobZOw82aILGrk2VcEqMQl8pEn9JdgpH2jOtaBztDmlnHpUFs06V4h7W47
rhW1J8PSRpxTHuNV8uFSKAfQ5C3jou/NWKw0zaK8X/rkcEnu+M9qNSzbiMAtlmmS
FUzvAncGbjF7j1nhI9DmZslBZFPdRoKIhbfFm1HQQDcGjjn/PFxFdbi1YWCRAKI3
8aN7wKvasBRoWmALDwycYyufnH+Z1m0VbQWgqM4VCwywYEd3KwksabpFz7faFqPJ
8qKfAgpP5TfVKydQVcLrqw==
`protect END_PROTECTED
