`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfl3zShaOQPhobLz5vqY1/Dnq5mKwWd50OFD8DhrB51UDS1QzQKtGekgd0p+r0AQ
wM+jt/n5pTgAxvXJqXqY8COYjkENPeIIBhwVQYrJPSAMr/CTI14+fihMD8DvqTeb
rxUjCnTn3w4RqUyR5BhStQzjZMAlTHJo2SQZQV5SSd/xtDC5ZCpZ7F6+NVSwYsGR
HE8nH5IpF3a3hdR6RhPlMGTJEbGdho3e2hff6osbMsldoTaXNRwnBPLXKXCLhJB9
v1rlH/8ggcjsjk/9JCtGauRSBREDbGEouqNoqYequUiqA9nVZ/aqQa0CgMbQZoeZ
vbUpd+pt177pm6fF0h/9H8RU5rs1QGCxT6hG7emI38egGSgXAHlQjghWVpNlecBl
4XYibO3YUuC5hIvgMM/P8cUmY8GtTjA43j/WQiMzywvm7PbaWmSUdAeHhVA/K9xd
G+YBmdOyfDZdVWmUpPbTM6q30VDgGc18xtE5J5Jnob+E6/Z0hgwSAzhb5J8TJUoO
wHIMPWPG5cGpr22/NdJtR952ZdfYgyF8XRecTeKps0AO77ZzjlcF3bRpRQQVPXwS
ERJEYDgg+Vtp+yomVsaSYKVGt10ykvCE7DNxlD07L4RKyzG7nf6lMme8Yd0UQaG4
EPgUnOe0fEhvw7VSn2ZitvaJdskO7c6KZb77eUMf9fwIH6/2sX7HTpVhSWNvuQap
rrD8dyM1+9x4BAb+e454aeyzvg1PaWeeUWVWkHnDBv0bgWABtenJBOXrqIyOcGBr
MqSw+RvejQ55glmrDdZ0oszwLyJ2xbPtHBb+CSufHfyY+CWy+VHlEPxCRJr5qTBR
lYDrpfb7gTCFc3tFR7fEAVuSDsFHveeltnN19wMRAvfV2E+fe6lAlMAcLsfC+CwM
yqYRNk5BzKxqpErhHbfMehzoMNelPCQtxUg2zlv0tkn6q54pP/U3KiHOkWFXXsZz
`protect END_PROTECTED
