`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHVJr46Ei4jCggj1mUY0B8VAimgUZb1X7XaeDBnIeAjsHoj9DXuT2gw9XkBh0Cy+
T7Cm/u6xZ8Yr8UHHgotyg4v9WBBl/Jc7ZJyxKdZruBJXmfcQtrY8GraFItaGgljR
ybyzAB4GXUdwnjnf12TXXb5POIlzv1pl9IgL2vnDflBWW8UcQYBjNxHdmpO2Eb7d
4ya9y90+bxxyHIguzUC4clXB7dDp5PD8ow1gfJdmzFZyNE2YnLLDaRuETSxy0HnN
i9yLAaHPpExQ+YtL4fNBRxfzShnHD7AnRtTCwnyWPCqkCTOPxRmz1IAP3YV807Bm
gGOzl6pmKjeCgOVmQlXWAesM+kHNlxaVwN9qpPHECO2kEDdn0fTf4WqsVGz0DZcm
FvkzMrkztst50+OXlCA68TgRhaMUN/cV26say9xa24dvgU39553V/8Vs8gf+2hrw
P8f54KDVmLF1doPXijVH9sLnSqn/8r3f6HvTjxQmPtKoWNZlBQeTkeFTyIL33M95
Rf8QI0ResJO3cef4gLl4BtRW9IjU/skSt0YhXfGy6/WGPqHiYoGI77G5FEcsnFvF
IUMOcBNbR3IYBaqgKpMVZ/zi8zMWWeUk3S8HnwmYpcjOYOcrLH5gVjN7+hK0YuTE
QIZOokwbG4Y3b2UhU9k461b9OV7dvdSAuH1AjyfZxq99kqiKlQTnrA8OsC6XcI6m
BfpPPua0L/yLPofpEZi8rEc3VjhA8sxLDUJzKwupMS7G3w3phR8WuAFUfk041cW1
jJi6z9z5X5Jo4j/iWF/zbfAFiwvMnZ0gdVFdGRsrwKSAkUGRMQXZCBl+PzesTUTG
0pi3tAcxCOWNFgiBW3DMsBAmnnVpJi1Iu6VrpSzGYig+0nrU4DE8WJYY7zHpgMiK
S3TX+587hhZSoC14G52lTyu8UvvqGp9ukTfZS+LvjUbF8v3yqohN4BdUgEpzaFVA
U3IJMA+5fgxvmN5KJQUOfshLqfD4vtiz5KDgouGGkxyWlvacGZN6oGgDAd2Yo+Qi
vOcqJXQahRlKhbngAg7j6RUHBnMl4QlvSCx6mm99qply62cYWHjRYOOrKCtGuSCf
yOV7pMEFtB/acZ9RNIWkhsJ17QkQm5ZUVw53MYpUN6TZPvFiaTSp53UNEtjWtSuc
vV/U0bETfRIilftqZhAbh8XFyr1QBrizCthPE7ghG4mJU4lTEvxy/SFdBunoCeTT
90LpbZDrz9F2odnunEvdcVUNHe33Y6s06MgJLK5AMbP2/UJzscd6Ude7EV4RpWOs
SfHjcHjQTpDGZzA48iVXEsXUXdBev6ElVTKooifjKlQFGw6iWSKaq9i1vT9dTbNx
0ao9o5orq4NBKfbmWoE7eBr0K5rQruRJvELbbGm7rRknb5y4zoUd9J2UPlS5YVvg
OrbcjXTGxR9D6tB7wnzpV1n8U34E3fojAQoQ2xDRAexXUxo6v96bk5hDTk+B3Tp+
Rz1ZVKe0L0kgTWlsFurUv1truu9TAR38WxaZhe1kPSn8TTskD8TICDcdfBqDMmmc
5J9F/Mxo+Y0lW5t4Pc+oxyy8la51eu4RN8lDxXl9EpQgxmmUSZNnpPWyYfCIg8PO
AHRTfvYlVPe+vtCASqIP7KFl1xTSINbdcYK06EohrQ1M/cFzoYewAUwR0uFcC2YS
/35rXBqHXH1N6wHUf5/eyA2VcFwG2YcLYVfjhMN1o6kOLnia26Xj0sPeUAxuS64c
9t4lBWGRLQWBYYR0XVnIzJfYhr93qfnOjRmmNxw4eje4lyp7e06atZOZSok79+CU
ZHboXv0hqIVvMBTj577d+2giDTODnvkQi6JiuOuaVQxiKqZpZS7NM7LWoktQ7N/s
mI/jljFQmd7JlBYdgtjO/WcNeTnmQ/R8fqFzRA+QmGVU78Ecq4ytbzr/u/hmQlWc
LCj/pjMSv+TfLvp4RMRUX/Kwn33pmYiHBQqYtJkgmYBh4HDfhUeHGiQpfxhBU4ok
e1i89zoOQ/PLmyM2oDl7Ij691EE1InqnQDtooJrBMNe7JBQIiNmngfBq06oCRGR1
YVC5KHOE53VWZgncEZAJHX6lBYAQ4cFEpwv3/JqP54OlB6NdbZQh6Hduq5EmexTJ
sHGDRILhTwH/vX+43RsSXY2x3InzPtFcWLt57Wp8ggtFlVNnnELm9C49E6Z3X2zE
ezIAQSUlx/ezbaO6tyvDSAcMLhYxEMBS55yr/XbFK/6TBnY5hrFNDEcE9UXwmAqM
2FllA8nkxHQ/hwgVf6p3UQH/sQSV+oKc4m9ou3NgaDgZ/b9hdx0q/GkpMOhvccC3
CNSQ/BQocLj6GhmKO6XpjStcbjGxgyomvg/MkJdrHPI+0YwMWNTa6hCxk046WgzA
c5bk9l5gCGytAg0ZzA95rYfdqC61qQ7skGXdoZ75K0TlKS4kgA2b5VlRPC/YV6Cm
p9XwLTTZBEtEseszuO1lOjI2xnDHQeuq9MYyGZMWXJKvoBIxtCRFf+lRuRpwDtqq
t33LV8BtMunpmlyTOF6bBamv1Uko9EHImRgapBe/NyLn5hXOktdV8YcYnvjzu68i
R6OpfuVrBK8gRhM4pcbpNruBAw7AT2P1ETDB9cp9UpdbMwzspqDedZKCIlffBfSQ
OC4h2C3ZObyLhFBaxvu0GS/VRMR/ntbg9JhUmaNO1f3JGK0HxceJFdz5JqxNTw82
5e2SEl+5SKAHg+4c0tIKdAuVqAYVS3O0EmXUatqtbkpI/42OssJIuQEJgdyPBOik
wN8ZsMzc00IypjPNP96b0okiqrN3WDnzRh3TaooT2yn8z2tIQd3sAJe2PozKvEya
JIBg8u5pjyU6lQqDt6Tb/qXgxmNT/lCrobuErosqZK053A1jff91xUeb+1qr+/h/
hb7ZrHsQNbmrBKJ7c0FcZQgdwE5Nt6F0nM07+e6WlgxOOl9Pl+yXQubpIV26Gj3J
o5B5qVKlxcx58xXESDo7fgef/Tg1tpVicOxAoYizgoyt5mnHesVZx8fIt7dIDaOG
tcrgK/MK4KKvs8EfT+99zVaEzuVIC7Df5gCecCf41EcStLVRtROOLzmIBIycs3G3
hHarZKE9eca/pUOfxnaf4aO1tCtmjDHsRpvEsP8HLYMEebR4kYexz3zz0T0J015i
HMb6vJPnkNzULombGX0QJdmmb1JmeKh4TFoaLKHw5R04yMrwkfLYAzv5gYTjIDPi
XxsomvK0YJOwfcpSyHENZzIR55CSkIYWPPF2+GSRGCrjVUhQssrINTnUu2gLuOiP
v7/vugUPQNxmcVscKmLWxgNjwVXCPw5ZL3vH54nHh2PcdJM8+QpVOsyIZK5cJu3m
brbbY1B0+CtLR493uc59zNy1VM4pAk0g1z4r+WjZBbmMT4Ra8uZEbVbUgFNU7SdN
E/qRbRFR781LzRj39259xrttv2q0XJ+ghoO7FdBwCcpsYnr33TtcpF/zNPbebZMe
ZyqZo8as0Z0C61aswQfbSpT8ybkGp1TlkM1Wkqz+B6zc13zUfvYSXjkPDlaOgDA9
M11F84KKHJ1K1pOeNMmcnB+vWydbJLrSvEGFZXtxn2e1jax/yerCiWYeoLLvH/xm
DXaoWTbJEc0RtxDco0h5UAcXu48ItuR5OCaKwyLSaHJztUxCW6EpZ33J698M3g2w
TSvrbyO2TrTzbOV6jbjSrYDZMLfEoHvQ/iJNOo86ldOQIuR9c7ptslut/ZCN6CAR
1cJLWwrz3POIr62v9mv8WgQIVKKD09eOLcNqp6tErZK1b/VoV5E+k/zcOSwwtOGD
ZjmnW+kaiQGgBbvspQE85TJXlkSztDE9DbZFqC2MSL5NUzRhLea9sjlaAQxjkOKg
vbzJdyI/bix1RYoY3I8OZzO3EeqF7Z8lHGHQNwlFoWxzkrbPUvLDUyFpbFojvf38
/jv/JEOO+yPiduo5GDCC7DMJ6h1ZMSJhMW0xH9oWykz6xoUHUb8TR4zKInHPUrPl
74vwV0xAJKAEE09VOoO2SryONkYCOBiui55aTFGn66Z58s+4lISMaLUNcRzOR657
xqfhw2MtoxrVg6MD+HQB6eCvR+YxPBcrR9qUoUeFbmiSj65xsNVaOLv7Q5LEUEp7
mzblxPFRH9t1O0iGbkwk7olrVEdvXhJ778cWp78s/mdatJFPz9XF7FYJWI3HCxvh
8NIQAND1szqTXWevnrQWX2ubX0azggQQRXuT/vtkIRbG02LSxIwluvcAEH/W0T2R
EGjc8eRyz60egH/n+KuFOd4mP0ojYvYH8ST8f+VcGgc06A0c9dkWXXauekHFlMpN
4tGzAq6+D2XWDY8V6R7GrjnQaUXt5LvJ5gzPrc11wsPr+wWASagz/skYoF9cQH2Z
FHn7TMVgyfOw/FTbTemw+PepJ/H9PDQ53wf9vLrPDHT5yJ5AMO/NftsG+l/lEaVg
7PvC4h39Wmuue9iMJKMRsFK6DOPiiPPJLHJI1HFZ+bdb2Jr2HxXEnucb37PFJHAL
zN5Ut2ieJuEXWoY6gapO1OEhbzev2h7OvBnJGxVDhi5vWSWHAQdP6n2cokjsSZXc
DHyyQWIwvTxSRsNsqFDZuTPoc3AqimVlQKOAGr6DqyNWn71fO5i1Vo3AfqgPW4qW
py1lFmkuLiq+e/gdv4BVA6l50Ph8i/g2TqJ7mNwf/ujsePWCfR6C3zKlv2kGlkTS
H43/uSZNQwfvsXR/wnsm+aailgmpN60/iwChRr4Q0tbUYf21RAQ+3avx2OuZ/dpU
SwZ1N8q0IRX6i8B8RakGkDZksGHOEkPMLFrYs9/sKFanOcgqAHXtIv++u1EhONB/
2o2and6dH6fVfP0chj6UYx7GNxsNpsSgs8Ls7gnab7HvXgeKc7FPjPi+binOwhdM
3RgiJn5V957ykn+OMvWayNBf62wBcgR7n+ydbrptq3tqGrv9rS329UM0EEUzlsts
vIkO3KmF6BHjLbigetaC068HpdXg4DSND/VkAP2JQt+GBEB0HYQchJ+TU9XUNimB
gLTZcJWNQNyEX711P8RKr/6ezudlQF7kugBjQYw6IQC0dmUtnO+c6eDPKtHOvOwe
wqNCQw5i5W5EYSSBkEdWeIwRglMivdBawM5gd93ZlhULRBtZgGUPPRVBrt+CdC7K
YwNynmb7QV7+3dKxI3fqC+IlRy3s2t22WGg+goZeb+JFtu2vdJ11qi5EzG53qGde
p9pGcPTGwgndmoC9nMY6CE9+glYXq3a+RlSDoPL31VyckN+y3vJrwwtg4funvito
V9R4qVaSjHI05r6oltHuVEa0nioJYhHgneCTqisA3p6UGhphroTNmGcfUK4nJyvz
TSxUkoDtKJ5EPqHQF8/QS8madRTQx6Geuen8kuAD8KGEKL6IhGpFNZyx/U7HhO9q
pWR8KfqknO6DauW1ylgz3e9H9Dtj+Wn5qx/yx6LbV9OCAFtaoZml+qDAccORxBL3
tqLzcMx73p9QZazVhshPspkuVECC6wYaHOM0QddBs7dRHFXQbnn/+9cnYCm9vobz
IcMpHlftJtfe+Ygun2VfneYvweIDOysD1TgS1RQG1vC4c40kQqO4TUKd+EAJguoB
J+QhH6l2ZQYHE7QkAp7qo6ofgshaWZ08F8SqcJwylpuq5QlJ6MuZ5FqTrWcEX7/z
VwPMVZb0Xjqgvf46s2CLK8p1rTsttn5qnDWHb2vykIUAcxfQKqGosQpUPWLMX44U
nncs16l00JtIdRPb6ATsI/RNAnon12m+Qx+CwYz+4Km6reEP5Pusa3/S7BJaRj+M
3VXoSViFi+E/GMTy/8zihF4xbaJ3Awv3LW7uCVsmMt8S27b5oXDI2Qh67OPugoMC
OsCDmBhzT/+ygL7jOaIcr4oJF8XRAyXT9yHnUy6dpPqh14MxeVbiBtUqQJrf8W5Q
IGBIDKWqMCaW7qmTGZ9uk6cnZdGy7Le1yvV+uefBS49YscqZRupxfQvp5oVF9UET
4d5ajd6Y4LF3W8orpz9B1Dj+GgvjatQitupKemR9P3PuFbZFFeTEF0TnSl3mw0Me
UFT8es1Y6abpuEOBHOAL4mqZ7KZo/XIrc36D73VkC8bRO7OfLUoDKkIt7tjDz40a
A8MuL/kpR303DaAzlUR9FTAFcoBYuu5jxCe4Yqt25kO/CF+19Vc3pbby2dtl8fVG
2ZP/KWzZXh3gehwq+Z7RbkDVSJon/sQksnOeaV3rt8jrwODss4PK/xL8sK8AhmBQ
7gNNTgMt7lNqvmGn91TruGe2W7AEwY5GT412w7QhAtAmn8Wv3t1+mQdydeV+jQxE
yMqw3A3gdFjtZYntySjVOlN1MwDQ+IYI6IP/HKfPZhlCs7O9vqk+X2pqd6bM1LD5
qOX/FHu3Kc1PiEuUwhbQvgP0MfDPJQzZert2z69ORWws+oyZVNdcfFIdU1Ml1nPS
BN5BbQI5EnbtyKoy7EvZefyQj9gTSBm/uDeJybSerll16acyt3vYpsBkDGc6wgTP
/h2ru2HFiUvnJpW7mB8kDWX6KRirX4E3Dm8yojBa66rnHvHAWuLr1JjhKWAovfkt
rIFf3o4q2/VO+vf1tb4+kFCLtLcq1VR4PJsUKGFYIj5e7t08kRvAgO8oeKXv3LIG
qYVMxRIod9qh3RfYpSchtjGMXG1wT4SEwAxZmjcEWOdF3csG7M+wikXepeFH6aNO
8Z1OLM+PbPvu4r33/eSUMlt3Lrfp1zVerNjW3tkGDLgIHoa/+gdGoWZAtd5Sf0ec
v5gLyg1jfUbQf5/t3Z0QnKLpS9134LYo4EHFDSBAZr2NC+t2alt42tQztQQ8Evyz
u8mrmVdbebw3t1zUPU7LFN3YfNJaxZ+5AJwcNPBbgMQElRpfdQ64M2i7D8BUHt6z
kWf+QN/Kzjyh8koeuUrIelAFuAfgC99yNnvBDv3hFvT1/51or/Cmjunz8XCvp99d
pB6+KqmCGOLYkS2jUObpeISW5yHpTxUm3Q1of1weZM1LiCs5Bs5JKnsaoASFKj7i
ZI2ZDvHv+mTTNZNxovsZQU8c9khEdvtYBkl+SJleQXftmtO7cegMbhA494zNW0Ch
ra8eGBZzkPjaPd4q2I2JN9n3KnVRAioF3VJi3bjEmImAG5mr+/w8qAX8sBzGBM1s
I7PpP4fpa764j8r6+s2J+ntdwYWd511g9HOnn/CKw2WLviz8MoMC80r6oor5u1IO
BTyrmIOZtWXoFFfS2kvEZDufOXMfivPFWxr4fMPvSwlVUA/DzXNTqoe7IMrNF/ag
SiVLBMrkDooXBC9Ff/zzbytNTTBU5F4ryn/3OLBbOg8ds2SOvvGYyfeqluM2AjYh
mLP/eLPyj5TOfD+Uksoilubpw+i/KeUwulu85j6V1KtogZFFouJ57tTyqo1W9gLp
/k4adQmWLXscZPZry3ImbFqn+SMRrETAdOMLZqQ8uI56uDrmkxdONjmNe7OSEvYW
ZfI+nH7TPU+NplWXAjl2j6yOui8ddGjRc67qQcFNrZxKr+sBzaKzXUyyyP5Nz8DI
Ojye82XBfVnF05PS+a30z1JiEn7pqdvKREfl+Zg5rh6SOKJ/Mfoli2WZ8FCyJrhC
DutEmvvAPk/75G2mznGNRMhBOQRYXeA6c07NcnAc2wj5h8nYhRFrduQzFuAKmDDe
nAvqjiw9+8Uv6XaJ2vW3zp9L3lcbY5JCOo1xAnhCuuubktqDAl+H30W49TESvMZ1
K8wF1jKs65rifThgUTG+Ia/WM9jLuCD6FH9WzsLo4u37KbAG41M2yDtHfEpa/6mQ
Y2c+uMo1WgPPUVbXzfe69fmkNzOSo5I45zOXRWitSAWyxamZYYKyoRDTWdg2rxDv
C/rqueoK4qJXkSINZnarsnMrcf33HdaNWy2kPNrkyJpDPkjTYtr2wFprHhc6qg/u
dGc5uBw+r0LJHTw3awurxuIrAd170r2nIELCT4fXqa3STj3j4TJzaMUb1bFJpTyl
2gEt/TkSz+Xkc3UeguS74Azob/QyHcpzwXqP8eHVzVhmVqb9jXt+sABWmfdo2d+X
XGjfRSArM7wrCXgoYnUWBneyNLXIcDc93l1hk89h5btSNTFi1DtlSFsRqd2J29rz
sdebPOT9am/KJWdgTZq2MO3J1R203x4S5+3CP4V0Lh/JOXxDOaBfExBc8TCWdoeQ
fLRR3s1mDWXerOH7j1V4F4nMARjFODZKYMccsVFUracqBkYGS8qDQTDarIsJPI5P
LWdHprGi+KL4S/01w0T+3K0RkpcQkVSwQPsmkDczw4tisM0y2jqfiQWz4SWg8lrh
R4Z5LbB62v4J3UZLqrsX/ovKToybEyJBfBWGfcV5IrCdflcfNGCBu/y6wXw5b7NG
3S3VcFWZhtmJfhEHUNJ2Vj2xHGyxfsxHT8q0RzQ/R4ZfO84mjhPvN6ZGxtvdu8ZW
JksiB7c6Q1ymeCeLltoaLGPxrhpqEXOS79Bg4T84W3sax8H9z1C50lKK+QqZVoOu
zoOoB15vol6eDwlk1UJRDU2ah839Aud6cIBluPv61ZB+rpt+AlLeBat01BDmq4Ni
gXP4GEa4s+lpd02id5ExyL8r3oW8c75hi++cHaKeISy4K80fCuDclMvde74jr2Qz
1YF889mOfdql4JsrsMAU8gw0snKag8l1dHfNKJqcTXpHDmdSFCqyZ/bPzOJGxUyA
J8pGuw2D2waQDYxUSJ4vObrDjwSpaC7ZAZ57SHItabhgOlveuh1yuXfi63ftG8Nn
7bMHZwLHDnApxhsIbdAaPzIWSKl9C1doe1NOAL02NKlrPdQsi+JnUXSqDX+QExU/
QIAT2op0S1L0xDI2Qw3vWtZCkM5pOE9ZUS7X8i/yp8TVPzmEUFZ7abm/ofF5TWzI
QLJaOxVOyLLisxMP/f5+S+9Or7ybCvtD1Hocgf102nD7rU8E+/tMRoE4/edlPOcR
nnvtVNNYHi3+in+NOs9j6XFGFGCFqhFtqOFU8RonqW9Us8Mjs0JSKaxVi1jfeOGW
EfSMt3hIVR+1ftLKc3PVXBzeboEjksg4GQdushQ2S0hDQiJW3I8QLHGWmDzyfED6
bjNSKx8vuugfpVUbB9RsXS7Uv7thaP0T7P56xumdr9rysMCTP+ggEgvbdcNq7duC
bnlsOK3ggMTcbkvobdYMBPEhgqorVdONz/M+PqIfMyt9wuwZ64jNQLTiVgQCUUhS
7wqBbXo5COLlL9XpczvDWMp3CZXLTemyer5ukr3JQdUtbcO4qf55hRdXXM2Av0RG
K6/jBpawBDFNzlFcw3it4hwEgyvPfonmd3a6GX9xeWmx+SYh4kf7/nxghZImcRXl
VNyXUOI97mukasJA56cieYPL2gbrZUusqrQuHRo5PGtsaqG1i8Gm8O9/a5er0zZ0
fdLyryrM1Jhxaxs7LIxSsLEoFt9busMGJFfGj8Y0NVy8f1yQRxgdIf0mypMAmznr
SLrDqA0bD9OMOgMMEl5WVcrpd6dt+TIr4UEVIxx0UfARzkw8j8fhzYn8p9IqH2jT
12lvA2XoydtmtJmB8kp9RXL04L41g+/glOeHKyCRmK5tA6nvMyzMf5zx1Q1fJCmr
wVu/ePrYwUOQdBm4qMTUZmgU+H0KT2QaSDutgCygRr1qv8p5x8afvKwmjlwrIFMJ
rk836j6u3Pcago9XZufWknjPnA60Dtrlcr3Nxd+lv3tXOjNlWtJEDaAroCQIA8OJ
mmGSY6GiZqYo8WcygwpIQKT1S44J//1lZS5lnnB+f4jL6WCWHBiDCHJcW1GXNAwJ
Y+QbagzoBe/F1PCgNF0m/HjIBxf+KWHBMoGz3sO9M1c136KRvZyQmvHGjAeWSkPS
lOW1ZekzE96VPfzcAhILV/f1QnbCsYrsrJ4pebxW1IWNo2hl6M89sL+NS1H2KmKz
BEvRsZoQgMOIzRjw2ZXOwgwuI3pdrkdqvXTTKLKkE4EqPAOEsmmPT4tKXnkMCxNS
LchismhEvSEXyhCKrwAWooYY6NpbD+Y0Edd9slGPtOvKI0QG8jP2c6JJsZMB1eqU
TSIrCf/pA1hlk+oROKcwmwzFm806+mOnWK4kHecmHU1chGPxW4KjUM929GjI1cyH
jeAAUGbwhpeQyEYK0wwiUVJPD/GXvnwTDAVYjAfl1Dx6ECGKEF8xddvADQddMvJn
LK765Xhdh6idhWI+vJYYKXBx/WKUWgWOZ24wDAJdaGTkgoZjdytNrohhrRXSERea
/ql4lBHNY+eVdQs+M1J1YVsOScENJW9DwXbm2JNSgfVTYn3lG09BsLuNrWTReY01
eoVB1uQaf0NQOqyHlUt1WnHeTnXtGA8S+0375zePS0pzxZUQjywbi2jh40NcUD4X
b3hIl1LdVcZlXvcXSEIDIVRcaYE3MTG4xtTYYiPdIZ+K6O4Np1XbXPeGFDW9Ghxh
dXRh9ZqrZlQrDYRE+SYfqv2TfFcjCUsDIDVTUqJNyrFL6Qfp4f3lR85/bWoWXKy6
jRRJP51A3xfXjUndp8Nh54pxU5VRKd4s59Cm5LtKFYidTufVREzlpoQPCs2UIaRt
nYiYW7JVQK3OrjudZObXy/U1fP6sLfjFYlfNN9fLojflpTIPeHBeBLwfT68UPbJP
/QzPP7PlkkNSjNVx0QgEet8+XJ/eZNAx8op/v75HNitmu0ayJylHX7VlbMdp9Jgf
PITBFSRakSq9Tkr9uk5/MAICm/MCCMWbU3IlMe5BcbbiPhNf5n/pJrbodRlcLwQN
GPQz2odmig16n4/j4Cil/SrOaZezWWPe6XQWYWMW4+OhfH3r/qeXCuwWUgYFZQy0
EYILuNgkXuws3KlgJudj+jl/XxN7DJ81Nbf9dqHP3HwlFGHUDbNVPd4LVJSSdOFl
GmEaawQUbn5fZJd3nBp7ErIOulzqI1Q6YZfSyaBQAUUhn3rYCZ08mGd9KaE00q1r
CZnTooyF1RWZMSvETq4rPm97XGZ00l8d/bC1vw/rzO4RH4iljJc7mxBbtheRbdMV
3PlPuUUSalpu9QXyj05HLsU6KHR0kAyafvsTNVL/iTIb7YxeYiCeuPhTwlI5KOwi
pbp8o99RtR1bgujSsd8uupOXoZcw7OI9j7B6r3S3md3TP1Z9GIvDrCUfXX6+DBYR
TTt4hYlTcbNtKA9vMR2GAla/Kpj4mPICgSkdSU1S3wlyaYTNu0u42KkDaNnzQUVZ
I69pL9dBrDZ1zJXmFe/BID6OjQ8uvGZ6pW7U/MCIqD2n7iD28vNoryohDByrMpPE
AkUORSkTk2Sj2mE0e9mCGth2cFzl5hPvcYCbmpT6vtk3yORq/PEhWm3HzbkXsfdX
PyovQvtCmD1g/7GCv49deo1W86JntMztFePhb+vC24nWZMhERwnPWU2AsosCuKca
vmlBvVKu9mlKbjbAmu61OkIYu67MCgjNzlyzYmxUUkSvLy6wxriLcv0lCuXyuZFi
Zc3saoKTwjCNq6BpHYCbLejTsTIx2uEWO2kNHv2KKYpl5DH+/rZRD/0m9+fPiSkA
PR6wPzCYtf9MJeqZtV7rfw/r3X9nmnP0v4ri1qshI2Z8UA/Zl2KtiLDqhsL48d10
dYIZnvhQM/zIn8RS8TAVWV21GszzvXi2Eja83mr6u4svN6GOqqFJmnSDQ78Kscj0
/l6qN7l+0xJ624lChsJ2XEbRzrtnhod9m3iXJRGhTWSS92p4MDyWyGZRKB8dOX1Y
7oulgzazZx/VRgag8hyaEA+1KuxdCvxuZXsWB9lNvWHybCauc/NWm6rDEmtO3ZF0
WbJt8zUReE+rFrrWnNzzMwXn5QCQEhBbyxhvJi1C7QyarNZyeSY9GDw5DQu+VCd8
rXwSgJSN6HFjAQSL97jeoZO+kGvXVxRTV8poDMUvomjaLhhzU1GW/CLjndsOeZRq
7W2B5N7+dLJHH1dFYj5AEhYOWyy1DsMUE+1TiA4R92IsByTF9Feursf6VtvF3l9H
9XeRD+BBt1h537E/THOKvPNNAno2FwEGxTwjPUlMxoCTe44fBQBjAbgLVyNUW8Q+
U+hQE4NKc/kvE2PxttNiO2WW4X2Cp1pw16f/Upe2g8JfPQNYFM76/aY/4OcsxgAL
eWkWRGsLrTJ5Kcyc97HLem4FUqusktSTrpnM51Wgh0HXiHPrfRLYkuHPYuozOpNz
qQwyNL9H8u1oiYN0i7M8OmQkIY257cU4UNG/8A4djUujyVSH9fkQfdxGYOX8L/N3
BpxdkydA++sJaHh9XBeF7yGO30sc/n7WICUF6E6gUpFWJhGdTVWXLgAzjB9HNnuQ
RuEQRExzMR30XKu0hB9TEzujfwgr9wfZ3h/Gw5OMbYxvO6HOKw4+Rg2/T//kc4vq
a95+y36CxlFKZ/HxhTbP+al70o0r/avlgirx5mP0hXqXRMwaVDPsFUKwQPcTQHEx
6IBdOCyuLc5BzuM2FIwkOWuIq/shtRfsc7FK++WgCrbn8nZOAuWRKxFVMONKVInR
bqMIJJvqhfCGpAmb/hquV20bLplxup/kViOpuWg2O1lw1X5rHVyd2saavFlok8/j
ZBuiNrqesRFZ3835G/LQilVRXl+kNUN0I2NO9K/RKN0hop+lUZXSYWViPiZnl8Gg
bb/BQfAPdM7Yt3no4d0lSucxx/nOPHU/+4aQZEbs3AwxVxgSo33J78MP3/Ns5Pew
EJcDdsabBMfOT9iLE2q0/iWeu3EFrMeCqcEZkU9932prkYf9ct7jS2y0rjXaaELo
kqunj6q5aXlhht5ZscNmDK8y4LeJw0ruQLjnAOUtxw0OUfTwsMehZUf/+OgDWDUE
W9mxPzKBxyjyyYDz2HHrUANouGS4eEesXpqEkQIP2VIMqLoemx30ctO+jik3OqH/
j5QiA0TK1IV1K2CxGgvNcUFLCc1pZtnTW9eqpLGYye/d8RBR0YrJGL5pJtfatD5x
v91/IVsTQmLXHZaOJrmWo94huJwHPSFTZG6q7TBbYVGfYFDYvMWWyk2z5+s7rtKP
LCUfy+AJu7Pm0AC5B7SroXbAi7Pnnr63QR6lYHvSt3K+SgQwo/a39MyCK0JqudV4
hNneXSWTjJEAiN5WQaePprMCXew0NFy8v3rnuiRDkd6vPlM9dSHbuH0ef9wvOyYI
lN8fSeuw+eiXL37b4HN9XG5X3zQUA6Vegm+vE98qDJnY2jY4AbbBp8Zz+wYpra5C
bY12lIdrtsQnTObO6dB5RApAyWi1FIWRouYPCWRTn8VXb+YFxhgOHvCM++nDEdBJ
NMfUreiRrC5NfxxCax46o0Ms+PXmmw6eDte4vJUQJHL6pV+iABJRo23M7IilVK2u
zDggd1T7dD6E/ucvNkaWggiL3V3ci5YgYNlMLUrvc3F5pm30BlpbXu5Dw9UjrLZm
KJ1jEo17Xr1RDIbXO84gak/wN9c+oxTqAu/5I0Rd5PJdu9tbMUC0QVL1f+JEuDvF
Obp2DTEAr8NK9fVyRMcK8byJGi5MUR44J6N7VftN91u1ur1lOv8HYbJQ7qZwE2QW
reVZdhz5xjTR1cwuyTxrIRGQObl/9ZjCo1NWnjpepITXgp67t++Z+WEQV0vrL9IT
Lj0lTdr++52OzUOYKkQcavjnYkiK/VtHbSlalf3QoF74HeaQ62PNuGFwrbaeKba6
j4/2bx6b4+Y+UCF1h++h1fw5xmG4HMBhXJBjk/yqdVigKosTp65C28zDBJ3V/Xh1
R3eTCGGdLxAap2DpYiRAnH/sVMNXcTo5LYLUBiCY8oVEUa0P7bYOjW6iuEPWEVwM
nrQbtEi06Kj4siLDWbs3DdlpujboV/faS1eGA7JphlhcHDQETZVt+ONGRTLT5x+7
44+0mE8zeOKrpT/jAYiTB+ylwq0SlZWu9lPhQQt675bwd+nPj1V7xBKwetT38FFI
xq45h3PSIb8dA/aFplsHvKsxp2a69AwsZrRMnwnFXZZAt75m6uZ+c/4AbJGBwp/y
oQsQ1vcxALkSsGlTYkXyRv18Lgr3XsIshMAO0N0ILm4CbV8s5/RVpyWnvEhYOuua
lq6FRynOkyadFGGv/gVC9LB9jEOyn19R8M8LnkGUCHahpiOAyZgbV+C814xz6t9F
2a/JCxV+CLdKMp7AofPHgxRQd0vE+zoDT1A43GlfwylkxQXoteKZ9lV+pHWUb4Y0
nEMbt8Q8mvFBpGs2iukiBWLknvgxxt0PxDXqx+yJox0WpGW8/Ntw5gZzoTN9U/s6
hc/tXgWowmRLiuF0iXhBBh6a+t1VyhEccraYvRvOOLCPLfQg5SrChCrqPaOKEf+R
9w5lOSd63vp96A2CtPny1IXKt0NjzxZ9ilAp6Pamsu25+Eo0ANPmW9d57TzdbQHC
mN+lPUHJIXZhY9y9XMKNX1hAzS6HYygu9Jjt0beF3p0iA7itY5I90g2qBya/hmgw
X6X9cpPgCwconIxU7Cgq3oBcT3EzZk+NVmMuicOJ+R7H+Gs128JO2PF/3ZkZHEfq
13nJ3rhH/XxLCB4yXMioAOx5sepNdGpKohi3N0jhlINloZcYKyI7R7o/3irz4kQQ
xf2NhifI+6Ju0r7uAXUnwCGO7ZMXhvPysCWH2Rbo24awq+3rvMyHbFzDLa1RvQse
707Qx54kOii1wyf1Eb5t3Lt1QCW5ZRzK1bPLqixucStbG+HvyjjLnt1S77zUBtNI
A5y9qsB+w1an4OQygCwO1NqKa3s6DABVv9nCwA7Kpu3DmKcb8vYpZ6djhywEG/IG
EAy6Qsbn96KxAviHcjjTHsOUgr9IbOJ1in3gp58YPG6WgHSjH6Jtq0KB/66neotA
tNlU0oVzMdP4GVywzb/l1Ru6d4IcBjsbsTwv4rzfSCCwFTGFRs8WT0/na+DhSpHE
Sh72VAyUQFrEAr801Tf8ooQpgNuGK654F3B16hg6nvbFJnKbQm3jLZsfaY9qe8jA
SXpVRD4rF06sqXOAkYSIZi4cI51wrB8OXi5uMNpyqzVhryX02DNmRZU9mtujE0ix
ttqb3eBYzXdo7/2aTrxd70F87EWD0iljUVp/voWnAXTQ1ZZtuZhop/HVf0RbGXip
ydOxe3q3Of9K9ngYDgPcOteIRnJaNI7mC2zb+GWUuqsMmNmWs228dWf0ZEvJwC3S
3XlIGy3xcfa4vpLN6Xgky1jrpndUepw38T25BDab3pGYrud0K2ZEBoAK+gQZwvke
Egq6/RZ6uNdhYQb4iyXFW6cfDs+l02IA+v0nFHg2PrSJOr+byl/+S5lcbEGX+8oa
7oh52BHhnNH0oQQwBsCdJMtGKepr4AyL9oee+knWlncfL2GU0WYMBXFTEYNodQs1
NWuyP5zSBqcuz6zCT++QuGR+3eq82kWICYv+Sq2JLbcIczdIUKqUrUTjd65sOsxz
3PK5YuVixlyRi2afAzNLIlbKqdbin6sAMnSTUtRwA60XSw0XVBOF9TjVwU8amTg7
mZvl4DDt1rPr+FiHIpk4A2/EncohAUuGV22cFOHC9uWPdLmNewRtqlhgQi0A+djx
bG51gh5e700exyf5KTzKY79P0F831cQ7thCTDEjySeXAdNin20Zt1nQu7wcpS3w3
uWTxBbS3sGyvVUabQVZn4RpdSSniKZ9d8kqK1J8fAjmbf56a5f0H2MKDhTeveB0N
7BWrPEkurO0TZSR2VzV9RRr2fJCIaj+t8jdJxxKx01jcZmDj6tCTYQWxCPESMip6
KmLToL6wBFoxYAUiQKaHjZCOO3iwCu1F9dO/1zqdEnUWB13MTUdxpTJY18WVuFSv
S364npfiz0FSZSTIh1AWzymeosnl2maSQARft947AmI=
`protect END_PROTECTED
