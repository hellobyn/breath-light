`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RHMSnaEmxQTQQWaq9Ar9+3IsucIjz2eo16FuTrH8wvEq4Oe13W/B06ONjtomkT6
kbPGtahxAk4KvC0KygBk39JfL8ysk6dZQIaPSMC8eQvkiEt27o2ZQoEbawpqhIEd
74a/F3od779yoP2xmm1ut2R3glkR0m1/qVXxQDXouG9BzzGodAttSI+iVnavPBAS
mEqlHxhGP2UXxx5P9yzLLx2QTXZlzgeLlIT88H9U7fQqh8fI3eeRhMWipMcTVJJm
0ERtrLACe7eeNTVeQeLDEzLvmCAY0hmqk9+9/BOsP9gVgXi+3OUNlFlZP4fWs+uA
koqNdJBHk5/CbNpA/r7z5jlWruxhQeFiBW95gBJSP2EqOaJaegt4kymjS4zu0KCS
zfAElmRpiUMZ9pSAnOM3yTnbphwxPav7t3bM+PxFzuSlxEnbRRnMQU82tIvre+dQ
Symoe385n4P9tOQTS+i7UMviBY0fy3QJVyt2I2o3xivcgQFIcA6GkKGNfX0VCb1d
P/y3tpiLaVxtxLFHPW0VwyY1irNTaJqTBWtTImtkI/P/GZCpsYDro8gbBxZF0M17
ndMXDveElxVbutyzCimv57Zqhu7wcMeqy+wizcpO6788mYHiFOReCQwxJk9MQk3G
SjcW4Ehtjm05ZY4e6GBaKUKUQm8EvAYq4TIf1/nvaN3yQlY8GyoqnoTQhiHGroeE
y9OKUyp2aW6OnZyKvbMdyFgTxw0n19bRW2qrCSUEXRju/+GHGddEk2FgZgDp5i2+
lnbS4DPq3wU1c+T4CZP7Y8RiHF0TRe44TYodaP0oo4+S1hqHweRvF00uQIPaoKdj
qneMPRI8bpdIL5XoAZQoZkM76jr/wVZrKKq9Da+ZgCCt+diHt6qfez/4U+C24hKw
r8/CuLs4ClWXFbQeqhQccu1WbguU5rP1iJZ9pOrkFIg2Urq2rCAaA40b11/X5qvc
NVc4XbRsf/AuaHpv+Q+OZvVyaCoIIGm9zuSeJQJ5h6C0VM6rOVfAF8UKqmNzEBFk
RQQaAUDN9nmY7/ogD8I6wjaY1KujUAvSd8hEaD07X7XvpreTdD0ldjxAcaGpcFBJ
N2ww76EICk2ZUVcS7ZABLsVXx1PAYUhHYBkPS6iBwNxaHwrMGMQra6I24W3bKTPY
soxThen3tSaISLZubwiCmhzVM/RvX6fz7Qy9t+XGiCpKIOlzyULzo5y9U2bZsWYY
Og38vMhmtliVFtuwNEC+Al+tZA9gvd257HYD15WoQ6vO6ThdFIiHAMzzz4tlpbET
UNjcQ9titBSFPY6CaxDIPJN4ppRoViWr3iEC3G0e6DHS71DpuUbgeklaoGEhbVQk
k8sgqn8dbUCs8ASTX9lcE8OS+x+wwZ5UYo37I7/ARUJMzQR9KcHX85mewMKjN1D6
YtpdJjpRZAGfH1K1gCwBR1ovTM7Q/kIG0HBPJxNZJTTpqpImRX2GafpBeR0PfQmg
GufzOTFnjDJZSzu2eM/+iklkyBiJhooTtELo/bRQsvriuZrThJ9/WBGA6nCqi3Mn
xLyD8kfGs1rBnWVjB9lIFLCFxADvKlXsC03/3M6dwqly0m2yIBTu57asxxyq6aNC
GK55uTEQp6/Jt7qkJsmeoQ4pHp1ch/w27iKHyBc6SPX692Mmz6q7JVS0HYC4fAsr
krD23K1oUfAIE6LjiALvc9pMGwl3WNUdXo1JKD2qju3QYUPBsvzmT+B0OPAR3SYF
NFwoWNawhrh4tQphr4qUAwJcUkFmvQX191biu6LTPPm10E16SRaI6eRgr4mcjCST
n7e+yn+JfI0rzL6mV7AuCH/wydxzixkEwRmtu/6g32pDvuQK1XeI4bfSWwGO9HOn
A3SgX+guZ/LsQPcqAwAFqosJ4c0gCGSgTOQWF29OduzHhT3gSQgXeBq+drLAOBhK
jTBVmEm6xJKyI0KF8ynXDy/dmh7ob6ScxTeVDnc5Ab1uKR4sktFlX+Cqv52tgZn6
ER/UldL8yvlzXqlB7R/9F1PT/g9YgBiKkN/dZsdJ3f3DJ1nPPIv2NFfCf2MfFss6
`protect END_PROTECTED
