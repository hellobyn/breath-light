`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Djn8K9CPh2ByBm5jWwG65FI7wfdpjECLIPYjw5WhXjPldBOphYa0EvtKKOm7ES6+
1eelNa4Awotq1G/laISs3DyYI/grGXHA4GnqbVELyO+xErS8L0/z8M87IRakJ6gn
VhWMZC1LtOG3AD3Dw3ybKwROT/miPb91zI3eoQjg9oegkPEV4LMak9LTOkOZt1zo
R5TmXYj8j4wP4Q433BwB3aRVFonT3c+mr5svPrUiRgln/fjtYTPrYIrefdUKSTmT
NbRyvGVq/ptzDcZCXgMl4RngACZDLYOWMFUPWhaogtSDCZhgKBKbcB+0bonSthlI
NAjMCtwn1etthV2Wx3pDDmqtdt9SzPe4++fMzZOclr+iGlVns9f+mAebS+fLhSih
eUsx33whfC97fbaCzRCU7tmmrslmB34EBhyAVZ7kTU8/FqC8mR+iG1swu+uYY0+n
hm7NM3nNgISw+qY5mSPqj7NeQe9uq4KeIIRn2tDyQEOgPi5nIpncVYYSaT2nXv25
`protect END_PROTECTED
