`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qnDTAG4fBwbjAMbCOrDqqjfWuoFcU1WuLkLgFr1ZQtDxG8g7A+lbTX9jwrL5nVd
957KGGHrFlAxScxNE/ykar+DVx8mNISbB8n29xp0CyTUM5eV2u+sl5pdpLLOwSz+
f0fP+JSIqGeuOtVHhH+DfU4+eAS4kqr00fJ0V97WOvzFuvZyPWKNlrwC5yoPDxNO
U7QMHuaMSWy2Lc0ozPCfieGb4CKXJrFY8bAIC3x8Jm0/yIk4mNYsW8pGaZx0FkKv
cihn7nSv2DcufVrn40MTIZCvo6E5RF4Kn3x4Vz3I3C1wtEqkVRzljMvetTnE+mz4
wgdHwnDayd4vfkGvqaaESDHEGUt3jYTKkasNDbdCvRS4SUFXLhiKut6C6BFFDTvr
OmpAPEYbux10BZck/Ye83Z/4ubAmAv7uQzH8qTdqdCVAfszYralKKyE0EL/k+hkm
FM1a1i0pmT3VfZAWWlJ/AcHYrHtjM+oDJnqzsm5jCv1xVlwHUPECeOkrbG4EwPld
UnNNR/iJ/+oCTHmA3uKrDI3qTcptQXT7aQZemNviPL3liEniGBE6raFORoILpY91
BLwJAwjA2OESf/JnlJNH95GOmq697gbBZIrMhyjeKUdOJf/BijOJB4/A62x84UCM
ecDAGlNWG57CAH1Ed/e9C/WTN7bSBsXMuWdeBattV34qr7QQNS3XB+Q3OXwlrsAv
9STKLFvlYFBGT6kdvOjTJYmXOowHIvpdVcSXTZxBEAfgNJzNSD00Rvpu22G4CSSF
RKM/F/Sm795A2IbtHVBzSdmMdZ/VimWClmpcjMOZRWSMgjiv+GJi3BcC8n25Q1zz
U4BQPmkX9KS9QsRGGIn25C6LhSFmwU4/HndVZdOZQfZ4PapFC8sdKHI0gmpUI4Wu
mc6M0CkJz10kX9jLNBVlAL861kSDFRN4xAjWSVPWTEJPpFfZNZgpAfvelwDtVl2F
CJanXaYXtPA2EcrYaY77Hfwo6ppe1dbmI2+Ouyro55AX6huDS/OyXLKoiRkoJr24
MJ+c8CjSEgXxZCWkA41NBB3zUl0LT7HCdn6Xz+j5yD19R57ujEDyLaTObnLr4YyM
KvO6/6EkbgBJqzJdddZCnHhUsrmJczPVNE9I7hqPPo4knIq9XnggjpIwrgOCIWhM
BvWMRMzxQgAvqqrrmeJa4yai5qKkbx3r3suJvf2eSUlhJFpFtN4PIFdePB9ztpzt
sZ/o6ZDE7L0xrUVbDzM1RNfXZSdvuMim/7v7nZWFfpBDYi8mGaQEbWwEIG/M/3oo
VO6wnAAun7/ZcmyVL5DgeO3jImtNVUHy5Zu4xVmSoBs3QEpGmxDDhfOcDOBTNC6r
DgaayrOXf+49MizxrFpGQCj7X8rpq1R3iRim/m0oguHLTxfBHGdBbrtsFOPmCme9
nJ8QC20xnSqm1k/M8Kiq0ZJ9qk8yj3yNWAspVQdBTwFtojief0TUG4lQWS6SAVZW
auNB3xGHIJ+aQQkUZOlr6g9rCPvMjiWmVYtNeFkhDGOQvNsPHlU83G3/arGGPgcE
ZpJofMS57Qy7JnJd0ZTrwYmRhHat3tf1Ypdhwh0DE0BCpe0M/951IW+9G530Gss3
hBieaP0aklXKvD4y2NUj/t0pie7l4VxMSqa0lYDSCiceyFY8RXodmOlQHG8I7egW
4zeb4Nji7Rbs1cqdm91CZw40OODYQWMULF48UlAQcc73LXn5qUj2X6OBP6woTjNv
m0aeqqdbwoL57tyPEALrcOvITEtdKPLvGb52PSWw/2YZOFNqAq5iWAf6+bCwOY+q
5XZLnyrwpQApeFK+j4ozAZfbo3Rwaj+a121wxRY3maiuFyqBkzeCxHCOEra3Ga3L
cjq4pN+1i78pUePpaRqNJ2wXcLHJe+y/OBr+OVo0RRk2+n+WDf4x7rJ/6bzIx2M8
Cs3PsRn+tGaJR6L+0LAp0Z57Au/NWpKlrJGD0qwQtoivEmFYJEeJPqEq6JUfWEUU
1K4U0ec2KeUYIoyNMrAN8rzMULXQzzg4+nlWk9/exHEYhjPyDIbwbw8RF/ocYYA/
S+EHH8IohBxk6hMJSy+Z20oWV3FmD+YmYJZYkd7qXFPx6lCDYAwogC26B7nnySJo
MZQCCOMJuCAU3zOHkHiVDqfuxY8Irjhhdn+d1FQnaRDRlOO+XNjB+sKMNfO516bv
//9Y5PoML/7PBPmatmu2tZ9vVt4yd6xjaXDVerHKLYS4ad8KonTxgrFKGz2tthEl
+bOShR5StHot86f4y5l2LGFuySWlEtawlTVC125d4cve8apRSW8qvQ/5JCA1Ey8f
nCxnoiG+jnq+tIt0NUyZ84dpqEcnOFSrnzIgkZamzh+BErNx72OiJWJS2CyGs1+o
zTIAQSlxUXapnIUl/MIK8M6aOKnSwvuzP5yhrc3Z9XXVNq8N4vYVDEE1hztvpMk6
VLK/rhZA0NqoUPBAVAudNmv2I5MXrA4c6Bwk1WUU3m19RlZewU9A9hF6XOY5rVAW
pZdgeY39bML0SelIb3CE5Reg8FZfD4G0xJbmxx+nfPJ3Sf8O/B2f8PBh0BOTvjdl
qLw2ZE0afOYm1g0MKSHrjOzn5VXq9qV8GIk7mlxbuEqQNqAXQHBtMLC526csTE1P
Ocd/NUTyCqfoiCvKBy4doXrJ/qKReIiKPvo5/BbQpqGZxE9kEsaLF0GZqxOnVLCZ
+7YIRJUK7WgiDeDb+8HiYWTxrzcTUURW6HsbM/8AP9eeAE8kgWZEoigqpJfuAlbt
RHBtAQILnkg8nhIHbKPvyM/o/es6EERIOnQgfnemQ9PXAcC69yBqJLnrO7SfJkEI
idjB9sZhe3BJzcav4y8DdsxD/7SC8N/ZtORr2jXjWcSwvQ2XI4ZgOnCftP3z9F8i
+6C2bIeHnUTSBl+ycL44E5o/w258ftyHY69CmNhgZjm/gsLEeaS0pkp7kp2+YuAa
GtfVnraFvU6KDqKkqlmuxlfJE4mXxoYs5fRI5uwG8tSuo6SBWg2HnN4x1POcNr6r
llsgd2FcQwu1N5ub3ImCnBKeRfNLtl27fHJXjwJ5YP2sw7MsT3zxZ5PETrfPjDYH
g0JLEQxYKeeLdvt4atsZ0WYY6/4K/+od7lt5X36Al7b29dmzNtvRYhjUEio1Q4wE
V8Fy7sGFYpscOl4IOvNsKWVqqHROTlORpbQKTCQcrKm58SCG5fbcar0KJ+BInedv
X/uDHB2exLAd59HMenmML6hJyLC2qVQ1g93rSfj5QIDpo9XBGPQRgUDVJPBJgWGh
0MfB0hPVPGLpiq74gtZhH5g4/LxoYICw2egBiB5hCTEHWSVG/dm8uaaHg+HnHFLZ
8RxwlHBq9DoxOtAbA2WBY6XUowY95N4hLbeK2ctuiha+3tQ9lYhl2oWDLB1AjBzs
Tr8DEajSIcnLEN5bPXtBUir6VrvzA8ryrYt+mfcmTzKAghMTU9P8ekYzh2N6VHNo
Y8TfDZ/40UvmYsxXiuFIs73XceLmN6yS+KIFC+7DTegpmz7SJ3ovlqKmofjLbv88
ZbxAxXujPQZ354LKw93eyR7JXlDK0bFcY3WlSDWE38b0wrddZmE8JLLu3jWNM1uZ
fnPwrLbuUjqXcnPJ63sc9Z4SdLAQB1IZxBihYSnoWYmhbaoFkbaWHZ10Udm5xWix
p1eMPiIZv185tH/3RT47hENeZvtGaDSddpqvsaJagq29lPwSCqXyiHy/u1uLgapm
ekGX4v7xMTgOgJzstl6OIIX7vsqP2cw50GXKXI3TjfA9O9CV0FWoSw/IxTdI5I1o
oq0smRbic76ozwh1B/2k+p5DJWxFl64iTBFJRudtQtmu2o8niACpBWecXSDta5v4
SAX4NM6AbFd337t7+xlcGu1sFDfOvcPCQiryrPsQRCAl4UuQDQgSLkHJYf277j1E
3NsAAT1bajze+XHSW0co9+tn2X6iKWdsC42TlMgp2fQZLm5qC0Zw6733hpWMVt/5
P1ixsz+PyGF0azj15Ekgwa92OiuEmpPjEDw4kft+Qs+0U+rPpmA/lc03StRgfVcp
GYxQ02B7CpwVsAmqbhdhsdovkQoeE98wdaX9XNxtjBVXJHg0VBFqv0VwIgldHLu5
NyJtx+6/YMcQKKVMT9j3kur4c3nvL6a5VHDXx4CFV78x3C6dxvcZVyLM1q1GUwEQ
X0rpX/9w2Kq3XTTn2PjfL42b4acpLrKBRcyT3kN0iC09I7rHec0ulyVkZsMsV3nW
YZfgaGGQ5uy17w1vb9aMsPVmZ2AsysP0eGSPikd9bahtwIuqKCgAqOgHm0ja7moe
9Hw1kHaXW5fVpvf1janciCFfsu8qQ1k2oouc1XPcavIs14rfvJ64OGyU7pp/u32P
qUNl46N/ZDWoXrmp+kimg4QBh7QbgvNxe/zsTbUX2vTYkyv7XyOc9aFC3ldyrXtw
Y6JBTPAhniAze4gg9LEdp/ZmwUFZYO4w0ERTBuFeSBoDayt/sOKiyMU2+51X60sB
/J6dP05rrBvAMtRrvQ6dZgdDBP61tg6Ll8GaGkj4tZigpYJJFquQv8U/8/J74vnB
HV40cBjkT7fJ2MpSNvfLjzP07qoFZUFr4Zkels2hmtmddmXKgWAnUyPatq8q9U+Y
wU1ZKCzjBJvgumGFdMC6kup4Cio2yCVVg0tKneLF8fCW+GPq/28VNF9ohokXxNhR
Tz2pbGuskxUzlTTb+/hZLaJa1ffggwRHNLErs9f2btdXAZpubjmoL+HTSTBli5uZ
MZuZS2toJbFFdWghmJUlK6nHwxe6fZtCGUqatZ2zjOt16GNn36fm4X1lToznIDCu
0qmqhhW2RMz/VUOex0KcHk7M57kg9/1Vv9PLqa0zNjS5q0q6g7zAVkJOgVTWPIup
MKSlI7mBU8Mc1Y49Rdv4lE8mWiUnzinnCs3WtqPcPEh2i1Tn5ZNPo/TpKZ+ag8K6
ybXzhaDFqK9iChBBsq80OR6z8g+1kKYOLxEq2/FwYB4AWo3zGcBytlH6pKvY48dw
R/5R6VoGkeCWZSWJEetDWe0X9LQmHqfl7HMAC/f/0efCg+R6Whzzz9CA5serXrr/
jnu6V0LhhH2eYqBUuBbkUVOgFC0QOtKuCNIguO1bepbS8WAdVgdsxnjrJfS8JQ5R
1jpKcCRvSpP2l1MmtYl88LukgLSkiUsT/hYcQZuosN+fppEmTJdDlCc4rvekZL5Q
Zvayx3FXlhoV6LhNoY2vg3OsaFgZ3zviOlYO6AisNsLCRI+k3oo2Im2m/rpSDUVp
tooVoYiTv2TtSAyr19nUzLMp4EU/shTdVDP37ccQXQA2x9skc/xkCEJ6ar8Etnxx
NCeemFo2uvBl2K/Z3UzgWX90vtXyOpogtesa+EuWJ7jl+4/6cVZFWOgKviHPMXdQ
vLVBgMFBqIhcn5v78JMZpJ3xdyWyTZIL8z7liFar+NGApySVas/t0g3lCN2zzprO
QzFHP4q714KO+0ejLXT1GoHBmM99REb+qzjJ0NM5BEnmfWnIUyIFFRQfbhIh3uCP
SO9mGSyvPEy3cAz1bxHN7wP6csulMrTL2ss3p6x2OXm9tsfwRI1NcQedmvgeAgZx
Jm+85jzQEU9yQkrvE4HTypCmnchBQ4jywrlqshGZLzA2hQQwAN1mbnKxJhX40Nko
7aP7ZjaOf9NtavATjYT28wwe0JizgumhrgyLBredQu8vUjN7AYmmHlFi+6ysqqsQ
FklH55GUw5PdYiD+k7XpKEJlhwzQ3nQIV/9IPOzpVWUr+q95QhuVkEFsMCBlEyMM
/5OuS91M21jvTP0Ifeu0dkCwv9Ko1U3bDZGxGEvKSOIlSzyWNsNeJ4FsL0sBBtaB
r16bkE0HekXukC0wnN2MCdXb4b2pJtYtjndMcQVIg6yAdFvtZc8wFSC2iorKbwVr
lDo6xtfmowrsc/Wp/f92RKQFuNB+tXmoKKM3qlWwNgR7wtJsIdmmSP6s5uVD/Mr8
k6VeCj/HrEhdJ3YxNZe+OnShVkA0BWYkHVukIG77WIQikLLT6FqV1MbP/6mxM1IG
fVnR65y8+FpMzb1fhpaJJFtFSpuqvRO3+4uA0Kh90l0gT5QCckZjNvbBe0NGKJKZ
KpibFom7ALFRopth67+CVia7l9JiyKRZtVLzqAM3b/XAtJ13q8du6H7Lm+0kq0Lx
Kn0f8menmQHWrPq+ek+9kqptM/POFZKzxufaMSMmll2QtXf4a3nZZABsEYlza76H
KeguyjyCYvhtdmZEoJyXdvkqLe/tm8G17wVe6z6V3G/2n1yqrlQnCieP636sKFc/
IQ5Z1VlsBAftWNU/QMedjOxR5Yiw12CgWfP6MdY2fJQN1bxUk3WuBCrbnMIn0o3b
dlsFKA8rUBJzQ2/yyeRdPmslh3WDO3kJtgvFGs7kv3pBh/47RnTIGdGuhFnVntBV
pUWGCy+MC+bAD7Pwj1UfnZh6c8Qz2F8ZoHX5Cd9ey/jsjYzajuoAD0xduoN53YOU
rmvwAlvDl4vDWPryB7bF6kVqJPYOvDzPUHlPMkWLi8JOStRcuR3aBQrl71yP5YUf
2LAeKAGVRxa2LlX4zmPG1a9g55B63nVvxZGOGZ6C10YF0QcFYzjEr/Se3pae+0j1
n/TLtLX3Ej7cHNHX9hn/c6us0qz5BzlCQxvvx0E37JsoZeT/2W20dZMarcidwMSb
oLi9HeAv/H/HC8XKZ++BeGyrlXEZ+QBip0qE7bNv6YZeWqA5/vGF+wwUqSOHyoM/
31yzGud+OtsXwxWZlEjAgnf0Oyy6092Aj7TxbAmK70ASyVtZYc3yQdI7TmmB3DAW
5kcI205u2vXUbStSUqQZLJ2lsNb3noYCL5/zFlqNRm2Cbrf8QtNqUwuVd/c4+/Pg
Evd/gWyvztc3a5bQKyfxwr2ABBheIgbxVlZwKuxDD9eFLuGxl/nnGXA/Jwrm6K+c
pGOn7QfnpK+0S69Bd9CHFxMFrACpQrRQAe1qbbkTGIsAwaSgb5t8mPssTGU/FWFH
DdwUVXsSgZApVKmTYUvB4mt2IlnpN43ZSpeeZFqqk89PQG2RTT4dbHNjMwNCehZs
zBxmG/6OrvHxe8tzaOCHKHbrWgauEC5Qib15tzFOyYALkMlDXg4X+Nd83Y42tx2e
sc5fwaEn8QkiN/oNnZdhuHjTwkpgnU2MA6wOfKuMelt/Kku5CgGOZg5xhh2+J3JU
VZ42Yq5DdBsnLPbprTQ8hlnFMyf4HUe/B6RpH9Mt+C2wXUF7SECEZsAoBQ/CZXqE
yZASeayXrH4SlTtPJ/AXfSwXnAPqpq2Iu8PQU2YuZGX96NPYWJEWjJ4KAo0oZaZ1
IxN8J5AmaRBVlP37D4S/LjQkZJIUgG0PoSULxg+95UX0vNJH8o4ZW2oD7pGSSHW4
wpGPAOh6HohEGh5Rruc2q6oQRhpBvqZLoHJJjfmJBJ6tEUHX1/+ipi6ZbFHTkRF6
nScOJHf49WO6ANz7rCon+1kFmNq04GCm9nD6eHzV4NS5BpyGYfvsGJ/bYWCBfDym
0O7K5SwsCvw7LIm7oDYT9G2WhKS+rEO6LyspgU7AiuEjYueGBIsJZQJTUm5BeZ1g
kJ6Bts0aDAxZeuAMOevmjr+rTHNA5uj53/X4yomuQTMzRw9dmqwuJty0Fuh0uR+u
XlVTyHEwMg5JOKrZ2KjAwlYrDTeQilt0NNgGWwXqILNixKRY6nxE8KJv/dZjTykR
omDzZcURXtMz+octjs0uazEhBCNK1vbFEKYj48FnVVFi2zC6NQQV1ncn8CFoe+wE
J8F/0vIzm+2+ngXHfWIK/42iSxea+VYt2Y/8V0cuNb8qMTXOVsK08NNhzeKL3L2R
k+FnPSH4Itjtk3gBgNwvsSLjTz541NxzoeWCJbcv7jrHMl5gDA8LU3W6SKB/Mg0W
tV6nquEAp7nQyAZI8V7edUep7IEY+hIxeiGdbwxuL6jp9bP8m6fNGgwuFTmDIuFn
zBAmaIgTYsBDTBrpZijY4dYdwqD1LTXyJx+tgx+20BkWoO5bj3xDxe45gNjbRxua
i2u+8LV7sAzLcmlFZq8sL3UNFYMOMNHCJ1DORuBPEzJgfOVXF6nTEBNi8DmYwtwq
IFEhtMJe4xnt4t8vzTIHkdyhFDOTHMrrsdB1MPXgmHS9YlbTr84QEMcTiElXRcgf
Mk/G11c87Jn+rh7yh5a3yTC2SzMNhAkOiHLZsKKXMYrxRvt9sd4tQbytKlKNwt3s
xnS+ijD6mitZ4JHEGE53HsScx7zD0h09w5mun8yxX78=
`protect END_PROTECTED
