`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgD7Q8oNlzNxxDikc63RqSiSODWeAy7pLTNa/i6gnJ7qM1od21c0FXP+U7nsBZ+m
sPM2cta0FsTjqQiUKgV+KZAjXnXBjH+AoytvXOch1UPuIoCjizW9WhBngJa0+qNO
/njwV2jQXqTR9wDo5vylwuAV2Hk3Zacxc8IpLNyYcDdEO2ungWqbwzHHyJWDrQMJ
fyaLpapNfh357TBYpkLWEkyJoAlmMJN1d+YgTS9MO5ZBA3Lr4k6jElw49aPaiT36
dbZtATZ+wCtxskSpY7heSPKfFv45aNyor/ILzfbpaaqq2PKT2n+55YJM2hvBg3jr
KVWBGokUdVlITGpV3Hzl6XTpPm5B7MAhiJpcankL5R5RIglXjQ/guyV7s3xZT4cT
efiVsxg97Ubk3lP2MZ6ijgIzThSWpYZPLMIxn6s31Gn9N7/ZcH/zZOYt1iUWkH51
7j8OgPsnFBBxVN1/0T1ZWqFEqQDaCINhLOH9hugvkTXjrqSJSvpd2p5EuCMZX4/k
PBVqClH73PMnqZXqoMTYB6R788loxQxX3l0kA6yPVVr4L0lwIdz96lfTpr/N+G2k
Oe7V3KUMnw/csL6XYx4k3l1oVl2q1C++eEuaySRE+6WAm4hZ0rvFrbTTxrOgq+jz
tFTpKMJRMWapFb/7+H+NWHDgwg8DNR5KFcSEC+/so5PvDlvhio5N1KaCXG8D/Ffm
HrpNNZTn/VAeVKae7T51u9U8PmJUB98ieFBi2Mb63oLVEvyiSWo2y1LO7Odte8V7
gqAdD/c24NM0vWCkkY/e8dHJYXV9sR6AcS3imSXMyqp6M+xVg/paMpxadoFGX44Z
U0PLj97A8/yWGm/cf27wwT1zzS1Z7KIwQKVnOPOVSdRWkgxAfrtbaXSDqiUMrkl9
pxkWnazfTa0GeB+k7XMCPjQx2MkVQDCUsat3wGlEyJYP3uzSCG5Ik/5f1S939x12
Cl5jQHiQriJfjiUGmtdHY/WyCRyfBmun0MlttEbQtwFOBybQR6czOj8i7mo+eaYp
/cbqCmiw4pn/8L9AAmcxnuOxwUS19hlYY/YmYrqiFTY=
`protect END_PROTECTED
