`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oceaghIQGPVvUJYTo/A0Ec4Wx55pDCwy+RPs+Rg0t+uZ4boEj1f1UynBB6jPivN7
y2VhHwsunYnZiuDefTPM7QC2w2u3301ptm8OExc7I2g/c//+s7SW9xD9dq1UR/DE
HBlvFkhSRRinPd+Hnr85QdWFJ5Q0yNC9tbf67gJFpVXtocnIKsVL1PLHsWBWpGKT
mmdum335tTuKMnieGm/is9ND9eGIWenqhlbtL9gIpQP42mk2x32EZtv+gSWhtuiO
H2ZpqNGbDyFQ3wkYV2TeLGG09I1fVGmVTPdinB96nHqmT5KfXt0nMk7tHowuND68
n9YmgxJ+TW7ILZ39hwxaAllERgU9rI0fwH6LJiUHXXHHpuzzd4HF9CaFmiJob1fx
+FHS839M2mgbEPbi2ej0pRyWDkSSI2spNE07+hTdp/v8daKx755DDuGEqqWDaQr9
g7aFJdTkKeWcHbfmLOpxJMn4v2LC1Ni2dsdEYC9kLh38MpbEhNpctYzQsXzu++Vx
ItMGCZJTZAev/OXQgaOyqUXQVPMccyYhwj6dhyNVsxv1V4LiDwfo76BBAAxfdUg+
`protect END_PROTECTED
