`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oD3JIFSJeYMiqtCsIaHEU98+FkTXb6xxFyw9bMnMhP4PSxs8sufxdlBsj+kGzb3A
rMBqIFis81abgHSsHzxK6ZjxEDqozuqoJGmOrZ0NZM8UrK+beBy9UQSW9w1UcRZh
Jl33nFS6bOPmUTYutP+gsfV0Pocsx7iZsobdAl8zWI5o/VySpxdnkMLDnGnIgtI1
a7uTLqurjsdyfFnVDdxz0LR/MezSp0W4ildgasDffgrZi89SY5SzyZHJxxDSUnt7
MaehokVxhtMrKbZslzdYzfcl48Q/+IbeFD0DAhFtlUuW4VRPtpoV7/Do7Q6hfbp6
tM1f6iPn+mnR1NPEY1yqDbOOz5ZQfhBmb06lKKJJzJZR/dYRpnKEKxEEGhv+hpaO
A6yXXXAgrCBh4fyw72BUymNPGegLgVhPUYeSZ7EMwJ8g23DzRa2ncnc+qsNaRs5A
gglb3tAnvK7Tj8vch9CsSWOPX+WG+k68hnwagX3abqFt1rhzdAuSIx3nP2laXQhn
ppA5zgXKJ3i3uDU4oe9MjG+qgQEtCDwYEWcYCDQcxHe9qkdjlFBJxDLKcizoaig3
Xhmuj7HW+d+b9yL+fSDk/QRhwCFeXU576ws/BlrSkcJ8C5pcnEHe0TpfyE4NjXKn
ARza8TTE0rBCGdAzNW2bT5jMfgLOwRd1vS9n2ZtoXa4Um/oLjoM44clJr8b71H1+
71lYpKA6zQ7JD9AhTBSa+I+OeXg4+tkMf8LDXO61WktWyvVMP2ofqVRoBkqV6SWj
doR/G/cIncLDnnqaiTxX7EAyRnTPcmih2GIybPVBV78y0aOMKeoUGlLzYvY+iGql
Ac0Pj9Yw0idvWw3joluDbwbAycvsCQZctKD3OkqQ9vr2n8B4dfgxGcNgoMGdkwMN
vWaZfAvdWOoICv/xavqz2jws7NZvPNzzkN7mJUCBexboqrNo4QSn0xleiPpII93h
C5w5pMaeFSZC34PZjt90reJVTbHiqt2hDF9eEZZJ9W+aa6SSJ3X1WGl0M5XVqprU
b5asbEHWiXqr52r8kDfN4z5++ksvEwDzh5JBXYmQbvVYzCpCHCjA6ySduKA+V8qj
zoRfL4wA+lT5mbjLxBeUZoIeUHEKsstPOgKS661OZkrm4ljMkBI3vF9MvtLJnGWx
h7qu5RBhyCxEmslE4l0NfvehYz9Ni8jjUiSNG3iMaqndCtWVoqgXw6vFcqPr0nRi
edPu7s3tj7kxBeVxEItTtWUyt/nMJqGxZfs45zHWJsR21TwNKWVmJuki8qLtPKO/
mazWIe5rAZYkM7SPdSQCtOYVX+8q8IiSKYRTLmciVFRFJw1bdNJviwXD8NXJmkv6
Cd+dMicoFreDqbOd62b6GnJpuMM90KdVDkOm9vhFWE/WCGPE35YC2r29FTUhhlOs
zbKlHa7eX+pL26CleWC/OH815oXl+eziTO9feiG1q4Q+JPKHgIoOK8F6BT82MQpK
I4O7qBp6gsbUhShROYh2EyPYuqODhXKZr3OBySsOk3X5XiG9EI5LzyMCQAFaIQ8f
L+ZYObBGdIkrvgwDsF8vr1EcVt3YNOo9LhFlhUKRtjrmmCZPaF7haTV7gPjDcFvg
nddXb2Vi8qwS8hMQL21UukzMCkTzaW/vf97HjO8CChjBRKa1uuhYPlaaWSJwXkVN
UZ+mC/STGIu0touifX6KC0RKDmAVjaVtAvBx+VK26sKKa9kT2eygpRm1H5unAtcN
tzgEoWSv9+JffV727SS013c8yrvogMproiJlRys410ngtUk/sl8obka0x+dED70v
CUNtfADFwD3fuYP5WnkT6Q/cDQddYcaCGiwx0zw+T85GHQUl3YGUFot6AKGqa6RJ
NTKO3rz2wXIN01bncFtf7UVs0FguDEhSwV9yZzhIp5Uzpxiu4bDdTI/7tT4t+lDt
XrX+i8EGu8B3ZD4GU14Ijvw5aFcVglSg1rpYeyQs4Kpzm/mcXYiap81oM6AQe05I
VmmOgyh4k6ZoMD05vmGTp3zOEhQSYva7OXqdt2q0xxDJNnXzBokRi/h972csSm6l
Hhw9lGIm6gNiWigW14oWGe8j/Gvbj9vO6l4bz65AMY5qLRnbDWCnCiEbMOr/fieg
O4wMTX/AI4xbNFQzKv2iKRUj2w1Oaa2F120eG5hHbpLKSvIwGiDKXnlry9tl5X6d
mExXiW4Y4pfOKhDr2gjn7nduW00VK/CKINbEJ2KxBUtx6ymhC5bHh8emTsudkY7i
yywNxwrMQyZQV22/AO19U5S1bq/wFcjHlnsPdIu/BhrGleOFgII46gneuE/N+G5x
MMA84bR2fCSR8IgZJJ2n1F+veygTxTuSU4ujMtPb+no9sbQtOixiAXoe9Az16fWC
1fssWXcCeQkgS9F18S/4uYsU67ALtzh/wdnmdOUySjRn4eIZlc8bYi5zsgdTvFjQ
+xAmPrV2kdQ097mAwcLBPrwmEa4bZOttNl675JIFRgWR53bolxvmLv72mq0BrvUz
QGxmmqmABz01QDvcwG8xxfGdg6j1D/53RYQHNCvlHKwiNRYMJ7LECX0JB7pLgpJT
7KW4XKVW2Aavd/F08ikf1AC7AMKdWagG3yePb3cFQXNTdQIf9pW4WJMSpku7fOz0
jRRDkQVgZlbwwQWbmcRWXBJGI3FLQLujL7L/pkIbZobIRutT9GvW6EYwDLHk0FMS
bkDtG+OJZgD/j+cko6E54L1yrmQWV7ucebyLX4CYRK37aBK4ANPzAGj/atS3EeMx
7LmPTRM5ndqoDEPSfg4/XD7TTK3R456i7hLiyK5lY75Azd3mYQ+8VIiFP3tgEp5Z
pfCoxGVaI1xAFpZHOB7ex+M2uL1JmJZS/KlW1ulO/NDdmfQgCxUDOzbrj9HlieUp
iqW5KxJlVBc0MremFsA+zOG/E2RAdEc8t/ItQCaqeb06N76cTlQGeVFvZgCgQjk3
hjUipyFNqOzBanxjgf2iR/tt5Us0d/FEznuy3Kif7ShBerSIrcVaWZNTN9+AI6T/
+MJdBaH14rox5p+a77AP0xLCRWxU7ze5y2U3RYTAGG2Wzz8USevGnyEAHiRr3uTe
VBmxG+o+z1VHzsU07t/5DuVpnr16S8nF3dhcUgmUI9WJEhpz9YpMvJNO86fyL5nj
tNIe1gM2u9qOVPIKWtEoSneRSd0O6WwTKx5rocZ6I9VvRrtckcwybi6iOI7lrLQ8
fTyfH5cw99wCr+Dwo0dDc5QlHh0RD1PDDeStUtT9f/EIru/REqjegXij1vCEJjgl
ly6MdIN+E6bTWNy6X34shOf5D+ohelLTDVJdfWFe66DyOmblJ6PG54NAu8Gsxbzg
zA+KLYNzvMY9rafzUX7JJ4AcC0qb6WBZd+4isgHYhyQcG3GxdqRrEz1v3VbGwfTX
7nfj17ZGF2ImfJrPZ9jnXwN+tO4TDeu2zpblooiqgsAwH2gOAZfOEXFMX+8Hs3tC
g+S1W/yYPWVSmRizbIQlkZ57T6YPMegjfd5erNGchyf6EBU8WnMMo5A7WOTCWVUq
q2UH6NhVtl/obsFP8Duv4I+d8DTVPfHfegw9CLxlwWgcryLe9uPysiHglhmhR+hg
Om6o32v9BTNfiIHtRu68o/ZXXT/+qfKLDd77ISaa60DEkgynHhG71HKSpSrw2p5r
yjr68qpqcheRKw9tT97C6f2uDTG0NKpRG8gphmgtKWw81fEA1qQm8iGelyir0lbt
CDkr3CQxUqzs2bvw9/26pFHS0RMse0KtUYAsh5pZ8AWRVmsboiVL0f7P1CdzifeP
vmGNa39/qlysFzS9OMJnYw==
`protect END_PROTECTED
