`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krW40rTcDC726BFBmV3mV/ZyBf+pwafF36QGpJi3Z6IXg+iW3IMRaeEJtf3en7AU
gQe2COYBwdYBeJGrIl2+IId0FXDn8wRNP0ec6+IyX4Yv6CmvTmEo71M8Hkf8HeDy
fhaxiy8sdZa8enQLB1Y3eaSJLZT65g9jZL4Ex6NxqkegL/aflEPvYa5kVxWajjU4
pcNPJs3DOSCZqecPremHYZfqGlWZLWgp/ozzK3YDI0Wh7kJuOWYwjgCPj99W2Ojo
7WZO9C/4MkDtAKksDMnHcoMJgr0tBbpJItNgYf2F1QFmwkkH1JJtJKdXozjoWu6p
NfQtQJSYP+10ZsnspptRUqnk1kG++0qGsxPOyXF5vdCCKh89bXevIrE/QpX6qQj/
FX8Pq5ZgSRlWLaPC0Q1v0dw1LbHNXyNc3jyANNG4LdISS3wlzVCku/z58Wkgyeoc
v7LGpYZj/5DZFsixwf8dcVv5JIck38zCcRZbmCXkm+uU3X+fomKNFqlRggXaVQ/p
wawMby5fzLfO8T55uapC3XEZlOquqiVAiaQ659hzLeqdguqa4jYiPs0gD+edzfdL
OAiGrdNzm5wsqydwPBAOXXiHwaEVpKjGHO1sqhUIXVhY7hh+j2txnMweKcH3X8XG
w/UL8AJlbQZzwq+A3hbaXmrRuikEOXzb1hOdwJLy+SeLI50pLr/qtYKjjNYCjQDA
7AC47Wn6b2A2TLq5J+8+V2AkcsBr5sWC7a0yADxECCvfAhLzpa75M3xFL0ohJhqV
7bpEPSwBrWGG/kB8HfN3f7YahzHxln1B5BqbNoBo+9l8sRToFwaM+AGSTO+tp3K1
uRNO4x/H+O11tZV+fGMxVnLOhm9x/k4Ba2AW4o0KdpY+cKkMQxOy+NU94/gZLmm9
KqJBBfuRFxYMaD+e7dduu36RJ+NThD3gWKBDSy5n19JfwBTHc3/yrUk58jtFLdWU
aHPyRb36pmOZU1Xo7DVzbN7s1Qkyiv4WIXCl7Fpx3d3tSazhj0GG7qiuDeCGxEec
374N830uOmeFi8zYBZdJi3Jx3MA2N47QC4mhCHxX0B209sPfD6SoZAjH842arwT0
mjCXO9yNogzUuLiva4YEcRbb3yp8xHmiaKD4hM2+zk8UcJqnRl11E1nyqmTldjU6
w6WMDxU+DKT5ZzZoUr7lWr3nLF4ovbs8aVzIZdg6RCRmyCXrG5iLIs561+yVS8ch
4K/Jb2aiYwShmmLMjqXtRJh5n4j5L4ATzIJKeLNtbC18EyVj3KmLOnjkZS4uiyGh
8fEr9W6WH8XIeYv05NdYvcJRFgrUiw5z8hMz3IYLu+vcdcE2R2kkCEDRqW7cTV1c
1M7+EGRl77FddVy6rAgOPwOIzbP4e4m+MzHpIXc7upk/cTJ+q9N1Ab2fPheKKca7
VKoEcotXXIO41TYV4+YbOypl6BWT6D/fxEAUDsOp7nUZvbFSnm1mNKt5RZn5jKkL
T4GnRKjH9huS1WgyKPXTJO7LkkI9hz251e/Xt7AJb6HIhYmvCV8PChIeA6a6qjDl
nWkD/+tZKqUSwisaMJ2IFSQtifKQJqLQqFBTHso/2ub6Xl4StkYTXkDVymKjPreL
bYvEtF48rCUBb/5PBlsFgOzZHXpjsQotONKsOmhy3BY0J9Mdr5E205L1FZZsGpI6
V/u5kQATec6TwxQLGeMKDGFCYh1pxPjgzfxGHAimkNUd9zLG3iB2/M0ge8tikJ+W
IFI0wqLunPuUmJ1SEaB6y17uqyP36qpQh9R6EwxLj3WIbDPlJyDTkwJGq3ofC1ru
OcnxZUVq3OmGFH6ZHgQS/7bPfQtNMxN/F11/uJZ5na2GK+h5yrFKmP921u6L3pRa
WQe94nJNJOCn1a+/YsAvytJ9Yp4bshP2lnVkdAeNiTbl/0jRp4SfaJSVEoTR+Hk0
C+tfj3IGnCgGuXvU2zzrw3htat4Ay1QmIWkmbcKIBl7dXQwIIMl69CLjbpqmKuKU
IIvrOsyUCPoHsoGZ3Y6Gp12RMYxOmnImlrBFm9ATW7Cm7KkoJXpytzLYMwY72XWr
ohnGNuUVYMZaVGwOPGgOKfpH+k//jITEDlmB8UmvImtStsxNSMAgfbEgobEC/TX4
QTxYSajBqboulJaAu85pLHW1UZm91fo7j7BRnrAAN7LwPZlDPagrfWOyVG4dtAGb
fvjtQ8aMDPD7zwNoxN+CIzaWa73ql+/u7QxTUcExDUfXP0IjEsEJZ+CBhrWLWo7q
Sc3yAO01SZnYNpfuyV/24ELyfI+2yMxTUbLiSX72WuXGKz3aCjOjrtC8q8wZAfxe
7pqOWBTu6A/vdWwshdh7PTma4XmTr+BFScBlJHHWURzZrZO3P6HoeUGLwvehMCbI
riILAKFrIQJAiNFwp67LONwbu4j6TthPl3TcTxD9Q8AtuIMXafVOi0/laIRrL1zE
mBQjPXLuiJkkGHX8JbBpA1Q2wn3W3+HCYb6N7JZRsVpGfqzFU8BCfPmNAfAkSxeZ
/hCu5HNLanq+yVgdFVPdCphLYCnRu+QiFsJbaVEHc1mrA02oiGqgmYmkWg3f8PBr
9QUjq1A0Z3kr3vYZvVMXq8ZqIyW5maJ/oNfGymktPGDxRsyOkjBxCNwImjBOES2i
tTlIu1t1WFyKDHB5Rg52BmuhyFb/s0tfft7OqavK5SOKWnucDeTn0sXfe5lIaS1q
T7m8qR8QtRUGNzixwB/wazS0cVK3eBcNgEa+bk5zn+rdJ0mixu8s6FRGDOxID4Rv
ePZ+0g7EednHnAryvHAUfARltZwVmujHBi+kBccBCvnsKTadJoKGuiTlJOtsRbVo
MyGWcBMnfaAfZf0ETf1r2ubZeS9I9RXbGK2dDpyoFbeZ6eDEIcLPZMRxr5jZu+GX
olzG3Z88wfCoMNPZk/16DWQEc5BBaaD6jEERxYxAAy0DLzqu04dAbEN1L1je531l
DwloWvwGj6Qb00s9BwseZtIzU3eVV92rl7Id2fX1m7cYWDOVUQhO8z0MAzi1wW9y
7b1Lp2Uu2rVGCBwirzdTJgcsbO3Q/ZzVjbifPdPfTIkMJvYTLt5OCXL/gH5YwCE+
6dlPoS4lZ4Eq1dpSKUVsZt4gkBCFnxyB5rRaWuTGHyhH8Kdvf7GqcaH9lMlaowlR
9QaHUL9FZ5YNxfngAx5yyKxA6Wlb9KkJSDq20vfGwB9Z9l/t13kxZi5E+E+T0LnX
wbsy/w0rlO8cXMmA9/a+V+ZK4yJ1aSbKpXYuo7/g/PSVY+cjUtzoXd1yXh15n1sT
vsf7EDUEw2pZi4iSB63HYGplIqwyl+BGM+FGR7Fe4/wgf72g1UbeRlmoFVO05oXj
aw4CXfH7Oj+w9nIVAZ2hSXcmNWgkwYGAHOD+B2BAPLz9RReTH9x2sSayxokXDtcf
B4j3UG+pSDuXxzyf5i914V7heP4lY0YSEhG3Dm5WhXQQkFqzxZradqKOBrQp96Cj
9YXpj4H9b+RB2s2nlpKQo3ZyuQyOfyiOvjKddb2whUeHZVZk3NJMOW7bm/NMjas7
cKGFp3S9s58vdtL9lTL0Ketb0XR2cbKJnxF+Lvcl3Gd5Vi91edG/jjyLvcY0bRaa
Udt7Is/6+5hpQ8jH5K2ibzmtZ2+lFUJaAt9a7WinSU5td30LZdQz2SJOgFJR94hz
xiqA0aQytuX1DfU25Z6V1THC5vDLh42R8ISfL8R3BKEppeds8UMRnS3jjttCWw18
7aYnMiRAb85vYBUib+79rY/KnA/yxqxoSV5M/E6kg0Qtr9zTL7+hIjYae6Qy0sNV
/YPhLUsNFTu/1esWczNoavAGdyrX5EB3DVuc1zkHnWta54qqynfdM+EsK79Cv4G6
6TW8ZDOJgEUEMw/noG8uS+fs5tpNUb+SnUSU/gT0KK91Bt8jvW507IZtByOoZqLq
KWqiVmTvMiGU9/0a7lHCHP1L/ehS2x9bq2PDcSxS0Y9bRU20TzPETdfy21TRu0BV
0Lg4rRS61xVLxrAdt5phbWNESw4xTR7BURqaUeAj5XW3xBFb/JvNoheXfJio06n5
+9Ptrhub+JRaopzhXEnjJYOWNXCRurCfXWa4cgx4/75dAnaP+QoZKGy8r68w5T6/
q08uYhDlR3RNmzOlGN7lxr3CesNuiI5mKKG17nTC9Md6wWa5IBmU//x5uDotoeKg
RMAk6CWnPditrFwcuaag2p0pwkJ4FjC5y36qTVaQxMXgaR5FbJost3Rv9muGxy4p
nHdRT/nhd2AwN16XnaWdnL6Mf3MW6UMzqQAeh8VkYnUN86wyn+HMNmWI0xfaLvpE
WW1J9wh8csSyqTB+z9rnkpiTnDDCHIfLhlaXS47B5iyOZUdS/bO5mACZtgEF8KSv
Vz85q7Di14oWIq/HIcN0ueyWIF5/h85lt2LMCs374IbBh2kQpTIH1IS38qYc/jLD
Zw+bUymAgOA8yBHRABlB79rZsihQEP2spydYkCRaHPtZxUJo65lHRmtnAgOJYs+q
HXr8lKPN+kMqL/vhdmHb3r6yR27ccbD4Q4jI662ntX2vmY0bdd1lcVUZWN6rZ/XP
tB54XDdRN7bS2+3UyHBeVIiPs4Yc97XLp0TOhmSGWDH2FcTXn40gsAX7cu+joyf8
qlUnYTIUUC+lLtAG3DN/kA2NCR5h/iQ5IDrrReYUKPMhRXSr/Q7OAGe6NQUj0QHb
/9yStlqlaU+qNOr321K2aYBRM/JjeFqkTG6EyDYo0VMdzEdCUou3OHALIwdSv3jy
w2KEsZjYdEpf0ayj60RgwE9G4WAPIbiEjDuznWllhOtsmGQrRPmmKKahfiLAaa2D
twB8CEcn+92QzYkR1yvJYRguVLXgb4G4SXnl35BP5LuL/MINf04ev/mNK3FaJ/bA
NHN1hfqK5JJa7aC8bhNd1qAjWxVc8oprnc8SwcqJ34m1VwHECmhLIKq661VzGhmr
CdKvaJLu9lzCPd/0YqXLIrXb+sN7GVn6sYf/EOFBMZNK6tcYiYXz96LhKe8+ssqC
DuysjKkSLqszSvum5PnDggojLU0ehB4eLbeRRypG2Na47fM4fGoWRRaAw8Uchq1b
DAP2dCOq3/W7qBw7HMup07bTfTPQ9XPYuoRTV+FH3KUphSnPPeq2k0WCnsUtxU8D
qeUKefGp3eoazCDZE71ArasO/bUiJf/z2cskjcqsxPdoVhcWbnH3NppRDRe5V2qb
/D2NqcBWjamChr1rAwWneRFwr/Q+1BaOF65eUkLqYuiwRs7jjXSfwHmFym7Sz60/
uRM84GJR6JoIMDODPOZFoL6L557zHJ2t2tIB+L3Pkw98JTX8Up2y8l4bf4Y3fwSN
YrCF3OiGF3EZ12ELIE07MC6yJ9XL5TAE6zaTqmFoeL3ijh4Iguv06910AGKINM52
2hp1J5YSu4T7CAvh9fPgCHT+dvrJpIUFSCrdnnV64mAt9TSbcywaBXG9eE7t73Dq
5Dy/Bd531qLzUb7Km2IyCxSBJ2X9jMctYCZ+bQETIYrD+UCSFrj55IJUlA4d3HJ+
00iqsjuxrVEw6FR14eKQMxwrVyttT3kX9YLwkDOnkP1aWSPvEIoBcXyLqAIk5Qdx
DIdOvr186dKNYN+xRtdfHb9o2sYqNZ1KOi5TKQZOcWZx2I0+YZ9hIyJkc+gH16kj
H74P9QI/9br1bKOXTxscUQ1K1xFkVhOB41Ty9XMAjUdc7nOCrN6mxc36Ggm0UF0f
R2pljaiNxmGkGB0PklWC0TDpKUewWYNKa6o5jJh4Ts1aZlG0rxAtV9eVY7UhZTM8
YenWrG++z+xRWz75569+Fu4xKNWdPJ77KeERvJva5qgRDaCnDY0hXXJS95NSXbat
1Apz8LMwzBCP6jViKaZQQrpQrywiYzGGWAGspSOIqOPb7ezYwcQ70CimC/Tedb0z
57GAVa2ND6NP1YcqdTDDFfH+QF1n5aPC7VpFop/tOoRe98EL7MHyCCaYPxNHEVma
IVwuVICPcWz5lSUPHDOU7yDSXS7xs5xALwm7RQNbySXh31OlZOnKndM53t01WtEO
VTKSL95X+Lp/S/V0Rv8hDGsU7uHTgoV+Ui1Ar9Lka5cAthEhoYrsJ54/GrHgX8jS
oeiRJiG8MvCcREggOBca3sUE0aorJHYC6NfeszgtipNSUHRIfarhAd2C2Ojn+yDZ
RU78/OFubsIxjomSX9BRRihUUZb52ZX349+zt12IL0CP0Yb6IeTkOG/A6abk8DBq
VClK1IpfORU9UHHAPrLQtL+xbJ67DI3cI2zrl/zIMNmXEIPzIZ1jGQUn43oRoj69
8ck/GpKhRyrpFXNGyY7H2QMqkXzEK8nSd1GNTEHPR2KbSteU312Six44cxWVWZrU
Rv+l36EzRT/1thIfmd5sd9RXpWZfZCglD29FWE3+e7P0ckDaxEhvWGyrbyvYg6/E
oX5eVAZINLm+IuA0CmF3GcovFrR5PJdVRC4xsI+vgS3N310kPM2szFWI3/RK7blF
7X+k8bxlKmycVWQhkfnoNjdAilqfNAy5F9NSoRkTPyotqHrweWK2NngZUUNYHJur
ocrO4/iZlBlg8Ee+upuC2gbD7vKOqpg9f2VIconnkcRWTZTlDAvV/pi2AKE+//ct
q7+fl+JdZfIGoYabrgPLpG4Xz5m5sgWA6bLKLr5ObsLEMJDsMZH5W03UuKb4Pzcr
Ye74Q/3GVqtIgCjYct+AyN9idwZQ0bev99tBXaIkveqC3cTM3XqzEy5gWHs6KFAt
TARObWWOLXq3x88d1QQqzxh75hYou6D4aKKBhQbBOuRKwGVj/relSbKJrh+8CTy9
77W7OcGmV6SApNQoUiNDGsxtH6Rmn8bAkDbmRiWDIvx77+6eEbZSaVImn6dig6Rs
naWekvKjnrtjPAVm7dqkVQp59x/uSrJ60c83haaD9TBGBG3LTlYLJoqmH+4MtBH4
sIA0pherHaGQ/ZJ3z07XItSJKlBK112tLaSJIpFQ7NACYthMNZ6Zwow64FTYsWSt
WC9N9AfQnDJvUAesOjJUIlpgQ0vAWCFbGH7+mfVxWTEZnljVhzBG64Z1OCWIPFvC
Pk4pOV1tHxIiXUKQyQoshLffJeNdV8/FDOGB4cfei3n336VZuVc4LGP5YS2uIRma
JmdR+97+xqd5G5UcTrRKePJLzUdapveBmYE8tnGYa1LcbyChM3AHFzHJfTcCo4Qx
EjTjgZ7gnpdpRf4HTPZypt586qy0OOr7aXcBghcPuBdWMpc9KMGt3g5ONt1Plsy0
AkbfFwihPW/oUo7JyU/q7dyG5HBdMxh1iixOtH7Dpff+lf88sGClaLFfYGY4lmLt
FPYqSvJHST/uEyHcRyZMqkXSCuP7oOMLQcEumQvs2lIoPjhd80aIo3LWYdrxooKp
bMCSuSxoXKx5bp1nnbU3lFqZJoR2abQSGjWTkXwu+87ketDU3cUUh0XTO8TTBamQ
zoSH7LzeEfIpzV4YNZGTIMFMk+ArXVWBumMiSolWW04HM3KPmFaciAArbUtDCBeo
KFA++hk5tvgXbxslWfFwp5HZeNDB29oajkj/V2EFrtjb6BtpM6LLCC6mD2Y/+xcL
R0DDxGaMO01mKMMGwRka3F0k1WXjLCAecN517Gjhxzk0R7Ib1tbkodDZ7IgTlMV/
YnvL6yhF9gO1zB4dGdIorWwtEs2oSwPatKkzPmGesH4gYp6nC4wk7K9Kfm6bXaBL
DaXoa5+fynE00G/K5OyGs3r7CNZfy9JezpnAFw8KSw9yMV1T06fdSTBnJL2UvjRl
dJW0VXSeOWHX8YCQ6hCtLCpSHjW4mtGORWdLmJXvp/g6e/4u9PtS25ImoM+Ui8CG
G8snoBNqa7GsjI0QL3t6KlpoiAleZJr2oxjnISbXm6/EdDJ5z2UHECc2tA9OeAM4
HcwAnRabvzCVbO+RoBKb2FFrU/9RESxAXQn2tULUqzbtAfS81gMHPBF/IcXAtTjL
7GfE6lAhC1yiBOu8o22GUrhmGAp63uIBafDCR2Rib1KdqTe/yRtpenF5CllR+Kg2
ufWKI2qTH9bQBH/52e/H/qdiQ8wUxtpTaGljN4yvVdBrJ/EeUfmotdcuqsEUZPoU
KghKQTSkji9627J7SVC9upXxso3o+LAR0gxRXVx7u5sW8ZSCvrkZcuUxQtcP7rX1
Lj8M7Ejxs5+NmL+TEdz0uHSrBfNw2hdKtFj6Zi+j+j6dxdv1m6aSEnjoulVGUcd4
M11f6ES8ld6BTPY15wnjsQUgNxdz5XO8syu/cT2daqT2igdpla4UmKcYKlZ2Ri/m
//XLXKi/dfJZOtzEk0a8vGfmKfdwCZnYPwcyXWug6KpTT2UyxWoggeR5408sIZYL
ogrAsgTCFpL3ypjq4jFTuYT7HNwQa2DdWf3v2JUsgfn6KRxZc+mxBJ2UKxaKQ5Hp
rhzFxmmvn/73cZSYQZ8sf23NxlHDbhZ4O/29IlaLdEh4Jwk8Hp1j13yA9ZiLdthO
tvTcmRZEZPTNh1ZNRzIBagQrjSyqAiGQz0Dew2ndh2CCI4nT63vuumJP1dcg/XaZ
FLkBw4SZPFHZt3ADPFfWYOvyN7RNAzLJFFdYcDA6DMbakShOYZ9hI8dBPwqNgliC
HNSh5yaUnYvrq7IcEDhOEgn705OidWCGtIM2F/nE928vblkRU9E5KKcvgj90KbqB
6DQoKJ7TEKBijhqhudoJyEDMFKaPluo2lui519rb3ju4y/3bl+dcNH5U0T4rlotI
l/WQIM+QxVP5RcCHAu96wtncUgPKGcJY5UWKWFgYlAcb+HNWBVA4mwoSnKGuMqFO
lJJVM7MG1EoU0zZ38AlfN5V4hxI/VkaABxEguZJ/DkA19HyTKGJuXzBOYoeC8aNa
DFe4yP3FkWc+7nud2Z93aZIB4+HEql1kIbCBrugQ7e0=
`protect END_PROTECTED
