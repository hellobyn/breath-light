`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1t38Lk+5RsqegPJ2cz34sozY+nKKPi4rVcRSNfP1gAeRGkxYrZ1cbRs34PWyQbH
OWFbcoNjaHIT1MNLB32dIPdZUgmkOFrWZKTWHdJj6ko68y2S2/+M6AJe1GU/ZWm5
+gQnSjydHmXOtxsxVNmZnVVkFy4B8kwGeg97TOksed3BvC3K0W+V0FPymh88I0Xo
IHcpkB56Fp+Z4XH1RYgIqkmKvni824n5toly89tB19WpNq80oXNLK3GiZu4OHjwo
YCsKQQe/b6sLiTtBuRiiag/OpELeh+xXNYZJL5JWYs2L1diSR+D8nCi1Bo+tIkQr
JMjet1lqIXSglg2FdzsAQ2/b9kvl4UhY9inl1oTeV1NhUW9aNtc7Wkpv+xMx5L2+
mB8R1mMSzNPIejlvmVCh1kVA/NpnlhxLI8Uf/X2AJToCEcQjw4VrBEcMwS2LtPjI
QYl6tdiH5W1N6tpWcVfZAT1HV1MPdFhoAud6gAsoZsrzlBngNcoBEgn32ZGnsPXk
iR3gJEm4Tntf1zGXYIqc8XY6s8DmtrgHsElf9FY8asSNbFdRnxfLhcQP6qjJLwdE
sjbTgnCKg+fjvQGha7dg+6zC9t/426KGy2Gbs3fm4H574xyqv7WEInxUxH6cSDN4
/HPWAit2E17FSvTYs+0PzWZ7BkGFXb/tSoXuuAn3FHIba8+jJF4JXnlboITKAC8O
TorprbtxR7InoePhBzts0n4N7WRL1Ud2eIaHUl7hG6pWm4R+MY/whdQVae8JPyaL
gLF7AXq9AsscZletaAEK/JwkpLk97+K027eE7sruNEpkxGguRKAt29gJCXkvpbCF
fiFFKTFFwTwBoVf6NoIRerc87aeFdhkGxEEn4JxHIRy78zsS7G3C2QBitwfC0DgG
9NwUfmaLsutNik32jAwP6+sXC5qC/J/COGc4QDIRo/z96TBDNFsziU0953ZSksYL
R9WoS8rI1shAP0f+Y5DyyEplf1pHH5x3nDITMWFTbXR1gJefoMrvw/+D5/SahVbZ
ERTUn0YWJlxcfNXw/2+OqV5b3Cg3ez/Stal0RASDChcQu8aXen8JctFMHGb2uz+l
MXpml4ajIoJWvqSaMm5Zb23VU/64K1gOVkAPZVMjQEkh6FLT2SDlKtFXSYOdqfJE
PkgVvQL+CJOuDeU7A9O9GadQpUIGrOiAiTX1/++uTkKRgiHiy0QTJsdtQVnRVM58
pOOly+VlzmWJg1I4JJpqMpDfFjkiX4l4zsD0G/Ks7EBudgUNuuE0s7WTsChOa0dY
7wjyV0qFFPAGxqcE2CWTp8TO+7jI7Xhqzh5eIsRy8ApyB0ju+3vXuIy//K6760RX
QEdLpR1sV0015Pa/5kZyeW5dRPgBCWeI42U55idM7B+SYs0MqkQ1iHpxty9fGA3U
9Kw7CTFOZF/mTZFIHhwJcbV0dkgyP8albYpYdL/6yVrzlefX4QDwZy59WJZZk1rK
zXSl6nKEn8uQOFylLW/0rExqO/mjOI5n+sRqZ4eI6KH5v6CIFLrCoddzAQWUrlbU
S0mrFUwOkSQEzcbQlLroZ/7fXb/rfvn/e7dWW/RUou11AJ/hPqU1IbuFLQhS+LgU
ng48MsEThpcWjWqlapnO4CHNWf8VLuZFJp4Eeo/yjREBIZ3EpWaV1KrLruUBvR6H
A89meG1wWf7S19G1V6/C/g==
`protect END_PROTECTED
