`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ob7czZueSYFZu+jJP7lTZygVV3MDLtReQPSPmJbzARsOsyANt6c7EzizN2bpuXPK
EiJ6YnCKPfzEATbPCmFUc6/m05r+44C/2U3EKQBByS7y/9wrjOq2/GVlhdsehG0e
Nvd7jtOH61H9VmPw2WKzAyeGVuIpnJpVAuLr57zGzC6rkuSJvIcXGHFIfuBLUytF
PjwLaWycfL/U0Qa5b3qxwyEtm4ir9bhQ+5X/AqBnlhbBupfxMIEyN69SQbrcmdlP
oz5D/L2Xqd0FBBp+aq8OH7bNR2ZVHptRXBPhdPiA8HHfKlDwBYDcnjx4Jbrzc7e5
LCnupV73QlEgF84cdAWskYmjbuPj4IQiQcJ5/poTU+w8NPUJ2ozyAf2w6CpG77mm
ceijmBrVXYJxaGIkZNbAoGEZ/ggXY592KemmS9T+3WRUetrfa58qXs1H+DTGDY7Z
CJ9BTBQbnXfVBqqRwy/BasE9iw3/ora8d+d68OSMcot7XtdKgQYirfgOFmhT1hpJ
GyEIXf1OkkirUYQaGfRHu3VIBCLlzQOKy1+QnwgMg1G0k7/JYeddtmRiqV1p0D0y
fLzwfBZCA4Zap0TBLezCFZl5L/7rP05cYq56PwjrLjlYDa0n3ndMI1w+fRTiPCpT
NdzNXORspnO4fnEOBX77orwhkE5/arIJrZ7Io+oWZxtD/CDLHMQ8p90yQc9K5mR6
nCkFHLHiSzKYyqBPrW8k40VjCrwvFK/SswspUorLHVTv4NgPjwVCPQK+cHFTifWo
XDh/oYgYGB2PNLuTXH89NyLcnhooPCkleL2oArVtyYPkqHqj25BYNJkOH2tthIBJ
KqTr5McRi0vnA7eAANrJZhy2b2e28YwSLSiMuci7HV1gaJuuUdElm6oYyUSctqeY
O6b1ztlgmQj3PRmTBbTtgyjEw9jwTA8PiBDnT8CtufasauArHzTmg8d+vEnZVpfF
fJdH9y4oIJpityO1iz8rOvjvwXl5hh/wPcVbGMWhCA8wq67IV3Z0YFh7/upThU32
41esoKYySfd3NRw5kDQfNWgrbjDp1wOFAmGzEky1xh0FkEM176nQBb2wuZGkx3Vc
wFKCVR3+SwtEApvOJUoy730+kNPJe4u+aHCyi+WyyhZO+dD7FMaooi7T5Wm7sIa7
E+STTvxY/Zys6LD2vGr9lQckfW/a3ayF00APGNsu3fPgdYzyZN5SadkLPLv+SF6f
U7sUHjn/ZoljbGqv5+suqUBRUHnU51jOq0HB6hQ53zt4RvUdIaSXYdhdq9xfL2jy
y0g5uRzCedUkYKDyV2hNVMbrfeJ1w3l7atorHiE61BeKQIUWT01kZ+MuCtxogpHS
EzqyuasP4fqdfGcra/w5c3aCvGbPZ55ruMEVu0FnHvH89H8sx9bPpVACa251vAAM
wh6exCBmvP4gT3T0pyuXAlrfOBTs5JvuUV0buocERjgp2pdsCjKTva/HIyA2oSi9
NtGsC5t3nIsZ3hujEulTOpcZaJFP+5xCHj0Bpd/EReJFwqpbYVRwktMK7tdavwTT
w2pldMt0/qkQZ2TcPEts0AMKVZ1XZl7J2pyGJMm1GVHX38X+l82rXFg8DoaQVfES
CTS+w3xcn1zGvCke2DyqBvnCxxHGHEDCpnC8gWSxCqhoH6fV2IXoZMVi3pJppi0y
nDOn5KkJ43lHtskVwG/9tfQVlTKK8QTJF6kG1JPnu6zhZjAUO2pCtwv38AsW3V3C
mQdAxjQdDDEpKBakCSCXAqRYlzSmDGiOE5yw3nM59Yk7B2EJ+RI3Z9PjVUP2zu1q
lCFQqHp/8KA5V2fMFmNxVaz07iCP+7s8/1thZChwsmcmp8skyLB+elE1U8s5e206
Pcdfg6Bz0vF1qrMczr0JVUOULWbKGOKOIuu0KCAAl+cvgCMeloWcGZZyu/wkMTBy
cGsoKJrNLfaPn78V0kQrs+KtE8TIaRdvnlFTAsZdWE1+4Ni52OS1V45JflDlrNXJ
N9a/VHGtZ6ZqIPBkh7dJtdalY9OdKtHMZsWpNR8TNVb/c88h0hOo5raxGmUMISVb
pb9qq6JkMNnZGFMlKRTg+qgwKkEn/eM1ZElIIDDRcxXNFARYviqJsXtco6voPAZD
D8f1PL85ZBABrLGExT1iTlc1AM6jenC4YntUzMMu12pqR40HqnIfnRi2hwAY8vdx
qdRYn193JRHE+2exbcloOo2hq9fJKFsKDcQouJiVlmkV5BtlbMsfXrLLNRq0CQw1
aaaq89mExkGBepuy5sXmra1LGWAkqGuqQtcH/nxoGQYqhJlTC+w/WbQCfQmfVnlm
EQiTyN9KrcsR6kmpub9X5ju3ESkbXQLgpA6vcJQ00p3uRm8nyFMFDAKpLUeNF/OL
63qPPPSDBTrpO30UP8obgb7gwecrXKVjMhwtRS9YgoGOLmFVw4WhuZZhMZJE7kRs
iQ+R3Yv191WXajIlzUwxHsS8JJqSF5xO/gf/UKKUrYCYm5ZtGoJl8e4LYS0itoc9
5tji/K2uFQfl/3V49GiJyOorBPnc5nLBLI+h7crX3jmfQ4Q/3UiqdkQqI/t+wXbt
LhyllgiFSfjsvLYzPi/44HYznrCiQegMTcBuyhv6xfuHeC2dYxEHqxw9fYS39hXX
6+zulCNIVWvMllHu98mzg9IMx3f79K26DTpVMA2mA3f/9FY6mq1Z7wnyqPrpmbKr
PA4Rz7yly9Zf0akantW8qpDBFx/9qWFfvvbckMJ/fVNVHq9DJ7HCV+Ll2mlVC93g
dCScWyi2LASk5hk3SP9RmUQ5phtiXqfgn3oO+A4oIYtHPDIPi7eCILRRzlNJPWFA
FSdidrcdI7mbMNQiybNvciciZApWqzFPCULfR/fJY9RRhAO5UH+FhSwQv2yJvjL7
XuzixVWErR0UvTMxTAz7XYEDBrYyiX+2/11CQtDiCWgBQWce5AXQmONsIpdB2TGu
ZBGEl5SUOlMsxpvcSCJRJb2lOe2M/OfzF/VBJcx3ahnCJtnmrQ2JzW5lL8KGW7bL
v0Ki+RXKzwB+xKI0msxwlsn30xmSUPIbrNz0l542IjOjwxos4zvWzZqzYvsHTRWy
KffBiIxI3frzHaGD3aqUgyGrWEUeNJQxGWc3LVIhoVchGE0qyZFgO9BPLVBDIlqm
y2YN8PkvDJuQGs1IftctTnkigPoYl0PHabEnKo+tShdvYz/T+RUDfgemkVl/ujPU
ceFgXxl0xRaIYFp5BVX2vPKknrOUAYmhG1a4/mNxi9noeqaNaIv0WwPC950KlU2A
/iHwuzN82acyYqvCQUZ69gzHO5wiquD+vSOioDLkdgrcskISyZkgHQRnUte6xBIB
VRK7CHXSPSaqjMA1uzSZMS3wUmjYsJrhjouw29oSnViHqrAvAB/FZErEldTdgoDt
oHGbC6BkOPOhFKyu3qq/bBapZyk7rJzLK590BgS93oCIcNgq1U5GfJUl0vwMnw+r
TmT9kwGbPq1ssMhAHALd7hUHBtfb0dEtMQIKV3BZT5kfUqlBfFOp5YQEtz4kaRuH
csy2nFSN8vGiOXCqkLUJgODz+9UVvmTwLf8multkWskvR7HNZXNNrsLCPiNWzTLi
G/mgucnicUQvBAqbMWvZMhfuimtAbUr79z0uv5ohaMZDFCdaeN8RbqA7MLEFmp+D
LdWr1vZ9FvYG6Xb9knwIr9MQgwKvntowj8l1Dd5+Kf3Arn6JfpGMsKg6pBxwe2Ew
J2WF6h1iUJTos5p5rK+WKWfwEOW44WgMQgsedlQf3cx2NNTGReske/xzPyHAbgqL
1jwtS7r8FdmHDyKGnfuGlYSpcFLgO//bSsgrA7aH/x1Os+X5XOYQhYUjdV/b+fNw
a5bX57fDhCdvB0IegG+kxqLS1bJ+3Ea76Vl1jPbgPMKY71gjh8WN9ni7I3UKYRTo
O3QXQO9DPF6Gyv86wvdVl5IgXuabANBsFzg/lnwD2Z8oqZ/FtkFlSNMJwNVTt0wK
amvlO0Aq7dQRXif5V3xgC5mUXhCjYKs7tM92TFFhcdjGxLMfHxKJvjs/sZkWa7a/
DKABcgHW4SMNHk+piXVZXnMIi1l5wJYcyVjo16oV7T4rxM/sbuKZelSXX2ZiFxGC
kgcqAHtvb7o/EsCz6sk0BTfYNNJOuTx1k+1Lj4V2CeTT8c4krD/nNqlb+h5tGdx5
jqQHCE/RBlQGSnPmeYcFFNZR+mA61jcwmoA/BNxKhwUs73Ub/4+mU0+XMkS3eRrF
Qm542OCXX9xcegUiKEvsknbUItqyI0Mv9LjLk6IGJ0/n2OgohiaoUM3vV3Grvh39
D04wp2s2OIEHUEBdxkWxKTMfNOyu/AkjIqCCJYRgYkgbbKhXibnZgd8MbxoBa7LO
6bLOT//tKqIlNJiNDkllJ4xCkEaHXNJEcnJUndkmQyzjl4//BckIlaC4HKcPEPJ3
LkkVfGbDLuAsf3W4527z9o908XovZ5G0wBdN38VJ/mZZ8mpmWL5tBBuOv2O74uXN
vmbGGzQZxhkJ+GRVSRUIM5eCaQXj0fr2fqXTpJcyvBrvlmug0kDEe4rSvEBvpAwq
hGHBo2HCmG6OMzEiW3NydiJ2q20YUTDZfemyTRcbpdrnEMUCpGcDf7WLFp7Jnvsb
OrNBSH+ILNZYIpqNfvlPbEWTELjoCkCZ6YFtSJ3tqg1mQ3kMhDGt9T5UO+WVy7Ex
+65+ZA1FwDiFRV7uZNUNZGXoENrFfE0UVvxDyFuanuhH3QnoYjp97wTP8MobtCDe
CIex9upekzZj0QAlLnEuei7Q0BEc6lATUAXcyfZbIKR200icxxOYGjWI1VOrk+6W
GwwtBgfyvHb1WGGcLACdWoubAKHW1Z8G4ml56nmAATeXJSc6pyHxjRUTxZQDTxZt
7Hjqe1J0Kpp3M51IElz4iNz8HhS0JqJWOrsg53y/mwfjphsGEPwzJwYVZF4suN4J
s1b+EVJJZGaUfslFt4Z4Va6CfK9ZlZ5690LhFkiqGnki55FR1z9/MNVcEiZAoM2h
FbN1OstIviCeDH7lrcZuhYQmel6dQnFML5nzd4jAS5HCwwZzTDtjQ659IVeF8ufd
hCIudesMpPuNWLeesITj/l/Sv6Fk1cdGVgBiOR2muSZQuESFqpTED3pLcDdkQ/Hm
Blvd8RNmqzSDTVUpNk5yiLNaTBp9jmBYifi/+HmRAGlqrgNjHkeWPKa4rEUKJe5k
FyQUAKXt4+o2WvRDOTb7KMggkwmJ0fhwdQV3Q0MYuZA3yMoWANbSAINVnvy9M29H
uCfHWjxTKkNs156Xo6wtezzlZcGIjKIpnuoRJeqSI52I/40rNA9W8HdKcyMYD3YM
MJvJJJ1RnGdwk8aX0X9KFEjEilIhGCq5vdLGoO+ezuvkqu7HtHdfCtbPhGTrLK+Z
9Yxo9EKWiaVf1yJibLaTHNrOC2ounwNzQrdF0iQq321FqJP1Ry3n9jp3Sj25lhbx
eS1ezSDkJDh8tIWfgEW/Jvd3HUqamDgmW+/aAgm95Xp4khmnJVYATHmWuwwxKDpd
DRVJAzX8rcR2I/YvruuXHSxeD4AbUuruUpHmYZIK2rnz4CRCfwPkmgM7p9qyDN/F
f+xwKrNeeKvR1nKSS95kHNe064mAqAIqnPpxVvXg6/nOTE+j1kYsqLibCCs0KIzQ
nz2S8sOdsitgKh4kRsfCe9M5EOnjbPuXPvqPlw+FEK5uGja3a92oOGHnGtTjj7um
U0+oH56voFF1yFHi8ZnwuWYyEwcgWxolJkYky9wHMH4nvGW4cJZaV0z9Cz14Lhsq
4+fs5/paKl+LW1wdtYNwBir0WW/4wDIBW5nisif0/TUuYvSu5Y/4gU+ASanIDBnr
m/xgorAqJViHQ10uo3qtM2YnTWKd5zLUIlDoviHv8EwAKJvGrX2ZYjgcRdWbL8wF
xKYB1jXCk26rwCcrVirZBqTGDJ97cuVhgpkXFcppPEqumVhb3+avORRj7LkNPOU4
iTz8h9m+jybO+qBE0VTyYN37YzAZTBusEEOJhLHtkJhVO87xyKzgwmEigbZs0mzz
2efjZKclzfKkhtuo99i7qwRg+DslMH0aNSl9hOU4B7F4JRAArByuYbUQFhExWOb3
oJiywzrILsJPOmfxqk1CR94MoFPBPPI4HHENBo6oqcg00Lc8M/0CJ07UQ4HCkJHZ
JInCvZeYbXplLFiat+fsTqqPbrTWLdZ7A6m14sIJOKxz/pIJ+TPMgIwizEmxUGba
ndrYpAhLIck6DXdig01Se5vdxWgRj9/zkmbQ6vx4DpnrskUS9/1Z+JekdtLUuuLT
3c0PDLb3xNpWPWHA8KBm0ShDY44uwxy44yYZub+X2hMx9wk1VCrMDaVeQVIgHr0Q
MGNNQ4uwzG4oXBLSibigyo132WfQKUPHEk79sp8VzYQpcviTDic+IBe4OXnpYdOS
w7t5H0+bBNUjpFlB9DaHo8NLtvRAKmh3ym1kRVqLPqKKE51CCZk8Sv1l+56zzEIM
BGgjxqbkloyxzQaRSwPYRw2kMKgvepCpbu07vPtEu0Gp+hzBbO/IS7gVTABdQbp9
6QlTQycgltsCqVLMJsuNap91neaVnB/w9cVifKdIJOzkmFHGYfJZU9FUB8Fk+302
OcVYQx4OY6E9rUQBEhXyBC08SyFM/mRm3XFIEWprTQ50WglCZCj/9z1alBs+08x3
G6dPaj+bl4VS1SnNWNaoj7rX4jYBFIOvwJQwQBrL3THKE5Bo9lUHcmpB+g7OP3UW
plWGiKVtDifD/vfZ8d1IOldN7wctu+XCADGXOubMzQDSi01pTSRvREaTgDZMNDRV
u/jGU9ozMXFE1WWhtQzxbV8jEtW0rw+5bMdaE3PRxEzMOxXFHO/oCgdd8vL5bC5I
AQbeN5DmGl378W1G78Ohd5A0/oj2I7n5Lcyd6ZHtA3sN3kTS9QKfeqL+nuo2Ax1o
v2+zvQqZ5Q4WpTywhPMg5Mk6+k8RbmSoOB0e8gQ2t6azGAqacunB3arcSsdZyw1g
kKsviHOQtzIaY6RzwSiupj8RnUhybObXOiPM+vue+PG3XnWxRjREFxjNmva0GIDn
RVrjL7gUjPg80hDRpZhU6lA3Lphofjrrl8QIXCHnvGGgg7Os6WlPaClCKL2EbTkA
xzOKEundybES284HlelUybr3jwR20ztd4++96dzACluLoG2Sv/uBrrZ64vIRrEHU
BWutIntGIdeZNblC/APo1yvfMmAgJDbNjA8SlW8p8NHlBZdiCH6PGVS+aMx71cD8
vNVkr/QSAFShqk0h54RHdDmQsg2zIVf6ZiVzafdUDATp6v1a4wJjYQSr0ks5yErz
BM7wHDtmS7SWkkMf7b07YnQ7rGFHc9MN5KBFvcm19Mk9NfzVG9e3+OtEMq7d5U/r
ZfwjJizMFiOUJRmVr8tP3TdYsFdLDQHY9Rga0wQevhwENCoyEymVNfCIf2SFxSbR
92PgFM1AFM0/oEYieF0INdCt69HIgiCf9dUbrctv3ej+xeGnSwJWkQyaYoMaC2wu
Z89TfzNv+5sQ1OYpcEEEbbNpcNwAd7isO/0ANqKWJGwspdoK7vtE/KR6RsFRTvv9
pouVBrNpp4nWOsGYFcc+K8lJdDGcd6erNfSKenhd5e0dbrGfOgsj0Y0RZUYvni8j
v10QPR+1IxZ9RjtK0odPLLkJwHYyXFA+a1b4rgitwQhl+KcNN5ttJx97jL3H8Nl8
R2FPorO3JMYdL5ig45PggxBKPGn0NAeZU2Zev6s94UlW0jspwbUVi9Q5ibSpZvi5
pQwl6Zt1PHD881vo1fQ6ZCyEzAdvUfVeKY/ofYnYrZljIDfyGYdzb+DCJex54k4q
SzZsyLJqJHn9VJbAeKKXIXZ78VPOB6xOx9KwJYfieF70yIy84+FmDCU4YzddS6PR
Xyi69BvtnM9OctFMoVfbvLwkMnILa+yCeCrxdtDjHPuZ5d/QpeNvtM7ILKg2An3n
EgZ8P8gfYQyCXr6d64+dAaeXVhMkSXtMQbGfOaEoAhNol+r9FljbRMd5Jam2I+gD
iw95J7ivLtreVcqCOqOqfcYQM6BZO8Y58OoF0r9nI70TBqWDvaCiwHhRBV67SKa2
tw7WEhZfd2+0YrQYXevQN7bt9erqEtJ2V+5EmY645+jZPWvFMyX701KFOVM4FQU/
+TXKmL4slXmcnte/MhMqu7YC7mcca0WOzRcwoW3gDLP0fHIvw3Xyj8EhohJyEUs+
ROeDOjxaBk5uD6FbsT0respkpZKe2B8CcL/JxhspfPDqb+Exs7+jEICR6xP2+V9K
Tl561KnkG8G3mMCtUpjLd48Z2XxyGJqnIwOdEMfDJHJ5Y1g4JdKZglLXPnsKZiRQ
tznHYgMTR5fdp3QuAU28KNfZVZ5la5xyis1Bn0f2qUXG3gOOVnqh95eSgl9zTZ1I
stT7HRearPQ7Bk6PojFjGTH4UepQ4Wyzfm7r5FAra9+ldEEQO5xIdvWv9H6QOTl4
shRHCZFsIyKuyxdslt5BJhN5WTEGYUZObay43ZefYvUCPbB/M+fuZMhAA9d9t3Vk
E/4ezCl+JplNH1KAb2y9L6QuezJ8PZDrEZv2vr6RrBVNDY8hW9n4v48YyZUlnTje
kQk2CxJSmfgeYebxWczMA/7NKwKGY3SRLoiUWEKJpOK/4vtCrT2XH8vETKB1Gj8x
etDBhRTyMBpVEOaWw9/+inTkBZgEho+aZLwxYnjn0QPAhREHRjazLBrZ84VkoMrp
MSkunUnUyXFf6FuHQNU+dNCESZG6Nf5ctvUSBLqUyhWFb8nTpXPQ9DPChkyNTlSU
6ZSTAbAbvut+Twr4FT6SlQkfb/RmCNbMtxV2FkEnD6rluI23R5QyT3SJukxTtCp4
S9Uby8T8287GbI8JXte3IqHHTsopkmDq3WzxjBiQuU7cWiYK645W2qvAXnZlGetJ
UcBFk4aTKIe8T+siOQzlLjR/TDIUJ5Yg13IDiG66+ckVvOed17jCVbXolW7VlwaK
9KRxKcb7A7eq8M0/5mK/4Ot/F0uxC0ZqDb2rgkRP7lRVOeW71X3XBaUIGqIKXFx8
A2gOVYG1g+8xNCGbyLB+kWXDESW6VWnTY3nE6fS4zv02sJdM5r45Z+mKzqoNh0Pl
BSkzrcpMPaoctiUwZFDTNa96sBIrsd5J9rDRepPFRZLE9GfNjRcK3DW2evw6kI/6
w3mD4KwevBfHNOscfUsEZUmr0B4h5Ffy+OtvSTeB4MhBjCclsz5PsGKNgOE0IwVS
J+w67moCzna9M8GVRa2PeaIOlNaBY9f6jF05b1UBYiSF0bKXfm9WvPiC9eTJXV8n
2sJI6/j8JTr72sBCDEmIUZVGlJhHMR6TQgfmbXWlm1oJywS5qf02rTFut1Fe2HCA
5vX6+ia2EIWuysZC9myxlMFiyGMLyfGnTm+la2ocPmfSarAsCNh/NId/uo7mPy6k
XNGCemnnHVjSEwcBVZ6OJ/MVDPAs7EjrvTN2uCfF6m9vFXv1Z+Ai8GabwXiBjBeh
3z4XzkYtW2MjV4ffYHunS6QpqtNIeFu5dmX9FeSbZh7TeEK+lp/bm6Lo60snDpXJ
5cSBLy/YYSuQxT0ITS7WxXOJx2jLVQJ7v8wcxRVKAXnJlsVTIw6Pee/aH2Nv11ds
tTeTt2e96cVNAcvinoMwKNF8i7bS153NNVvpxtj0m9WAg+vv39NC/NVzIa0W2paX
+jWkKi4GZFJDniG9Mc1EhsFwa5cu60n/6/SpnBg2I+wviJYl81hbgv7AIPnPGlOv
fvXcrzytbfn3geemfGxziEJ952A5pkBJAjDKS6onA1A7beVJEKmhPq17mSaEJLEk
DZ3fd4Snj+SlSZLPksoeH8CJuKIjdrCcUVPDCYsts27yXENmKwTlCHRF90be3Xc6
l9oJVwolPGIxxh49U2NDalyAqc2j5LO/1GY1zToOWcdehv2po6yM7j0lpuPvssfL
uwlC2NSprO5XsbFkElZpwAuJ6WjyRQpEov9A5OypPRQhuJugqUB/4Pl/7QPgLi4A
TWjPr4tzGN8d/GDnvaOeATARnu6epi2xj/uPqx2qXTJmiMzqQooCUMPx2yc25aSH
fENN3+VBwBf9b4zsuVyQ/qz/WjLdinTrX/jQ2g+TRW151H4y3C6lzqVVGf+snDIl
oOGUmD6Xf0nBb3Yg9OEgORqsSEss9pOwVRL9VB1iRP2Q2ADiLg6cx+7zqaaXVnGu
CN0plQN+3aTtQtmlacVfzdjMXuwkbhUJTn4AAWT/i0BOszSLFE3JnycjS4TDDkmz
5n8VVLiXiGcIfUlRtw5+U7x9UeEarOVqt5dz35+HENqQ+JDThO/Ze5QzV2vHTV3L
wP5t9qqUZ1219fw9B9ebW6qmE0p/RNJtbru2v5iDBSuJu8h2xHXcFar43l5FZMPS
2WxnGuDnm6YCZD6WED6Z1OKjsL4iXmJ5jS1hpDUQHIjSw6+D0/EDe0emaJirN9aX
FGVNekoD3XGTWO9TveJmfkDuuq2W5cDOTuC9Hh4JvSQmhKDEajoZgtHE2Inefw14
Nh9I8wLGZMwi5zM3cEhCWCWqVguSEwn6bP5p20ZlE6yDYn6384UthzuyfpwHWTFz
bZsqUb0Rovo7E7LVJ5upMP1XMvL7r19O9V7v03VRKkND1ypw1/cmjbQBI0WeK8UJ
KN8I2YkeR2YlGa+L2zCi5/xood40x7vw8pSblZ4IaPfQLZ+tDWVjMIh5OaqwCiSN
H3YR55K6KAe67PawLIqPSG16tGwZPDqQepcBdpCp/bMyF2cdnlbmO6LcosbIXY/k
M5F1cZSpDRsoJrPFjLAPox6tpIgcNEIoZ5M7qMpb++Cyg02409I9FjCPYEdgda4/
m6YYkeKEqLZlALzIgGqDGVaSGnXnbvGBZAZ7Je8VoBwzPnvKx9/T98/6i/DfpMwj
aMbRaLfuqTTW6+ZBP6AWXRNOXNlGomQTl4KWfiVstPkpuRHyHoXlqm3hBKAuSaad
2q500C+kakzCQY1aguc0C0lqEBDtVtRyPP+VCYXi6wgNfWsX75F1bsT1nkkmlTYP
pcK/JYw7CQL8dvhqY/2/GG2MXTaoWe7jOrYfybhWe2C04Jhef/ieYv38p+xFQtZ8
RM/jhL6OJADyM41byI0gh7sc+df4X2NwpeToUp/686dtDWsdxICEb51f5NIi1G2B
IXBr6/LVMOkziCeYu5fd/NaO7Lgx9MMgKAkQ+kgDzlROHKfUKNJdli53e0Lt5jtn
Tf0Gtq7EXndzBeDtSoyawS222m9HH36Vvh9WBjMtQ4ZZMelidLsUB2lqJKXmDWNk
qNPd0mVY2p7IwNTSaTjsRmMekSLGe0mP0ejSy+wBrTR7AGh76+3GBf0OGl93d8YM
uUBzgkpPloksOSV35yJncs7MkWvlOfQq3psX2VztK+zQ8eeSDbLU7d80MOSIe+4s
N610d1sxtlhSX3p7MRzwSpsrx+P8NKFmwrhWjXMub8Ox8mj253RJLi8wBRouBrwN
tpWeaKclrYYVCOH34r4mzxRS22wRpWqhbnJITZey90os220652O4PR2BA9MOIHBb
YLanOktFLApNJr+DqpoXEkQbrm/EEl6+iP2IUqYTxFZ953pTVX4G1AFFPROS6F14
4hiScwrOPs2VG/k23mcJwIgTgfTapDqy10ymxBZL4PWMCquqR0J1pPpQ0NQVLFVs
8JHn0C1reqllkt0vTR6FJJwNuMf/zzMziu/mGGccpSgMX4LJMCHK9Tih1rtkFZDZ
WWRLaibQXYoR0wF0NQcHt4uQmidohNnJHHhbN3VmC0AMG+/MGinwRqolN+CqxUU0
ct3GCKfFc1cnRgiNNrdHjDxiokQD88JacMNfeQ4TFtDwC6+qRz5I720KAkSSbth5
kjx6bUsnIS5ZnMv71WOEibWfEF02+QWQ8vB+w9efhnnr8pw0hkjbJ+nyCM1jNw2r
fzT2ELUKKeqCaYuAEPpTN8Vj4F2iCBNDaIQ4h3wt6xvrxU1jyQFJsGtSDQ/YBd+9
nqzAE5tqK71SbSNf1aRjn2Snlh72eui2xXVprUHg75GJPuX1dZpwMU5hvy7s56Ek
oqmrtx5ighb3EFnBqjxXukRrIDlvKTw+NVZAbnOe5Vh/oTkN7e5gauvFlVJQytOL
YWsfvmWt5tqQo6rxL++iRjD0Z7qoDY1CRYzbcSIELIQ/B3TSRnV+oRBlX+BjQfVJ
BdtszKSrGZIV4U6HhKoK7oX2m8HJ1c7aYweBHNJTWfp6wu1GDTh9JPMG46toTOP4
xXhO6lNIlQG3XII6tSVnkWwXR9lYaRr/yMSFo+BgpXEbXmGL+rs5Zo7akqbT+2MB
05ZJobc4kSkHtvHSo67E2s0Tf1cLzN4G8FDmrhoASou3EySy3OFhOvfXqh0jaULM
Yz+dHqVpLjF72fmvkdK+TI8OS1yXoPVuu7BQ9BojdrWGmWzh//bQOfxPLT1k1uQ5
HkNtvvq+EnK8Jyg8chx3Da6PHdwBxSTXAGjEr60FzYVIj3dQD5Y3+tcsO6ckf8TI
YAcRtO9VsbD4TU6eFtsDg3D8drrtEmLpXeJIkH68zXs8U9dfA7MPF2aksANabM+9
oXNp14d30ktiWSiKitYgLqTCBM/IxlA3EKsvvIjYL8ky8iDrqSk10QvGge5jFZZn
83LlwYfOTBhOGED+aKRWs7kQoXcCrvd39sW4KW0ED6VbuBZMf99HOpGJj8kcjRla
unpTvtWIusknEAro0x3JaWJZuiq8HgoWJVVvOvasVOkAjjDgD7FjPWyNKhWVy/RJ
LpS18kcoZQGBDuz/SkyQJyHv33zco8wsonh5LMfs3FXqIfudqjCGVC3wqVNzRjvj
yJGatcGx5zP5UoBjuV+TJWJgOg7nCDdDK8J05ISg/FET+J6HmaNWl92afBNlgdju
Fj9qxcTHR00swfSBWXz6STrISHF6y/49FS+Es7dQtHknPMliBPDK54FMFsDLfYyG
BuXPGf8n80kQxAKwjkaqqrahrnbYKGuiwJ6VQN4gpETJynD9iYrY3oPYrV+gvyBS
rWaGJ9hsn2NnfroNYpB0pw4WAg/bIN9almVe33baDbKo94UFr/DJq2AJ2NPjzdd7
R/RBFs/Dob5vxyMalRyESG4OsdcPE0L7OGPNUsKjbWnl8ZsjcNoLWX6fR1MdNUV3
6XgBngEyBQzT1R321Qpk7B7M0Qsf+l52FC8uT4+nCHu6yapd+PvWV66UtSV9BbJ+
dPWGlDfh6HrlXfKFasSAB4MvpB/upTmdliakQBOI0qnFeN1NFlxScEqsk5vxxlU6
FYpJLBMBZCw2g+RR25hl2uSkrUTXf3ALpoTwnTA0acVex0brJejWQjIa/NeHpZyG
A8kii/iFcwVd9Wp18hgiGdUX9nwC0CMJNo/hSpRKTzjhzsW1WSJx/tb3iz7nB/TB
fblxZyFdXR3TdowQAQSGXbphwf6XjQWKl1Ft5yWN8OpWtAvKjThXauePpdXpQzK9
3AHDerjziG5zIXLWK3ahSeOtnlhOdS9uujLLKcSC7vMGrM+/TvTA/2KaTilMy8KP
WwicsI9JKpHcV6eb2KBQHlezGsTmBkNzWkeQYHKWubU8brOcCENbRor4xqNUdkEg
wWNh1HlLIFZLzQaHFpefYFg4IsYoIIZSjj79uJY4bAuO//HM1CIRN0YgJWXLU6QT
M6Ncu9Lumib7QpyUIsr9QPce7aW/VCtB2ZKHYHqoePOgnTDcuj6dRf+TxGS+OW0p
aqZBAw4AwLCY6wIWTlNLCp7JL6y/UDDrbzolTX/EKT2I6/dtuT/KbY4vHFfCbojk
37pkt3ZK8SUYcrH48CjoqVwLGovI38YG/t/zwNEWWSHF2NSweXsHzX4brgqgpxnf
h0FCGLHCexItPFAnNqDp6AJyIAASgD/+mijxV+GqZMvyyDm/pLRnTENcCjRipet5
OtD1D1KVx0nJzitcC6a9+GWuPyWafR/wnWOeOtUfB4EQvY9onQqFwdrV/Yr2I+Kn
0GL8dytKpQSnp7bNBQwrmtHqV9CPndTcOAo3JAYYdPpU6lykEjFvZjvBEI++lQDY
3fzvS5r/oiVthTz5SjhO/tbcPMpoQtFKUg2XDn4A2qzneGsQz195ibytXVT5x7mR
10qCgF8FSTTerwX02FoGXcZpx32ycf9GReZZoIWYCKl/rUjTDY8x/gAuNPAdy9pK
OzXkbfPDSWkX6L6EOWAJ5As378eEOaiM5Uy05+et+5MSngf7ZQfb6W+pWePldB3T
yQWoqw/OFrssgsdVjnvk/mjriVbXP/V4n2SJD3kTaN1G6itMmOmtcYstGQTj8zM8
`protect END_PROTECTED
