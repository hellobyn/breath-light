`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdku42FF2apWXk6Vfy7KwSHe1UGlOPJheVVQGRbEtmwjZ3TJZ+aR3wId+bfx0Loy
oCMpmxY5qsmhr10a3R4I+B7dw4A1saUgrldvrFxa/lkksuMDGcreCiWrkrKhfj7U
xy4xV7jFwfUct6TXmPIy1gPuGkZonthnz081+OUgmqVzTC/wtCFtpheHQpqMmylx
Dd4DJ5aZhXpdSAPY/WE7js9n3JAoW9P4/AefHfmrReLHOvu8mHXVyEYQcReitWfh
w7xoYKpL07+3QTZRHUKB2f4E576GfLUcpMTqTyHsv5gDlBoBM/MZ2qQvP9Lp/P8m
tc4gEMxwvcr+9CH2riu+zcZ7aZuqIDY/Lc6VTaH+KeKIfBwVVT2cw1Uw+XpZIokr
8klkbbVKvISaeJI4dmRHhaOjl7rVZMLuW+kLFZI1CY7abI4ACtgh1vfIa9py9m0o
3SjmgRrTFdorSQ4EAl8h6VnAa+tGAnazKQRDQdfS3vtA2jzgzmBGXmTiO51Xdp7r
3f7jn8g3fzPPs1BWyaz+fBdRdPaGzaOdSUuBQJT4bKYRsG8DVfTP6LQ2go74BbOP
yVEloCWc2/ZrYo6y/1TiQUPCdiuGZpgFxUv8REOprmaFWLabRTt6LUH9d6/jp0I2
M/srGoEBCnF3s3Xbn0NR365qNkhj0PQZbaaQy3JXOWOXyU2JtvIHl/2Qx+j3CiHn
LxGKNHnccfGz6/r/ycFWkw6ZJvJPDV8uev85gt/HNWLkei7bSE4ty0Eap1k8DUXz
5jYtP5rryoBACz6rw7o/WR0ArWTrok3u8NQIyhzXQQ+bRq0sAi0cBxYEDTcu2Zpt
mhuBXmo2HiKkiJ9geFBdMXDrM9Sev5cRzvAMbWV7JIqB4pKLzuSkB+OvCEapIiAN
Lpv3dP9CCSsrYZzmmgjjisewaAxXpi/0j0MPgM2uumuF+j4TUxRiAWcfr3rkgOaO
D9saBHrlPTCFrxqpP686OH++nnf0LHJmwGOcOKWBdXSmO7F9L01CL8JWwFUs53yN
iBUy8q5Tq3/FgrZFWTvUlVUjJOfDz3P85zqlA3P674yhdn5AfCFHTNgOQuerSY7h
GD8NxOoSIXbaSwciL3D39w==
`protect END_PROTECTED
