`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPHJPDlTdoFCaD5qXnqfiga0Dk/K3O31IQFrc9AFFYuDGlzF2xT2IthpZ7WoStXZ
SoO6WfFtEkWAT0BhfBrDxnPxo3NkqhmtEYLJ0wBHkhabwQDEe/zU4wbwPQQKIvD1
fjUNXQF8t8LfAILC2KpXUrtEaSmo2PEha+RNXd3TcWS08BdrWYMe+n5VlmvGApVo
m8h99uhoJef6noIW0qci2bXh7X+LyrGKEB+BZ2woPryNW1K7yPABw0p/Z6zhGY9A
Rs+Q5XDdngifhS710381XFKKJKhngj7t3yQ6ewSsIy90hxOhneRnnuev8If3NhIW
flQJtEl01/GEgIV7dUl7NImJMIi3BkJzUFwetGI4A3lxmjkwSjYXnMhLJEljWMRc
e6Xs3cuXvlbSdmfGj9quILnU+u0rl2pXogKAQskt98pPfXNx0Ocfgc5WY0CE4I4e
WU1K4Cml9i7kkson4+niuBABqo1p+/an5jcLqJVG7QX8EK7CvP++A1JGkpu98vJG
EF+2P5fMO70sNDfFC2V9ajPF+Zkc022j5dTUllHuR7X9TjGTjGxMNSpLwVonffZE
DAY9Y80uUcI2+T2afHt/6gU2qZeHjWu2QG+TndtdF7wNezbnhHo0bEAtFQgsFr3H
7iKkpDB4iS5qND59l2ASIAiNrKwAb9TslWV41IqaYfGXlw1+Bn3TEncSp3aIpJGo
s7IaY0QVXC4mx09ynDzQtQ52obceRqjA1PSTaXJmxVxN94+6vXdxKpluRHGAqwVe
BVYe9rseTckv9HV3UXgbrBAb3PnTCCzMgfi4xi8jbiI7dKARXOMjtbEwv/ohMJb+
noObQK34Dy3xEhW8dY1Zeq/atgDp0x+8Gw3pzMx1BwNOQU6QBia48/rdbew/wGJI
FXxH9TZmokxVknRBi6ILBHr+p4oUdAhf/ce+T6p05VjZze4GCLedek4jPScxnr2I
wW3+O2FvsZ9SYHqupIvql92AslDrJqQxWfg7nP714Ak8a1IVSnMgDDXTqkzZMVr8
Obz2FL+FCGj2AyunJTANBr6hJfPDS/biUJzHJYOinoc+VArVS2nIhTO3BwIBg465
gZITl4OUqols0hAmGZa8zCGU/P1VqxJb4G4Hdds1x8M1G3tkkxKascWX6+FfokM8
g8oB96+Lhdfe6Oe8bIBfSdEJVfYtHcOEjFtAVUZg/HiTgxV2rXeo1Yzlh8iEcq9A
t0CTz1OAM+gsju5G2LGUXWsNinPb/R4AqpHlEi2QrV5AIPpkBW28G77uEC3/ZRc2
rgyTV6zmNKCaybQD/QvPBGkfnG1DYFSmlRTo/jr15VM+0PjnR3q4337+xyMGYXEj
B8A/3093MbAdga9d+0DIpIy/XIuv6rvDs0kyGxRovUsmm1plg6OlXzkreQTjpwIm
7MzJAqxPEyfMWtJ2nNFMswEjJDBfRzNoMWAPJ606ArwVxd6eMyCGopo3G52lLqlk
UZbCR7N1/+hhu6TVYY8KJepgphV2cg6h/mxRG9peta+tsHtz7dxxgS0ppbAVfcnr
MeKmGgqtsyE1VcffumSlTv/xOntGciaDBtq3rhOzLmz/A+sVaa5fsem3Npy42wuz
5QOp7TBBmlQPmhfHZ4WY+p4gSDVECfNV8/XES0r/sdu6+qNzy9TUxJG7inL9Xj+l
k758Z5iiFl/3kRi1gynwg/yN8kfJvX610GtEpEQgGQBk4f7ULV31H8EoffvAlvzZ
RGzC6Ls/BalSzj2l9J6pG1yAZnCjqQw+PJK05N1Cs5Ajxuzu9b2dU457JHYmoHE9
H+2lW1wLF9pcQxvn9l7akHSEDwIDfmFF9GDxgtYWI5YWWFdZzPKfMfPSsCt+qleA
D4ftP/wnTlbcuhEiE57af8KxmznFVFavuMQZMTkxU1xAgBrSzq3UOepfb5DZqvnb
ixHDA4+nBSgH2eHwcQxvbmcErSRMIoeHGvB3kcPcCn5zCaFWmOwJbyVzX2YNvW/d
Yso5c1L6JLUHuvqcIRCAhLTu1bq0oGzOl8Tnba/lh2ST1NH9DJ08rG9IUScBc1Ge
PD9VFtLxwMjX0jRpayTnTR2gNbvOF28I/3RWTCgtTTIPug0AT+VtB0jK4Xk02F0t
A9YdiWbIliqgb6cI6W2d5pROXWBe7TcJr4Ya90ADOCG7qQ7ym+wfsq+ceMkXjAnZ
9qvbubmTqe/ouLu0vrErRU3jdB7MMNhaJM2BB2HOmQQkC/5u6UGtlyCjwrnCM4x3
KnTEcNcWa52Ckks4YWxRRHJLk9Bcnloj0jmj6dLoTRBx3tSJw588apnLt0sDglWQ
uYdJkVEZII02xWlACS0gM/UpFohz6FIyVan5D6B2Sow9qaAJalo4lmI0DWOOJl18
qSNBjJVz0EkXLiPN8JqUcMRuZG4dqLLtqzfpIit9OEEIfBJsB6F3K9ksN4BY3wiR
AB1HmPWO/sSDd9qd1gfdr0DXTuceXSn63uxsij0L4AD5nDdbctxNxenqd2oIZFG7
zeFW/QDscbuiRgX0DuYl/3Pwtu07h8dPXvW4lmE2zgpFcG5f10qH0/XYWE1s4QHs
c//yZ/HYbI8bDYiTOPNt7WMnqwItzLlhyIc6zG/0QChw7RbKxpJ0CoAN+7vcc4UE
tX3EVFrH2leBgWukclufMxL0ulYXqxeqDuqaWoG16+7sEs50adIxdTwg2qmkr/uy
HG8PKB66eylqy4gRCL65dINkJw+nvFYQy25ACW/teVtTkDtERnjGfTOPKXawnkQU
otN+y5bEx5h2WSb7FKwcAegVngVtEOb5vTsIcaSXLNykwmUdVg/XSMCRXXJJfbNS
f8HZBrvhBaZ3lBWwI3XpghqGfjZxWePtQQk7llMCeRddROczC9HEf5FcAZNdfgB/
9caUOYrMtwLpCEQIMgF4seDx4ON2Iqt22/kQBgU/WawYB6aRLXaZntwmv0Aw/qoF
CfPAX8Txr6UAo0BeA7QTLwq/qcrP/aquQFZDSRHyMrfjGV4/68MTfa6d+pUN2lSc
BggY5iyU84sUOU2A4gLMJXd+/p+YNMwN7FQpJVELN2IiKHCRV/F3MtG+XAvZ7lcu
gipi1o/PyFUsDHD6XWx9yfct1G/30WOH40JE0MOHuYG1CDXsrhmsrC1qL2rh/nhD
A+R4gLn81WT1iijOGVeUgwlbot+GMm7vFyNKYeATH5OHYxqUz/nG6O51hj3arFeD
1t9BDYC3d9cRgLDuBZWRwascNZgrkHS0UmIu6GAXgoOICmb35tmDM0k02muBWMmz
lSsdF1ovRElRwdTGiwyTnalW5OLFgeTRWD7XXNpk4Yuf9qhwx1fKnZv8XWSZsGpo
vmsmlGcCMANcWStIOYm7p97GvnzWmwgj/xzCeVM9vJDb/WeiDXb+rVGWVxaL9xaE
ZXlnQNF17RXpaHMDjNfilf046+txUjiNiIEuEESWKk8DT4n1Eb8j2w+dS8heO3iE
W2NlgItxNvRwCmiC5dxx1IJsG+GYdLyZIbXhwbXEdPuEcRlwZGbrqsmIxCaNrWk6
Nll6e2rsubAhvm0TP8E54ZKcpebyMrVZJBNkOSffDzUU74tDVKu62emgQnBcbpsG
MZ3c0ktjlordwSQYAQcr++1N6wnkGP24nTx8geZqxUe/d+lLSb9CFFQGZTcY6vEV
YegT0hxI9AJ8TBcRdEXMjUfHS2eeepzndGccSuIE/ZYpnxzqPgmdTQ/iR7QvpF+2
Gw5uynLr21hVFSL0XCINbeMYqUvxx8J7orS5baaOU7J2ZZUiKggAPo0tWm11UrbN
p9L3ccZ12+ZueCOVH/jjLl7Tzwxjo+wr06RyCzXVN4jdxSVTQkKzogM8+rOYBXQu
CvEgDdqWfvULy7BzpG0ug/nIWp2Zb3XTKcBTwS3WKGIhnymxHzH3G0qJ3gFGptnD
gadGAyhw14Iv16yzMSkf1lGnDc16LmY6Dw1NZZdKVawhl442EaU+ZzX6jraprBZm
YKrFV6qYMgwYrDdiHchaqd/vPExOKLf+B2e1ITkPmrGlAkfGKk+KdFUO3cwLieBi
Mop/vHsYQZA0GhP1YxKwdZADkbd+ci+qpSE1VwYD6r3Q+IXSsuiS7/z3BY7sx5cj
0rVElWbh48zXMV4j50x6sX6eS2qQchR/K+hJGAJFRw4ON1KF1SHgceNwK1TLKZ7q
PrMLaujH1mBaXj3kSPfep/oQowlYrWoG66WKI2yYq2zC593pBeUKrPMpxi6h0ff/
qPZSgbCi7O0DBdSozjJGE9rNzYiSGwZohaS6sEHjB1B7dRQeq/ap0wRAB4DIDFsD
/4mF38R8ULzrb2i75snE5usKCCOpFgAqpbqUPGYkeUznvYNNpgIUVh5s3f1VhIQg
5hzjFWNFdp0shPvUa4ET11gLz0342zn1z1bHhCn30WzP3sGQCDOyzDgAZ7Rix76Q
S3VCHVDjWYwNVgfYgWh2xcRzWiuF3g56SFibJcHNfBLGeoOChlExVHjFgMlSpg/3
G98uDwrImGZQrSouvwXyCKe7kKVxcQhadPqi51/KlGy/n6GRkOtakWRtQLQxmjZI
PiFSAR1r2FyuH+ehA41xQ1O7bZNqgh1X2RWTxT/QjT7YEKcMkKP2XsjRpMTH65NN
944fifdjfo7U6fxnI7JfEMZ6UgMbbYaqZfS4dDzltNAFv0H7f+ij2CbjNPPObmis
PuWIL2RpokS1Lm19SaaY+VQA4VUrd5tBifesLLEGnFlDyvHzXV3EnfPRqBuBoIc7
osoi6AM8He3VUg6YRIRIPuVxiM4GrWcDy5MX/feU7NDss5jaQG8IHlARw+oNp7hK
uwvcpM/MwPhvRkMKGrnW4AOIB00UvdZN2Q7cKDw3zDya3kHMxQmSRpt/ZC5AKl7k
cHG7HVQRlpIOJp5A+ImK19C+yH8q2OOabO7917hN5CUcUSK50r49KAu8bc7ou5hX
4c/Q5YyeiLE/OaIkyKlEUhvp5puM0eUL5N++Dv/9GL7F86MKDSwJEOMtvD5IQLfw
qVZ/fqeGtq+WnCFZxZmHc34mP1hj2p4df+u5qHTRvSWfdZIp4YxinUA3NsBC3KgZ
5eKORUWBBpO+dbCC08mlA1aXpbmyTAQzvqUEc7j1TvG+EnPb2CHYliLWnfIVEZwA
mrwTM/ViW8PXauW8Rlsnj1ewUbdUHCP4o9Gmm0rVV9grXAXd2BkReB5Aaw3zRAot
xBtggK4zvqartmNEuM4gCinX7rAQ6DxqpAuUtsEr96NxOpf08hNqAwI/gOVBryIA
S1Zfbk0BnmAAa2mWnv2HtwysMqmaF1UFd8NN9AlGnY20odMekbWLp8qmoOthrHgA
ocEW4t+wHOXG/MZvdRuRVL3qN8AFioonCtbEPvVXcp+PDwB2aL14NrhzEAs2SbeU
quECo7k1LP8NPFuAejWqL/cXcuFfaYWPLrDlfDC4VxATHZ+8MfYWUbtwRDxY4ZHK
tRor7EE7cUiybU12Ob2j/iAzLlmuAqfvt6wOv0WNi4FGcAZJTWEa4GHJQjTMBRbb
6/6DnLDo99lrcETaYIhERHi7dPf8hY0UL7cceUBC1oRLWFTTRQdlw/FWoAAI5vTd
ZXwoGpieqQPM736WzIX2/Ex3oUbN69+s67cUmqI056SwfplkZzhCuKypKlSdRMXX
Qom3DRaYuDJI9KGRXbXjn2UGo+DWd7RToCySWsU8hrF1LlLQuL9aakh/YA/omHo7
IIJRNINiVuuoNxkXdV3tFlu4zIgViQAn0Ad8FWY3izhtYviiqPTMEBlVPvEhSXZx
jAIP5i60lj2YjvR/verUYtBqkwOSuMe0vIfWG/Ssbv9s4EwetqOAVp2hVn1aZsty
SgHpx8ggEPmqKmvBYMBfqlTP8qDDPzvc8e2llLVHgViLZNxOVM+mKb+Wy37Gq5St
hf007PGDsnwZ36gtqmImoa46++8e/9C1JMd1o79IAsssuRcjx04s71nJAVYxuVhY
8lySrdzazUgmlkX/4Jol23VsesrqZmyLUfTWh2xQQZ9UCPUM7rXZ+ye7PcJNRC8/
KcOliyLAwUHmmG+A8XnIeU4nO2PYj5rQzrCSvwN5XCci+h8GfLd8N5Z8yZPMQ9+i
Y40oT8If3uG0t5XTRSh6Q0alOTw8BCYl6gmo2XaX81Dz3+nSwzwupIJvnB++vLFl
otewzy1vmGeuPCOsJ32jOCQoTyNFkwHPMj+mPE3GjL4h9i63JYZ7qzUUG/Hjj28F
YhIHjsIx53W1n0a3mV971LDIdzj6yl1SRHPNAmgHgI8MXzgoEJlOZoySj+ZZl5Eq
sYTKYzqAzymT+o/pR6DUOFaNHjNIdbafHIS4+NAbHk+13frC3mfWbswFk+EeRxue
tyyWUAyOluIVDDXidGk2SJv/NqmJ2TDvoCH1AKDIfEnBAqCFujFDWs+mnuI0bCiZ
TvjKjhYhkEG772blT4rtNHoLfJVHtcGLkXz/TMqubb1S399U0Bco3tglS6grbzV2
7lE5as2QRCBCGWfkmkR8K0Szin4Q36Gbli1cQBp1ziCcJjaupEenG2kHj1yyXOyh
6k/7oVIr48b6jXGra1z+A8dQwFihkKwFophsPa9SnhklAObDaQ51gQ6WHMg8Cs2x
U32rlfmCWYk98q2nTCbvXLsXMk3jmRtthTnevoWCrCPfVHOhpkhb95hl/isW+Ygk
m4uYpB3Hs4rRPmSdwpttvNLWBKh5l9SMG25U/RdV7a8Z8Gjr8sZ0QLpwbuXPnb8m
rllhcII77qVQ1xiaQBKgbVYms+qOgf2bjzXyopQrjdp2xy8Qjdt79yN8K1UMDDPA
oIxcgwd9Sud/1ntHW/qNwiQYg+tbtEavmTmG69XrROsaBoNlt+hhDsRqyYE6tcTA
fHgxA7LRJUx6H0z83ykgNXXXgC+AICTBub63KHuFZFrfefsMiTINTqckIlc3h+ZD
JB5hJrJ8jP3VLyDCsHxprpJp5NFgZmfERjbTGrobIKAHz2wW+Z/usR04bkEPUsOp
RDSDWkmFUDdxnoCV2sPow3imOmqqfVoQ/095YYTcCkjHj1GGcZQG5bQneqdko4i0
7IvZFZey31bbQYIaHF1TiYcZqWkjtmAXikGnkyS9ptf3aYPUKnUTjh0AGINrOo1S
K++tQUSh0VIHcQrT3Ndq1qgv0HALI6ObcnzYCJhfWZWLHJcNKZn2jyWEowg1mnJE
uPtNp1Ka8j2zGRIvORFA8UCNmjEazpVcjJxoLCX90Ukna7hbDMZZT1mhX2YsoRb/
3isIKdLgcLuHMuvSaoW0mRBNZhOBLb1mLPqueVGUDNanokC0Lzrih7JtNbDBHPg9
gRt9M8q/16y4zxejReNlCnxOwpxRt8aJvrz0z7j2vdp8xbYBjJs2yhzm+ZNfMJBK
Ir38kjpEMCYqNtqMihwpEaGb2oU89vLHxqgg76ms5B2FXe+Z79PwCqTLHj7LDY5w
1UNzwn2+nn0g8A6es9lFbHSbZKKFCXiRIMT4Vllhm/vYXlv11owO28VfSBk9i9RE
1q9M64SySRn2xD5gSMaSjsHISLL2V72+e4yqIwuNDvJgasF7az6TdzymYzZmp2uL
AxZcNUqZFKmy6FFhlxJB+mxjPoIPdReATVaW4bwFhzbpuQhFwx4RVPy6l/HSnxgE
cvd5YIdCGAeGviNhPyrE5+QqQgPB27p2avJ25PaXK0vwF3hQV+tuhWPoyDKrvZAf
wOYyvo4JP8BE7VnFsYh9D7hAcCIR0hfIMonkescs9AQzkzi9SBohCyH/TvJVOpyG
5myolNP4ghsScZmToEwqIM7EVeIR7B7n2vdfAxTQWl5/zVzAmbLqStsMgS8LpG+Z
FoKL7znUEnzlOtIePma5XCmV2lKYxJgGUZDsYLn63/qHXodl5HV2KhkKqGg9jOEJ
5aXtkRuN8Vue+UPlposWtNo8jzQ+rQfjVtEYfcHum2Q/G3fVLVtcJ7i+gNH9fTyz
znUqXusIilco4c14WJSWnHJZZrMomXrO179x0uyTfR9+a9cb31dPerqOuhSI0i5Y
1vNaqJHxcIPFwEWeWJRJO2YVJkErHtLFQM49v1UR46geGhPyKCE1rvcrh9i3z5xO
EdQPa5GUwsUVYm8I4Mq5PPLKihgQ4JTavzWCByZpxHrm3/JzkGqCVykAtCwN3vto
daGEOyRYCJjJM4bVPGkqMW9ZomMd6zqihKZVy12zU+uBjYXyJg3iVtdz4weSdAFx
t7L+uWJ5chniN37kYbSImmG85GUqsj/bjl01pU/2c9WF1o38f0OdYx1GHcSj4nu/
foGo15iRc+sh1wFuUtp1Xfkf0e40Uj3UTF/11Kc4oWHLmd8M6sgr/8QsQSiNfFMV
2LlHNUuu9ac+x70dDYHOuEQZm8yliYkj6f5HjvMDC1wvKiy4FRGPVWkVvffi2NrJ
T6I2ixsj2vP7/ZT3kKDffTKuc5UYwcNACzOHrDoK+l1tXf3gZHOyVqwAZKB17jQm
O0dFIVJ0G9q08ymktqqGGZzJgIu53QF5ZCmdZvpnSltgHxpRKdfvHcv7emHZ6WkE
bbwvdmg0emxnGb+iEnE0+uYA9p4TULQ+HblNOJWTlROZ/QhfYleJ3/Zh0aXTcMsJ
pPpcWK0DJZDEHxtMGqb0f7haiJIVXzO0R+GVFHZwKbMQ8m3/8a9nBiRSsOQoSFAe
5Wa0Zhfpd4itKOYSR7VaPoNjNzTKAqr2ngYXW62KU1u/5bMjqI6Z9Y3HMHPvwZm3
gYma1g6g05U/xn2lwWyQQl6z6PoQAnqXdX+MhKWpd06fCkDVlvdIN2MH21ynolkH
I099KLf2jxJfeAQ1zEzN+BoITyypETI6+OkI9A9IA8T1LebYisVHTcPCPhLrnQRa
QAUiKHvOLkiPoOpcp04Hq5oj4T72ou1ZrxVKj0pAXS4Lk/VBp2fftXzkS9Sn6hYf
7IEe32RK8M7z2vM95zBsHFFEkcuMj8OxFj4kB0AKCMZWZc/6q7/kozlXeZJjU2Co
3MqOd8+KLAWr1k0FeeBdLHnaZwjqOf7bd77c0HsfANgnKb+z74+c+bP4PqjSuT+G
GmduWozWqe2EnVy1E9zDdo15HIFwnKepC6psjrrK4hctXxiamDUpOKKgtMAzKqn5
aZ7N37FsgXDm/BHH9axp/vWYrzT9AWamQ5vxZPfmLsWb4A6fhLA+nLcT0IyMpdL1
uUip+3/xFXYUU0yZDYvsfrSZinbeXZ6I3+2Ky6eBHTMJVQdb9sFv2XH8/T6BE7zY
dIV8mIoQx7PbRHKVLgOGkGV3Oghr2OPVKQHwY6ApLyOCVzeqAU988rNh2RhmioFD
Q4UTfxtQC5d2lZXkRmW2z5xQlrEm+Ehw86DWIDXInc3wzm8nZmRNlRZB5YpkalYT
qayLXQz+B0l6e4uOZ1V7Q1zfviEdzepB43JDugKS49JQq87V199KIVbgWtmw7tgg
VHow+bCe6NvPI3lD07JZmVM4OJugaSQoxgVVYWzwo5SNU93R5TuWKEN1IdkuZukB
u1097Oce6Ywh6wuJuXyvLhtOwz3CiTqHZ38VUsADtGgnVZ9s3RRfOQaYjJgphA/6
B8YNJzQ+mV/cRE4C/iLTUp2SFpWquj5MPmRDqqjQFj60J5ouXGd2teSmDBXP3pj0
iJJzhEvx78qWhALDsSA6xlyTBgDKGBqCGo83HO9tNbELw6+SFD6IshKo5pgFRRlI
4SJKbApqXnEKgZ6jiU38L+A/8EwX+Futxw+mz5uW6v0rEcsDoXqOVupxVbQJ9TCJ
WaaV2y2jq2hv4anytZfZhAb0Z1WoYz7A3MIdA1YTFNNQ25x+Ws1AT2RFG6x5+CHp
57Gu4SQyHcLvnDUsRJlo1ji2FE35KkwlmlSML5giwJxeuszXMjkDSbL3Bs6xXEQ4
8uUD/jyN/xB1aRfTR8cpRcb4NZ4+juYtrpUfQU/3p5qo1pCOSFVX764S/sKvFoqf
Pe2m9ONyYLDyWPIACCJO1/SN3fd7ZJsdEmGMY3qHvsheYQi4Pf4doEqmmiIV4+cr
bsDytOoyY0gtcm/RPnf1yb24sxSPJqD3xGVhGFl17DLrnR/BLcn5srhzVoOFH1Bz
zou+/BW4Sz1PmvlYY/+6FzYfFVAAxPQ2cHRMaB6h2qXt7NFMH4rwaSOpz8P1GRBD
asYbC94J+01XZeYrda7SeNu/nrGMrCjwBFNDX0sndOt+D1FgZm1ssk/HxUJcPHM+
41DgT0WqsSY1IbuKDOQxUVEEdA6zEO0pXUtug5T9RB4avDP/ILIgQeY1XMKFkkM3
O8oHt9vQh8KXtwyljaTe4es3YmtOdwSjMN27/Y5jMUpskCQGTi4Kb9ZBAONm6esk
BPM28NAPIhut39RJRxX7Titm4Xnh0U+3tzIquTepwoG6FyqqToDHl1Fc/pRXoZVi
gxpBT3vgGc6wdQjgufUIR1EO9Xq38vMhhyyObnWy9Z0mLg4LtmlM7UOuhKFn05oT
h7drV0RJ7VfWqExWmwGnBdpRoWvb+98X9DFgRXWAEhMl8dyol6k3Qy2+cCOdaKLS
WoXLh9A03yEzHOzTpX0nYdpSRogGDDwtMgJgVLUXWHnEHDwWXMElrGEbhXj9fgZ0
4VCKv8QlajIY/W/gupFqGFMP5UPDsRiPw8va5P21l5KF1D8Ju8kR13/hElai9m2D
Ba1mzvaxJPX+8at8RaQiAOldevthfCARUpOlWG7lt0Ecfsw4XL4mHsWBaeGWFL0M
BzGzVxojnJMYnghMeC3IoBA+FYzGSqr603M3PLStxmN4K5By2k8oClH+fF1BhzYI
UVbwro7B6jZsj4rtaVrPdgT19CkPeh0grL3Hg7uThCdV+tc17ieGHvE2hfvfP0d9
fxjXSUCRGmBisr8KTP1VDvcQk45ndvalkoxlQnBhJdPQpf+i9DzmFXiE7ZanFM9J
aGaGHst39xUrAXvBFrCsU5z1bp61Gk3+5vk/N5kdTLuH+nqM8+jYV5jNXZXYD2JT
qjAgCNGZ71FvEhvxmG/x7V/9vI/3PanVnydQRX2TpCjG9Y1pccsAS8MSyNYgVW3o
zQFq1JihFnu6VQ6sTVZPPJevAFjYrr3s2uJVY8+TxkH+NCChjT5x9qjnxUivutwJ
DXo7gAWCniGulHO/fIDEQq5QvvUPbyCNca/uxgJoIxeoI9Xx4lUQ40ZvtXqiKFm5
/Aj7JElZsqKR/ZjAuimR2lWMIP8DTq0qxCP1I9Hr1WYdvIgzVXSVki0Dvn5Mllw6
7oblFgIhnTdKY5ChvHAVUGEQh+4ESiK4mEtVsqtZA1k6zmP82j5oWMFHRRsMJGw9
vCtim0oavpp4FKUNm37Uz0rT4T0RCzNvwPg0WjLRoio92rYHEySGB2iJA+Az2la9
zPz8EQrYt3kDAVyg3hsRtv4ChXbFk+WHiFBf8pBzJ9Saw62IwKACwdbI7fEgbz3k
RtZL1g1Q6DoD1mSYQTcrWbCvSzvZBptzzJMTf3tfiCanc8JEmmZCXKVu+8S4hXU1
xKcvb0oEThXf5/CeZ9Xw3UPPnB+GA1n4pPbhRNA1gBVYsbx50O8kbnWYIWTxMHRO
a/Vy8/fNMpEsrBkbfYAm88lvXd8RG7PLYkvsNrPwgt2DlDCWFe1v5QkWfiAZllEN
rzOLQAJ5+Q2u+RASQ354Ftf1YdqoOzFXwnGTmQOaERxdahM/IpugjIbCHFEJ578f
b04KzVNPY//disR6B6OEX6UIxpxy81sFZCmLl5HjocSFzUHvHECF1dqNzqmOiR+R
5EpkGC+lEVQlN4AT3kRyIQF1dAkjJ6TwZZOLik1waweqW7oSDHjuX5ruye+/FywF
Ggwni2ASt3D0ZvbOdqFti/hf726/pT8UnZtGZkUY2W+2/7c8dLJf1GKR/impl+Ju
Who5VBQ4j33NXARtB0JWFj0txD1i2AaekBoxJwi3J5BIKkhb9OCyDgunxK86c9vg
K96eOaOb+glYZjTscq9gp92ZSOM5nrZtNMh7FOnbruB2EpOyV6EVRYwr5X/kplLM
a3qTm9MovVFpPFsRN5XO13p+7mXYP6NGFBPYMY2yD3BA6kelklvauGzN2P3xfUeQ
AY16Z4Hj2vu5HFUrnfZBhw0nKFpWIrObjtpYnwXFxTQqErkwPtMxOekvGFEIuB9g
+aM/+GMDjuTdg5vE0sgWiDU7WoHi4A7VXQKneVFWEy1qiYEqAhEc6piMlyxJCwv7
0HmQEUWUNocf5OGk2W5bwgGepts5HPUZwFmWlGxLVPxKBUY8wIIQTulm1ML+9sTM
HkHT9vFDOHB7AI6HnV3YSu1TO0p4fbKO1yI+xCDMvbuYSiGSgevekVB6RlMmvcEF
BNHhqV/XM/L/lapNYQG1wdJGgu31qprTizrA+E8EA+DBxEmvWO1vIUJkvMsUMYm1
rE198JqH/Efky3PX4GWSARRBPRp7khjpJGwd85cDu9GBjYmIIqc6HySY0ugz0nhm
22BYLYhq12Vzek41b3WyWqkznXwUq+APDd6iVYOSUozkv2qoTPFcGRQ8FjJShVe+
16F1dw4MRpVtlduWZkOKCrsW+wbFRTHbX7F99gEhKjNj7DC2/LdbJlNCMhsA5Noo
M2eOZ5F2Z7d/cxZVbdDnhZSuHxfSbGe/uPQGJ+fdfJ1FMsLxrzJYCWZ0hzlMJ3Rl
63YXGjaU59kBRKBUQCwuIWj+bmEthy4VeC6Qo0/Cpg3++qtk6kBBBAWrLPgbUaFx
0KUvqLb+P8XSoIWYL6vhePfvf+kvbXJ45wwwECISxPHDHgYLbIb9FC1oeHiwC9pG
hJlURMZe2LQkbg1q8I6LxxVkzF3BWxY5Wt4NLUz9+kHShMAMiXPvEdcNKcyrfUpS
ze2vAYdeiPQSsMsmOBLogzKRMq/EcLTtkfs6El4CGkREaH1dwFG2+vO0qxUkLwLw
ow5qBivg6uWjanH6/C47O94HJcjArT9j2AvudJ4adfjNqLsRLrRwI4Nzn5skJLFw
8HQBuN/ZPsVfcu7KMSKZrpMPqkfEY7a2rCGjwKIjymTNU07ZprbL+M7Ux/Xf47YU
kRq7Ycich/o6GZXebYu+tvUPQqaxwfBb/gfWywBcHwCXKHza2JRGpGxxl+P/n1rc
9EjWUaz1aI1OJ9GALvjQyT+7SCbsVlVdRbM2hNlI862mQ4IWfNvDevO5zadBsv1R
r8WfAnyucGbcSI72a5IUYcFSlYSrINdJfRp5QtsjCq7RCQVlVtiWaoIGMp0r0u+d
eYMXSmuTp0R0saCebVexUphnqNAUJ22FUfqAAMK8RujXtTPhZXw5jfTbYLSl2qM9
d51fBph+IE2XxvVzKvbJlqzCiTCbrf9HF7UkQ4RbGD04Fgtm32srg3MrfHL30POT
rs9Y3fogJOX5/zClugHQ2YcP835AAIyvntANC68OKAuO+4HgCZIDiLoHKxbprTNo
0fOFR1W17rwJ3DlcnrD5fNVJVG1NEwGgMxcj99F/ALkLGLpUU/2I1MHT0CpmBo3/
3lSobNEfIlEfZUsEIOWNqp0K+Hgu0GPUDJihtvpkTgYGDjMXApp4xfzSnaaaeZFz
GESZfH3iwRHbuxzBOAJBY+mn3pH/hpeCzp2xtXHm2Q4897VLUiwlZaIyugcaNJe8
+Hv6f+cJgYd0OzjmCAEU6nf+DeHnmPqBrFrC4SDs9XMvJOPE2XP10N9wMX8b/flD
fs+OI4JdGph9R4QdD2cLeKtJXJ1cKs5mIPnxrO+A+S1UXQvu9aEnbrLQv+7jj4z8
SqB7keVWGUQqJ6bbcQ8ai4C7ISQihqE2LmhdLH0EGU9aWfZSuQkDgGs/Dtz72MAy
q3bM21wBTBeVXWbjfee9P3mYJ8lmKV1sVSxoCdMTznw35iwSTzFuXwsakBl8uy5j
pj1FqSHBNEjy9c4kcNd2cjQedp0aqcYt6jSgJBit0ulVhMIOofolQIhNxP8ldZKp
MvIL2Sdwgv5VMlP54NLLREeUCg8rFkMalq7VQ1ydyHeZNKBmG2xJdVURqPk6ECp+
+6LpB6jUaFuc9SvseRmti4P8mqjhqjTY2imXGWiEGXmcKG/9JFUKMQib4h+DLC9P
PL0BrUrCxaa5GZEe4289NYdDRuGsQIWYFemONcEBIj7oNKm8Q2xfjO3/ueHPixNW
Ej0VXuEGgAwt6eturUH/0zrylQd/QY74fA7AkT9+REYzxESlQn3zzkRYUx3d3ZUy
a8DlR67pT5FWc/KI1m+3cGpTFt84aycHJbbuIGudrdtbndYGynWzPSqtURAebzot
Uc0PFSEZNtV1g8m9R7UFd7U8iq4TdxIvtIBZg+tVokarj7zGhsFuDdPsXARxs4zN
Ry5pbqkzQt98HfTfzaOdPZRKjF9ppFGz707a6bejt+v51TDJm9Zw5DOSa5nPXCoM
lpjyKah9b5PYqoWZBytfzBHF3wF/IHoIyfYrYXSEpj8nNlAMltmAW8Ef7JQXqk0n
R7EZsB9YUhA2TwWwAyBbhPkfx3Mctt0QGcoyWqHEMoryBj/Iq3TtWKVVQKKYT4Rx
3RpPyZblWcGPAT1WOyPYsImi2Ikfta7Mvf391wE5bXwhPecIiUkz54ttxWnKMSBK
DVzJAJm5vYbGRQFEqXhQp+efAAm9RsOAaiPJLLpxqDAssaj2WoxRzb2gegCTRcXi
AUzYLh23m90d/8ifBd1a8PNKfRAIMB27yYfNkrOVk7uWfikzCZzmg6R06t6W4nuK
40zqS/rgeVh54MErvA3FN9rX5gVyLq94Shawy93nGQqNFALPBioRpGOQ4DJMfrky
Ngm4rQ954EkheiXwokEvIcd+v7YaKKTuLBIWPIeVoLc1itVZWJ3HmNq1PKnoceDa
6VVlSmZtH2Tz2vHEML8fnO5731OZVzOFCbiDKzfY/ctYsZIr9oFtPYGsgxZW1Tb3
xXWs2ujEa0NGyK6W/4DmqqgltgAaIxz8M3b8nrLJEFvD/Qc7dHf+LhIPSdkFCymB
FDPJDVwN31OOxEA+Qg0HWbpbK7E/Q5m8npCiOOGt4SrVaGv9blz2Ut8NRpHEcWSu
HoEZyyhNont/LmvHVqpNe5rVbL65Ht45bIKCESSKlY4xE82hWBOocPCKqLaDPJNf
5SliAQrYY9b9gC0WaMgxm2DYtr7eYh+DagHn58kfu56fNOAcczUEGHWzF3/WbrUg
V16F+QpC6Cch8fCasZEwlVt4dT8povNLHJ2/Ui9C5smpMSwZiMfL/V/OWIsv33TJ
3PI5TckX4mp18PPFtkbfWqlA6GZmeLqW5OusQ1PjaWyIQhmjR9YAPn5d2yoUTgqO
b3g4oalqTupXFFpS0J5f07dFo+IWFmSpUTLgVru3rgtQJamOzhQ6yD0nYWKzW0dL
ZJ/d+2t3KpNDiBFRh9a6TgWDaWQp2Jaa87WWNyPmEearJzH1RNJ8Eq0Ob7kh6vGl
opgzW/Qy+RVMEjVyw+qHVS7cONKJoerlIIqkqukxDn8vN9ZIl5cKDqtTSUIPztAR
AhMkj+/9CkKhuskCqtDHDHNkW/hQBAlQ57wKuC7SpaE=
`protect END_PROTECTED
