`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inSujEjr9RLYnAZmmyvJcsdIW6bvAOJg+VXXotw/tGqNNX5REEoZPgaPtUZbxMY2
xXoeh6saAkxIQpk579p4X179vsx4sPcXR0JFxMnkcZKbmCeYKWxr7ziValwqKuRx
vZg3JPfbBzabvDWL/kAeOqGdfCWDrTW12+Gfz5rQVuH/a1eCVMpw5e+BXwNAhVOA
QfbjSCoHwF8fYnVefAYuQAGmBrH3C/rrVjSeH4L1e4vyu530/AsbSfhWjsiFJvMd
HvK0tdMpy0+SXN2aAWC/kEfPEEzz9m4vDY1buaHTcWaWsvgRo8AYzFpIO4wbr77j
3jbWrQTJGmHK2jKmdwj1rG8E7ne/Q/1HF4rhEYCk4ibMjQcVGdtDg+z1/nPnHfAA
un79ofpwmOPcZF2O0WfinDrOset0trrhpcHMG5Y5M2hJRgDaovxT2wqx+xIyKpCS
4FmSI94cG1GW1jm9g4AXdyv/QxMacGVVWFzCHDeb8k+BYQBXoVbu+cHBZWCRc2yJ
ZgD6lMFDf1UoNJgiFjzw1CCOOqUOH8GVO/LQgcBujbMop92nEzm2g5g20UJcasjg
7iTE3TJJcrXAITh0EQFeHg6Alkhld9TWHl9B5BuSJSLqhfExvwGt1aVmwDux/kPq
DDY9ZgNftmGzazebXqw67YpkM9+bC055glJ2BXFgFnDKHYjQdrQS0XG/GxB8wMnZ
L2u4H8AwnpRnP6/WmOeOT2CXj0vzLndgGQzr9aXVs4E5lMMaVuZRnfI3Rek37Yru
ifIRLKjTWRhr3BAeCchXnvzbe7LTU85S3ctWRHTY2KUHf4GprzZEMKIUjpAhdaaZ
A7VTpLanWbzcXYE2CVG90eBiUsu4f4KTGVU31FziPeqEaCgkrj/kssLjOp8BqHzA
oJb7HRVBIT4dx04FbCdS0+XqUfdBVTABrKhRgS4DxOo935TvSL3AIF1Xwzmj0Qcm
zXO1d38sSvqPF/RVTDoLucpzeansm4TGQmGkmhM+otuE3ND8hwh9+GKrEvhFrA70
eIIm4MMnzcxc01C/RvmyV/u4eM2Rky381ZuTrFi6f4RW2iHsEro0nl3igQt9CXAN
7LH0QYNxmhJUqj9Y3qvWE5g0I9B84l3Kw9uc8nmel8sj8/tycnuBfq++jt+lzIbJ
a7YxSjMEyjeNkM5vWXkaGLcfD5hw5quo3gztzmTV4lcs7mAA5sXzaqJp9NnYb9DZ
RIxvvgUFzFxxLfimhwGH1gvZSlnybyGBGNEscw+b6cwXh3INUW0vj2ygeQnynYyr
RZ1lDFNpm5DuxK7uD4aUxOsu5GHll9JYs0vGd/JSjufcXXrZbhezKJqywxTAErOI
7DZuI5Cs6gsXaCkMyy2jH8DuLIuVWhwh4+lIcq6VhQc1XNAJQ/GbvhspMO1Gc3MA
D+2vSyRUStpOTeYGAz/R5oJWChENe/JYTigEcWlvZSHh/oYi5DYxPcEr1uugsby2
/A3c4rfEaekCWck8EZ0ddcDNqA4TuyUwqBGNkWdoBIxJzfY4wPpGOdsxPD/klh8h
Up7GDbY3V+3A1Vf7/Mqazk9pdpZmHRpO7mGq3uWeh6PkRh6Y1MBFu5HoaAzShgO/
dAb7zITL05pFR38cvf8CY9isDRK/D1Iz/NBnkZHDEA5ZXmH9yfyQCOy3tcUZI9EO
bWAURj2wphXeiwaVFqQRzSqakzZr+Oz5TpCSsYIaXJbbVoAhHjHDmi22SNILsCTR
VFgRghqcA5TF7cf7El9XHnbc+nvsQ1YDp/BKb8HeFFtesed0qCu2SyTii5y0Y6w9
OJGFsjvZs5dC4nM5nPXMFiJ8Bg2nKbv0pesVcCMRGWjSiNoy5fN9GUsk5GGc3gFS
HB9IKPMeBrf8LHdk8LtJupzc9p0eCDRGgdsiCzN/YNLrm+oGwJspiEVywQWSosz9
jKn8QV11HLZfNR84nBoMS2yaCGgs5/4Vzj+VnOTWR+jdzEvHAaJ5KHVQmtuwsuqU
JHRfHK9Hjyu/qozAIhDCf/6ddmi1eAYlv3higV9GUAwfW46KOeNq67m1jl2mUCRH
zUTH3riuhnQqcMoMz/h9ULQ0qz/65mYhxKsDKVbL51eoxoZ00Ve3v3iEdZCK1oks
I3DRLvWePAYv0xtGhPhdBKqyuDvP4gu/e6Jx+XGJAz1wWV75Qu32IwuG+Z38EVcO
Y4rKwdkTIh4C8l+0baBi/BWspiMe3fKjw2NBsastnLrc0HZbCIBQRchaB/RV8+GY
FEhBRM22ow9JmbSG0ahJBXkBuNcmK+vYreFbSkBo66BrLBKYunNL+VEmyJPkGQ7U
cUKhYUTox6pWGRWncp41SGeF1VPhPdJHUf0mY/ektzFi9Lg5YXcO8y+Qll1/FuzT
Ov6V8AdVaw53hVSU0l4zSkIuY2rvHOPNaBFgGoa8BIXoutCywO6dQyrimn3JzBIg
NczuGF/De5Hynuis9JJ3ZjC4Nk6lKxW08olQnaHj2FjRhEv956SyQVM+kKIzRm6U
0sgVWyZroFu5u/4Tc0JHWmX5UCacEZSvrh3p+arfJksyUOYJRGqDE0F2KwMEhhxU
cXmYW5/K+sqNOOLXnSxD23rqq0If8T+3bXSt3MDbIfb/zQLVYMUETK6P3LA3A/oG
/xVRQwbXgNft2jAe8AFrZA4+wSHjxX8xFL38PPWE2H0+HJy6GcndoP/7LIGXrS8m
B1fnmIWUjMiS5e6w8GIy3JPQJ4s7yU8o+3X23atetJeoHxkl7Tv4eLCxR9x4IF8q
MEAzhHufbvdEsrwsef8XO2vJnX8CzHjbOR/HMgxpUVy6Tek8stcU+eQgsoPsGu5L
AfMt/Ko2nfhj/1pnXQUKhE8Kvwjf0kOLxreKDXZmPFb1ppl7mxt2/9ET9MvjABYV
b30LJMFEuYRgQ/k3htJO2k7CzXASB+RHxcbgU74z7uMIyElYf5Wlo8G26s68zC69
dLnrXFnOxQY/UOGNQFuO1FoMxC+/3ZUFi42L/x/MnuDCvdTsoY4wD+VjB00Dqgwe
sVgisWJUdDC2zHjARbnsQQ0gqGtPS/UrokugszcaNc+LKMPbaiqh6tS8iuMB7aqo
ys1QRfixJKad0bsWlwwoEhbBZHnQYCOMiD79rA4MeLS0JMRiZVtohovNluz+TMyb
NvEdHukgEnQa1FngpJjep1u6VbeQW14kTCDV2yh43/SR1NAUs+v+d+Ux9KtlNdV0
C/1+A+R73jXuLqhkziUaEMhTc7xZCc+eLRz79Zs2vK1yIxVJ72/rLQu8C1jS9lgP
XGiyvHiajq4PP4Tv40S6tXRp1mwr8O7+4J61hfC775VgvbCqhwqqs2XYEzMKHLrc
qiTQZxCt2wjZwzvepv7hcMQ+64UOYyOy1Icyz5A3qDiL4TwfIK8O2Dd7QA1eUqyW
j+h1B+DQ//IDNwRAMYlQXZM+yXqusDQprgJfTO8VlOwQVBAm1+mctVFmwygSpIUf
lwM9odrukHBuusOWPoJ5qkc+nVvJeEIPqAtEml+6qfuH+OyhzguESesm18quY3vz
723Deu0z/QeWxWgh/dgSoQbasX8Wrk/vvVk3CeHX5O/d5nulr5D2nC4t9YYHpTtC
F5sFhJzWGHiuXj29dqT8GhNYo06RNtWIP1W4w17Xkm4r+jBQSMKCpdlrx8hgj4x3
yQIMd2gav0j6gNAIoxOdUpHwy9+6/SPcN5YaFUPMKHX1V2Y+4T7mAZxLM4YtA6to
`protect END_PROTECTED
