`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UeExEUxkLEwBRQlCPfl2pExvK5oVPPclllinMFwc85RnyhVihcGSDCf8QOocab6I
G37CQRYqc3/wkHQ/H/sLn640upLyJHRL0IxlODJZ8f3vktVfA+4tZxPWFSq7JC/5
P/YLixvMhGBomdEQn8W6VSod42VWbNXeIi/Tfu/TXmUnk9qz/Dbb7VTEdqvw08Ra
Kvze8rBPhUg1WCjGudAChSJCYgzUXjpORR+VveewKqBu1pd0j9YULgizMoCKIiot
nQOhdeUR0Ce1l5EFIu0YnZ7pVbSMPT+q1wU7ZRIkvgElbN/5623o/zoVqyslDLuR
3jHtRKph6xxxass2uW7BmWfnkACAhaNSf+yLB1z5F75mYoj7yKbGafPvEqY1uiDp
ziolYkeO/zCPvvSqmIbfV7kcrG18Ur/vM0yDCBrNf3jmR+i5obNcfjiR0Zcq4BfZ
fV79h6cnu0GZ9trBEBq8O5/LkCtYVuXOO0yNeCuSV3mzZy/vr4lsJbKGXke6faLD
kOJ4pduhc9x6KtPhST4RW2gDq3srstuRFyKrLeuoyZHe+ynI6Le4h526y/K69/BG
lgsLiluch4A3JfmWnl2bZT3tHWA6VMXLPItcvAA+10z0pB+ftYmeTLX/7q6Htfiy
jlmQ0mxfUBCqw6RNDd+P4LA9qHB+Ew24e/9QShdvaO5l7snrdsvzuEqSUAzSCLL2
RyAlncwm7w610gSwvqkWeCvLmZXiP6CNY0r40e57+OXnSZx8KbG5mjjzOr38We6X
xUnQsBtHYIUMiTPDECig13TypHAmRTgDU9ozEyhTrVbuvq0y1Nf9F73gu8DrE2dD
HuayR9Tw/16jtIAgUQ68y+mCSLBMvqmTQ0opcOftDB02PapCj/BPqwTHyCJQyTcP
JFcZjLKS+7tfgC4NbrqzQMKV7fFmKyS2Zfc+JKaeOt3IbBPRhNgXlyTWkWa1nJ11
qpqi69x9CHXDSN1ZPWxyxoK2NNXnWzHWc5dYubVXkw8y5cjgGT2XaUD0faJLhvj8
0xgZqEhZFZ6SskC+NTyisJVcDASTniSCPlorvL7Mnzh4sazdWYpbjL1KVcYADnLh
ZEzSbsZVxgK25Do1avFOO/Rba8FGcXB6gkQbWhd4sBOPFAhRGQ/8UFQP+AS38y28
zgoDA51UnpBNxU3ptIUGKGjlnSnzNvKYxMkEzBbvPUlHtynP/3QZi2RisW51eZgI
u+iMGbjsHGlLah7CMsLyhjN05r9p2XZTGSwhSzZ0GjHvpqaw1kx9KPpUC3YD6ZjW
wQ13Kr3JJ0u/JPu4f/8I441NKfIbG/li3reb7XU6u4iFzRgQUEkmDV4q3wzP50Y9
d7kdhCXQ6N0O2Oq8ynLF7cpgXG8h66xt20GQrrPWwiGIdYNgVSAt9fudJsQh6gUn
Gqo6cy38HBYhKEdsS+xkQcklNbjM7RvLCRPOL/5YhfJdKtvhaaxYrZ8HZdmXhBTL
+gR5jRlrTuJxx1DrBgWhcbb1dTzSB7YQVowvJKUHKiXkFPeEfycUNBQ+oLoXTeDR
`protect END_PROTECTED
