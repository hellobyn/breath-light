`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6i9J3lB0/hY4VNI3mmsvCznGRs/t8UwcZ1xWYc9hXkvGvuLasBTMrAjuhSPJ8nW
I9Cesj7PqIbntKUrpH4X9H0K1ahNkR3rmQk8zNDOcJhrRHVdoRPBbIaqkRaSXEJq
aZXWnnym4dyrjAVGl3f9ZuxkCpXdSFcANIV7CE9bLSWC95w6D2NOK8tF09slP70+
t9M0LWIXd6X9HM4FR5+SzAWnzGXtbE+a0lofNrMUMPkwc9t5kDpkDQqt9ujhYiZl
PjNCcWsGwHetam2mKiRSAIMs94Ztxfwus1/TQQVuVi+Ln2tMG0iL5OoO4LjNsfAM
HGPq/KmbpCicUwUs2NzGPI9DvmanrhR2dZ98cICaXO8sqUOXM1W1Aiy50AikWG9Z
MEwcaFGtqqoDFw60kk+vY1pq80Im7UV6uvExk1I17+JBwQZ0VAUiuyId+t3kcDtr
n7XwnqvCdqpi01km1ozQhouteyGcxMK4snmf3nTNHveOPdyqaNy6fUF+lPPFcaea
2PnlWl+R7geXId22dlNCld5WO76oWH+bRjuF0H7hZ3+t4O+VWVacoxkreUCIn+QO
9p3Cmc1smXZePoavCRCJ6sMh06iI6KYnv+u69uEa0zvj1N8TbgC+3zf+wddSzx6W
od/Jf3GVqG93iZ8PbJsfx5fxmwMG3/UfqWLE5mRrayowE25rEiK8+fbgoLjdLsCD
2DEwma3szXhuEYpdO5lB0yFgp3Gl8k/p3ejnN5AZjqO0yeVOXHUaWKCFwLMxqDCx
14BT5EazjEGEIA+Tdd9FqsTObe1qftOggBFdi7OiHjAVuvZRzjhblv42JTcPpZNK
rsX1CO+oKFYe7FqJ4S725iY65a/cK/tlfaLsfHqFY5U1jJjMCGmBX//Ffl8l7K69
IBzOG4ArgDcrZltMLvcsTjNgP7WUjc5i2I13wrrgQHeua/yALgQC0KCqIoyue8Pm
Q9xcUMLpPVI1rSUMXENzUDVPrupm6aJzemwDYl3uKLZnUhX598U97GKYqyP4ay6E
TGnX7ynsFVSHCGg4gTobvOzjc/TK+ImJxxolU/PqoC4jLTwGp77YfTdpIUpinmCl
pCjWWJzCoU/iModTezeCxxZ4jsvmaTBvAhSgckOH+g0128odx2+8tV1tk6c9z7nv
kAfZVFN+tsS569Kwp9e2wgcTvNAD9ZcMYHx20XvdPYJYmEhyUPjSc1uxvt8Qd6DB
SAhsRaH1bM0Ppi1lcPLnJiTsFXlEhbjE2Dvdek4xRiDCLfqn3k63cARrJb1v7T4w
gpptgtjzas2l4SMnJxOJe04S0+MncOj+o2dXcSpae1PlpGcvIDmX2IStaAh6bFY1
NFpeL8Nxqd8QNsnp+4sVl7pjnBxW4UOb3IjEkvDQNNAiw+i+48qZrRx+8Qa3EyBN
HBTUIWs6deHB4utAFRgEipGrdIrVy3v9xsKPbMjKwc5B8aUpS00Up/bSTzGPI7qU
/NrPrMLUITJRoctjsgJcEBGco0VxJ2SCbAmCLptZs3J1HpMVjzepwKZ8Op3hLXIa
mywSS0agMQP+hC+GUMHHMTHExExndBEUIV7RmdW7NEUoMiaoRIQBszLTgFo5d87z
gTASpZ3/fc3gyr5lRt6Qz8FWCc4LXze+5BnA5SdKpc4e/zPWgoCIhCFW6taNtQYz
cWf7Sd1HhtPE0wJA6zxIIa+3+6d2UqJYAQtYrCSYOEpYzpcOYsckp1M2Eq7n+eyv
LHtt0Ka2AkwRnRAuijnCN1dcSu/4prjJtzkp4g+ShvIKMhl2d1X9lLiG71SmkHxi
+Pyf6SNeAJJpdZUCrO4GMYRUNROD9hqpUD/V1sdqzziAXFjD0Gfwo0o9lbjtGmuI
4dSRnQmm5TSOt4+8aTWaKCd10GcQ1XNxCXjon64nwo68n/TVXgCy+D0yqCQEA0r0
uoaI+ofuiLYu4vTxub5Kva/pfDFYUHRtOHzhHtBslIJvUSemIKqD33KnnZDki1lm
Ys+PLddALNR52eclDJ6CK96sdRkyKPPY/JBlIec2N0PgpGCzicqXe/ev6gvKNG+e
I5RpoEWGLanFYXj1N6kWv+z78FhiMxztLUrA9jVzwOWmibxDC3htjp7jfLTbGyfH
qLLP+M9OfEuuDM71fNIlPldIi0DmJ6ud5NjpxVbQx7WS3BnbQN4BwA3w53NRDETM
umgWoFUEEmcHOMue1atCRniTcuHN7W2HSbZdK3bGu1oUEVBA88CbEqMAUVPcF6XN
5gJaqe2xbjgKTZ+vJPHrxPgNEAaeCdwx6x1yWu2nVVH/yaUWplIpCmsr53lN9zq8
ZCU57unz8Ba8ufklr91uYHbTTDt2M5y82ZEojKh0fKmP0TCLusg0eltTBObQ0uvF
giAmCml1XRK8N2X3ba8dnzHfgOzOjy6UwYBm0Syyoxe92WcKiiPJCtHpz2FWQ42c
sFMdX62NJEflXr4jGBTyjC1XiW8Gbhny5IEQ59ZJS7YczWbNVH1J/iGm3OZFWXIj
uo1wZfWlXBo8OatWnfujC3MFODWDHchmKASVM/S2AIU=
`protect END_PROTECTED
