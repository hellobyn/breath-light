`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxcANzqO3gNYIV/kN5ZJx6YuAsbg+muC98/eNXhvmjRy6lUnqGMPDylZbdAgs/rZ
KZkYxeH/BWVSteyc+iy41TOOZh6KRVly8Iy3s5910H+qGbBNQ512vnQqTn6qb7YD
ktUd7WKp+lxkPt66TxaZq7kq0tlk2QvOIqQ1omiWQKeC3KyLqScQoRjSJQm1F9Xp
bLGkSRpbkir1gkZOfwsmj/Mlq3zjwebuUP5bz/LCO9tufDIhhx6kCBwgmxFZ+uTj
mlWm10AgquzE1v6UK/fWn3Iqr327zaiIlGvzWLi4I40rzBhPqrmtFUMwhszG4+XF
dnqnU9YrPMRvZfCbMK0R4ex04x62kOTfJRHU4nE0Emqcv5p1ikh7zvxPAMo0oPVH
418AEow1ddd9zNJrdnMkxlaDUh2vqzuGxxMwSFYFUcQqchQA+rU8WO8C2FK4Nyn0
Sa3f5Wc2w7oxrzr+4sLWzE6RDTgoQ6rHTkds8IIhBxDuokhkGCqNfBktV9cuUT1Z
ud63DvqPYzgwX38gZqCI/I57UIVJG6tSrvs32jQ6lgGP/X1BUgQ6rQdml8Xb8DDp
YiiWEDJ6/s+h45YgisTtyjZdihXQ2fZ68drbpj5FF9HAWUtW1ZD5l8uDUsfcId9U
h4uPG9lvkVOythtf6iQNZ1A70E5DhitKPeA6rBQmIH44nnJMmFTdoIywT8Pd0C5X
Ezk36FuNx9JFLSorpCIv4sHFSshWqpvw03YHbedm8qFsJftlDwUwmUREpLiurYuZ
iZbzTDsz7XTpXK/oPbyHfH5UhuCSIdsZmSJisriwWlDjv0Tecj7Io9dB5Hyc9hIo
RwjdaCMG2aeJ+LYYCs9zLYgqSinQfg/Cu82FGOcyVNRURLBiuM7pZPXKhi2myuep
iNlqC4Gg9YjwJOyiLfiR7+hpX6zWz29EP3CkbwXjOimsJGC0ey8ndu+dNek4lpPq
g7gfbPhpiiyFR0EtNOZhK4RpsiqvRfMzsaoRcFzeoVPGFrouFN7KZDoyJQew5zka
qzaKBLHD/CDS68zzDULP05S+40CPjUUQU6R6vo59nw93z0XX0udlPrV60OZV0lnT
5/DShs2QE26DRccIty4GNHXbNppN3gPH3PQKoO81aWXQfT/qRO/POzz829gmK3fR
Fthw/RwHYfd8edUmM13mP8izX2I31EDlosu0cm3H1f03hWmrHNyiw6/8ifYjvID2
pozzq+qGdkSmnCy4IH54jGWvduKF18cUR4m4qImuuaRqNY9hogO7nxg+UoKwYiJc
aE19dJiArf/BjlEuW507Xu6TudPWu8XSGF5hYllPcdevnkpr5/7F5W42etS8nS94
`protect END_PROTECTED
