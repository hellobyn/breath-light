`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDyK3pd7RHwtaIICfOecbhDm9fs54/0ss8XQKobfuTQz1ekrrqYmAs80eAhUwNHQ
XE0KBhW30x1zwvhd4fRgZR8Alc+42xJXuC8NmznZpJBZ8EkYYEkz92540OKqgg8g
nZXwcf/vkdNxSt8Xa3VIQ3UWAGzHa9kUmX1mVi6xjx49OPgg04EPzXenoQ7pEYfq
bQ33MUVyPbsSSDTAC8g83n/ePitxKV84CbhBcn7x2SX9e7eb4IppRAh0c6tWynyJ
xodIwRBHpdBPTJY/Nya/So/x5dqnPM1Tbo4n/rjRNtTTfssE2lc4JE5rJ+Y4kJ3p
IwUgbs25xuE6pcVLnjUsnyxkQyI0ZycNBuzeAxG+wGcKpyGo/mCt5U3seXlfeFZH
aWzxUy9jqEhIQcAqaRm76eng1qFaK6/5DjVbg8tQnScpX1+u1J76r0O3I2seLitS
vwpEph3+KisDEhyMl1xuBFihLD08yWmvTdLVImrxxpG400q+ohZZ8GAkBYVAzxEs
3/jdRAGCm/5UWgyoB2YzmtbfRqLaYzkoLM9QQWFThQllzFH5c8HLiO5S9u6VpMDp
sjcSVicZjVL5/80SBZZvQqyqk37vB8GLn5PdFYU68JhQWQedZ2LMyVek1XXulgTo
TibZ/v0mY/OOODIlCogPAUpyZDiqgEs7ghaooHUEmRrYJPV03ddW87AgSBgyibN4
UrMrfpEWDZUFiQ919YLyM1UHPvgR2lqLXRPJh1IaFkeZt9EKOqzXOWmllfhi1Bfc
YZZ4JKBWK5lsDLV2Tzzh9MbGhHf0R2SV8Vofs6fmLxtAlZgV0xAayXXGkH5osbjo
Ot57tHCeBZShgPt9zDNq8wpQSvKghfM7a0uQb3Jgsbna3q69N75HYLQYQr0hkULm
MTe2GUyOzTrdvLUPUOe0Rq2I49YWwqtGmqGitYYJjrKxojwfSRqy8W96vlxcNlGN
2fe9DhNk4sPuk7nO3Y3W67pDP+bYc5FcT42wYDCXFhrf5UgUgsOX+HL9Pa28O37k
RIwHcSKFT+B9bSTcNmnISlegMx5/ocmW+6PGt7olwrupUKTzKcmkeVfnqhL7V/kg
R6Vts2cdx1ekqKH4S70IJcUfvm7y5gk5Etn2e/vRuvnnbdyKSF+cOXxxL+xY/nBE
kimaBKgCat2n095iXco2PLBeDkFAVt2FiXFZCGdDIAkGvyi/NU89/pzQYJ3p+4dM
LXpept9hH16a8rUJ14tkyylezFrwkrVEDT5M8IcqLNY7qDtv1S8UPN2XIVE0X9Ol
+dV7ylbYMGQM4m1sI766c1GuyDbKa8hi1nHAkLsN/VwyN3JR/yJbz1lHYSqRAJiE
YsaV9RS6yYTNlSUva+WKokZSMbXmOtA5XjnLrw+KytNa5J6eouBNFES0qVxun9ra
mdLDuHHC3/EeeyqZ9Y3ZPa4yitRbhYnD8xyxAoOY01Ck3fIE0SppXtMkxZIY7zWi
UbzX4i2/1lwBRf0V3J3o21FOVk/zdnVbUdVPzOeFEtuZEyaepCs7X5t5tjWSaAbU
jzoPiUoZnav3Pyi8FrjKelRQMlYIXSORmAortqHqXhzjBJWavEtjP/aaWtIRWMVr
7Scr4Vdfa3rr2qh9+L0LPoQTGNcOMPk8rB2pyiRmODDzpOohQK9zDjFZLm53EztT
Th+wlYvWBr2XMDujTm05cYjDVq/xShZFYupaN21oAak0ebdyaALKNfW18DHqD5Sx
QLrhsCtGJQ8X7lttJdzMtIn42xBHeQUB0B66D6u2vAvaXaeEbFCDxjPSNQtwMiYE
UcmDnLiA7H0WxmwcbiPAJ+HTMXHhzVDyQqSaCa+e15UpUgrlle/rd6Bm3nu3U18/
1yOor9dAkBZlOTxaoBdtVbCmafV1i6KX2VqUpXTgRlZz5/Ozs4OCnX1eWAbi6U2m
kZECb9txBfR1rYd5KWcMNFCpMx2nOaQPWGGtlc0CeFLiB8PbPoLc9w49NHfGX5uz
Mx5L+i84eSWxns6OJI3OdLEgcM9h5NaUl53nt91uevKF6i8YhU4fuU9zqUaomJIR
qkG5k+40gVlXz/pLJwLPLWUBMXBtp26YPpzcMFntK/j9SB+ZW3Y6WrW4Lcb0gIJp
1ibSl/dn+EHhNeVshZ9Y0O8jMWgNe0eKP2byBualGyn3pVJompCe7p+Q0dqDqGUk
L1VPfA0EcSN4YJCuIBgSCca+gKn40R+3ZmjgKqnqJSRGqyPJycDCxGU5gk/HURb5
jU9PnjbBEURBmt19vzy5gO8AcTqkCAKm2vufdp7P0elvRCXvuDR0ybtGdS5AMI6w
LBzqsSTSAjF4ra3Az2E3B4nTdCEq5kku6qSrOrlHAUswKPoQ3RSNerErTDzaQw9d
zwXsK/9E0lm3POBUEmleVlZxDG9p2XuIB0EfsC7z3AIHWdkYyv3/ztSBVJX1VSvD
ih+8m2E+tQlRwElaQP4ue5yaYDBgTGqsqau5a/AdZhUTETPoSX9Uz5ggaoi+oYFO
yHFpq4xGV7Q+2zaXnCXKficID+ZjXDiJ0YsUIWx15opJKOKIl10qPlL92JjbvJuC
np4G1Jkbj2XFKFJ9/Wm6Ij06Fzx5Fc7x0dRQhw/Uv3b2N3Bl5QFjruuvACbVANgD
KrT5nqY8cJuYRSgvlRR8aL/SvZH9tnvbX+bEw2vtY0iaTPZcFp+bBtqvfBfOYyAV
yGnpvqf/fFy07pKK/dQG8cCQiMzYMxH5J4Fx9ikyAuAPGm4yCSYm6l1fCxz0NTyT
6XRTGCpvvHzCsYiuZeZY7kCIiOGsuwxF2CKrAF3cV999U99XS7MKTZs2YgfU4zwE
hM0O4ojVCtAMNTUMhrNc6mSSq96Qlaua/KGhRdnCeKzAjl0+MGaIg0vpt55/KZxD
LXvzOrscaX5o90gAGu5JutvT7enBq+D/hlsGsS5fYCefc+xM5284mIXpBmH+kEy2
Aapfo4SRCV41wxFnsmccvqlmZMdhNih78tPnCqbQcqsjFPiJS5HadZTSKpA9N/ER
Fsqr0KAU9PXbHoM5uHbyCin/mbOGF4AtDKFpy3vBN/1gIlqV+G8tqZAziS+fNGtU
NzA39MV7Zma5zWLxJaHYrbzWktbY6aYqozvd0zzs+Zl5RJi1GNpG5dgF4exeV6SZ
4wTIE4yvSHUWMVCb2cFCT91Eldt/x+LAcmxSAOgLVX7pZ5dRNAI0y+IBjBMHy4Ys
Qqz5m6VOgxQM3xcEvZ9/JMzkv9lV8Nd2z25uCetqbEx0Vbr7DsFvdKIOrpRswmFu
hVDp8Tbpjn4INiGx8ZgptiFp6fJSNhbKtXXAlOcEsIRjr+LAmHYLU4EK7vxx0teE
KPtr2MFamvrEz2xgA5Ahkqs5OAVWvCMFLbUth7Nr6GPAhKjzmnyTOw7Qr/tOFzmI
y+B3YkPaG83K57WQSjiNKQaVf4pgQA2Ggr6VSIGqlB2XcAt1pD8ohSR8t2GlWp8b
8xfuANFsQcUJbmqUCSBdfdemIwagG4/MsE6NuJbUGABTZmo+Ywz68WB5dDbEr7MG
rQqSQBunFxhKuAZqD/03fhGyuWcfq9kmWsiX09dxiq+XTu9ij0DPNUJE2DtV1+Bp
Yhh7pNXAJAUSuw40V0X1xAp+IEszzMcxV+R6XoSsyDeHqVSRivlW5S0ORL/pUj+Q
gcnsLgMZQWH6ftA4vl2J5MoX5HTxwO/3Bmcgdhckx5rVqxwTAOThr1LgtrsuU3cM
+UNQGnHS5ciWnavUeCaMZ5RAh3tPbYxvPNK4QpxUeb6E1pbXlHZ2UP27xqgy76Jl
IxTPMq3teuXqw5yWP3hITTX8PEZ2d+uuJs/yjJeK2aE/KY+W8x4HMx7+0FSZC5HF
fUOMc3YHqqRnUbzigw6i9eNzUofatJ9PDaSqDCxIgfl5bXbohlOjqlHJuQlGUwPv
DmNBZhkwjf6LNI0iTuh8x2+1s12B25CUWb/Bl97im5JDq9xon3OSn9SVdSsNywQ4
ZP/aGEYYwRGbwgpAZMlsxpqI7g3pgv7/gejuFgehH6eNlRUV1f+q6dVLSVTdavW1
V+Ztxo6b+kVr+dpY7fD5vREf0A/ySOum6BgOAamPRdDsmcMiqVryavJSXsu9WFF7
bjX4ZKDpWNzqokhXLegQhMSfIIdoYSPKZS+6U0D3j5OSgGgmlKIkYtlQmqIgU4Kb
zfccyk+fOr9UXdtY55FuP61FPdgAectx8SXKOAEDMr62wlyvWJJ7JQ1b2iOStQZk
bqzccxnXuWdoMqrz4ZB0sjLhZNBde/Rn7a2wH3Q7A6oCZfE8nfcxvDLd4jjegZCN
UwyXiyvoAOQpus2R9V4UoqfKUZoyIFg4EqPlOLtAZsj+beab/cGKX1CiTMRBt4GT
4vfbsP5ZljCkQfWa2E5uzDiOGzFvxCGBzK4Jgp2u2JFX524YB9TKsIiFvgY2PQfM
+I0xyy7a7ttKh059qa8enBVNpxsdGy1xFw69WruTggcTAQpgnByQRmBYVLSgdnkz
iyvvqz1Vt7zxDhmxrLkyP3d4aiMoZBYsYAu6XmxJ2hVlYFX+UKdfPu+iAWsAAzZ1
BQKnJHSX8G2UoE1F3Jx//5PGu1Skhyrs/i747YogsxQstk6/s4PryEYa9sRODqqa
AY9u+hnNHj93cWf7A/NszXCFH+Ex/Vdt43L8aqPN9uwVJAqfcENm+KB6UG0FieG3
A2J3bjiMnIck8dqxEuDFZLz+sc9v7s0F7u5d/ibduBJAkAKuel/tyqV4vYFxzRns
0L0pQlIxWXozS0VyH9CRv0RAmxUd0CJ1kXYPmca2R0edTE8zzqOtvbLLYFc4BTvd
1C+6rEOIXqSE5klOT5jUjcxr70OOcLfNELJsibB3/HpMCJ9moJEaIMtqrx6940UB
8/7zoYgSeX3my8g7Wm5Nl0MM+jpcL7qe8kE7FBhwWd+1+efwg41Xmxn5vqBoGvTX
v+URwncYRkrw3JbN2uuacs4XNHxB28PCDb+nAZ8MZXNsl+XviIACsIFUVdUyGR+V
Wu/AI1/EYNEyyR7Vv849AO7OqMTLjcU5DG3ZqF1fDTatfl4JQJBmj1yZieJH7vzk
ltKgIo8Wy8S/KXk7Wxul7UB1Iik4FlE0Garkdx9v1BhSJGsyj084K0rZ+kbW42ZB
qFh9wKLycZMq/60xR8emt/fDjLVTSMKAoipFmRLaMYcmpOcz4rThyyShmXhO4P22
ZkG0OaJtwX3EgnigZwKbKsV8Ee7L7s9d6DFf2T79L3c1aCC5AvE5a1prNgAdtk9m
agK3xBso6j00fo1mtWf7QOOKV9E5MCJET8Ie5T9UqQsb8yfsffGQyB5p1b1MHJMc
osp784DtPIZZbcPIQ8oUvUx40APmM4gggqyQ8vayQusSRZ6WZatSKJ61cnR7eSdV
/eKXewgdrZ3MdGhsmLl/7YD8sUCeJXVvrg/1oujRuAb7sgyuWGZY8bkT6igEVcEM
8G5SdDevA2g34ob5+Hl3XXnBCUpJ5vcFoAIShQz2QY+r5seBlLcI+aIH+xgAqloT
1Bqp5FTqJGwqtz8YPZXaq7bludPnGfuOZ+9N+OujteELoGxJ8n5W/21ZzDk6vh8G
appZhAuD5zJsT0FKrKdsLGE2kNna0qbuNyUNTbV+QFw5SD6Y4twUfdM3StL+FIQN
lqbIkZTJgHUFYB8C/AfhGeeZhdfPdvC2fMwxoG/d6S5hhci0+4c8+h4iDaP0Jbc3
6iXd5L2wvUH9OlCEXR6pGgtZT+OUFFgCjKkxBu50/9Y0b0VC2SSSQMIbdc1LPEnC
mrtbs8T/BQOj7oYG36cL5mnzrUxOqjfdxeYfGLKafTadRPBPABdYQZZeBX9H/cwp
XFNS1ck8d71qsLeEVQrA+SR/RbuwSF+Z5qsDZoepbk+q7wtYEghfBMUysqGa333U
infqMem1ZrJkRZQIgFodAAcs9khhA4h8vTW5OXxZ1zhxmkk93jIYD5odilx19pDL
nkjxVpdajQvZcgrSEibUZde4Jfv2Yx64dhRRyTiZCTX38EoM13f4qh8ICr7+dex0
JadYPGqX2SYLvnPQMjxmn2stjivEbVs6Yr/fLEwPxXmherM2QgnMzxbrxYenz87Z
MZAUbnJa2WsH1eb3CifQ8Jtw3LUCfVYGXtf4HoMvvoTRtN8tffwCOx2Kf+Ine3a4
/lkUMTnzzZ7cnDCBTXZv1qyQNBvRd9Nwad6sx92UhLC29T/K2mZJEwKju+s1kADT
unXyfKQCtPGTyUnur0ih5pMcsZkdUbdGvpYEoNGCEZHFgz6fonDhSkjX0pc4YFS+
ssNaTppx3vljhxXlPqlpKWEnvhE2JTwMdxAoVRlLQDZKmqMww1RZ2pcmp7u9zeaw
kTwWuMqVl5GQbBOTfmw5c2QuZaDMYS0yiaWY4S+O3wLly9k0cBLUUI8SmKX5li6j
oGTOakQ+YHJV/CDm5Fze33YmoFQXG+FTcNd5RufgQUygsCU2Zp10o0ayqpw904Js
kAFpNacvnCu7Efjjv3HQWS2VmOq1mfmNkdXzpUX/TyQgYP1ZkDNTFFxjv2cfCgb9
VXz+g0pxXcd4dGZmhGHku1wD/OhdK7DI7gcxDrbcH/RkFwTV1mhoODFfdaklPvG6
ddOnB/2blB5OQOolSChfyWQi59mP8QfvEpQHYtS5sAx6elsf7EyrZoxzQha7Jb6b
xEieHLrcDW+Os+OLfrEwZfK2mBVqmycUwMloj4Wt+XSuQ0Ii341sW8zLinT7CwE1
idOZF19ecNlsjwmjJMKm6+2KWpNU8KmSbdd7LdzEZ961YsadZjNIh61IhlbwYoRh
CClaA8Xt4Ulz+bdUHHxirjpduXoeiYpmOVWHTstUfdIcw82/pfw743LNsaHvd0Gz
629n7wJo7wbIT7TgU6/iAMaak8JYTBrcDR0+s/JHsweWEPG3UN0Q/JCLdh1ldHM4
RvS+Y1hAlG3U+45DceF4lM5eyxI8UXxROSaSN7FkryMlci4X8+EZh3abYYQJdwmb
EArspzA8yhm8WW2u1SOfJO14Dpg5yioPs72p4SscT448UcyzpBghyaXlq8CZsi3a
ldt61cjsyCABz7myE1nJCWGeYktYpNrj2hpQUU1jnfBNst1sHNLvBM/OhhCyNd4r
11fG3RoBZufJMEfUzthvHruf9F/2i7ydRorJdJcwfmxIbYkefnrhgvnBke40xyAs
NxMFx/Gg+I9OUut9104T1Irbqiy0fJytNtRUrB7zOKl6pH8UdaQBkmy0JBAcKwnh
tuwR5vH5mQATYPIss0K/1vGkS12jk6oxNQX2F+qY6A/ZWPMErZFCql3KNQ3WBrMJ
SMD+OgWfL/fVVs9BdNm3qOe8fNVWaopCKPQiEjMFY4gEoZh2o54Y7AcVI/WtpG1D
itf8GaTrcWMeRQs/ADVIloWxywey7+sdAzC7t+swixbogyw3oZQN6zDaM2Fxl73h
DIyuG29ctUIH7b4F0+yb66WVPsNwSJ1VTitz8oVSYMe0Mp0JQeKkbJLSIPJbTjgg
Nfs0qA2ZcXRYmESx1XowmJT7NMymTVhy7+ZmTuUL7+FvCm9nTgSIxLATK6b/C3yw
Zan/KSxa5w9DFATqfhXNWFSvSgSKNri+NdKM9Nn65xDHjJ+jr0JS4VCCRXw4YtPO
LrqdIu+EfTQusxoCINuAwj8ek+P6SCbNDWIcy21Urx0qK07BZOoNFdi6PJli/mRI
ESAIViViiMA13ZYwlNmmRXvW/4sfbyXSwZEdp3yjB2KWXkUAGNVmwF+drb1A4m9h
dtcWbXDz9nLLfD3OPwGlc9sRv6/ACC643Afxw8nxSXPoh68eKKZVsOttKvofw5f9
aXQK3zW5i1cI0iSZdwN+h0jQFK2ijl1XbHhZvzMxIrN5TX08oIHScxVaVzw9ec9D
+PlK/vU4IncdE4Csxo7jN7fXEd/ED+bMFYGXuWD5qroS1hAaoIC7NKXQ+2LNNQAj
GhtZ4XCdX2T/Ypnc9jgxM5ha+6Xmw+tknuGtWHGSK2yplf+wX1v6bNI+T5WqDpO3
qy0UyTXAaAINztc5NjgZqIwecGNAUIgG+tV4Dc6cSz9NQNqmuSvSh/lPwFu8BayU
cXcVry0tzwwXuuV8NKgYfWLo2Wo34fQQsTouzNGECSo4YjwGzcMeewugOfDHZevb
1511uyP7L0OXuIbS7xyqs9/HPTT4NH4zGVasyjsvYtFrTQfq3VqBkSE/MMatE/nX
ZZNG3L5VIKVu5sByyTq8ZKwAgqWhhXtQGMUPfeYuF5cH8vpDE5iukGfZHQ3OkIcP
8uk4re4on9oFaA/nOhnPL/dlDf7RxpOcs4tnu5VHm7WHnE0SlSWNnbc3JDxMXl8+
3Lao4JNcOBLtHGX2LGfAtt813QMAa3ntMfMTO3CwYKe/K5GEHluUNPTdB0Td5zp7
joSUumfI2RlfJpcgk6IL3/ZdTP4STXFm99xUChEVIvWMU4R2FauGhaEU/PrKJ5Vo
RbdLpYJHFw/kyKhaYca5T+Pa/15kcz4KHi0i3wj+skalwgV5bAFxIo2PIra5DIPC
/taHdj76/KjJVNe42G4NzJfRGGgNlOgvqw12w6us53pcX/d9ZIvh4G9+i4o/1IUy
0CF8wM3MSfZPoFAYlTnTtHocGVrEgR9mMrCHWAAef0S9xOXEMSeQDwljGQrdwU/3
IS4gGxjWqxFtA0rvB2+xHVwpmGBQhtiEDRrWCqe+LUIdbamIa4Mb86/pnUPkxD8Q
a+XAaxWCfXH64H1hcPH5Hc0OCLBSiwRECg3Y9R8SS9QAqPyhIwDO8JRV1WQY/Y4F
uW68JlL6Yaxzl2dpKBn9g3GfYohh/RijAiSz6A+ASewolz/PstjK/uHfp/N+Ir16
6xxPoEjS5uBla0YB1IlZt2IgMBTC7vhzD/HQ+4ltwNflns0RAFcsL/aOnftUCXwD
fj4ABjokom6PnyLpyZlcPSC2FUmwU/J0/BFgHkYeaz+Zf4i1GVi7qRf8xGaP19ME
lhRUOxr2Aqd2jcE0BuK2h5XzJT1zPVFuOECXeLQzTW1XynCJMCTzPBQIofuDZvvI
u9w93VV0q/wV2Lr9FmUC5eHf7Dq8EheQrhUFl4TqQRwFQqVkJmaLKBSa04qxgViR
mYes4HsU4ZlBLuYTTuyf4TEZbRGlnmEhwfsWktRfYLrm2J9g7Ewr7P4fIQ7NS75K
RL9ZGtPLa/5ySWqDrihBJ/2wOfA9LClxKRAtCaehCPqS5eQnkWIp7QkNer4MGRiv
niJMdNnrZk9ZGukeeobZ2B87SsOs+6BXekUbqvIL8on4NwfQqZ6YPSjv6B0l7QlA
ZUN45WbDkPO2nPXgYFeEN7YKxEwfljzPeRZekqr/j1K+OVQqD5FAkNRgS/rnaXku
yQVbZHN+Wq0CX4ERE8D118fAQ7cH1EjivQTnEdUBQOdht7MG460aml+5o6mA24o/
ncrwpOBL5+UOygMyN6zHiNH80h03+bGbS+tv0JtPpfrzFu3GqaUK5grvrDohjdas
alpOZMg8ue5UUlMXU4VDrUs9iKMCFgSqCf4NiSWqKrV/JR9eJCrDWUHmqkV66DO2
fj24KrO8j4ST82iPlKU+fG9t3W2Pyh2hVFwPyId6AFk2C4mJoSFnkgLpn9OTaJ6Y
Nw+spBsFB9GRrhsHNneNVRnoej7VpzCbZ/n/s5nXpnpIvCDNgXXIBskymYYxXm7j
ENGbS2R9QueiRF6SNUZjCRP7N2dhZRVa1rkPZwiLIMoyjRlDVW7/coMTfl1MGEmf
upvtTxxrtTCijjb0EncfshL25E30wOWmSzT7sBC6HoMo3ZHMseDwg3NqQgfKiB0c
+CMiV1lLKfSb0RDESyuheGD/UMur2x0uiLN1GSWUAdivO46l4LcApGqdNgYSM6Y5
GohNqPoHKw7iHSOKiy0rnolpgr3h2tVssmoTykUvswRlqzq33vHyh1xIzGqn+/dc
6X7g1hidJTJ/Pp+d50VDgn+TD1jMvkGHjzsGp9to/cCQBewjUVXIecafO8tTbK/a
w7mjYszwNkgYEamy29iUwcwwzRJHYoOVo1O/llwRwsvxETnIGTyimNoWqsOXrOOl
QgiGUNagdw7MtNcmAzcyOJi3jh9U93rOMQaCc2DMj66Ve+EiSUp2jdcu8tWTqHsS
aRnLhrhhmu5F0fpXuEmiFYWC9fVgt+h2G92TRj8NnpuTnlMElHK5W6TxY3Gkd4AJ
Mk4S8snSQVkJcqV2Bg1NtOiQEEWXC8O709iv8tvHnLlZ9ipxZov7TXVb3o+MaQDG
znxwKFYngj07W+DucHm3821xLojVZ7hXScFsj2EcbEx13mN5kEgsCy8wMH6QCggw
MHD21JSh5c6goiLIa4mRNCrn7k/VCSDVBoKB2Sr2cMh5v9nKi93Z/rBhCJl9bX12
OnN4ZC2zEGsBGUyvjx2TPTqq7fBjGG8ijEE6qktOxOI98eRd0cS/R+GkGPtOrcX7
R1G6mkNtYfWvsW1mP8Qz6k4ixsq/k3o8EY46YlbeeGJkaK3lDAPGEFhSv9nT8m3E
Wc96Ue9YGiQ0yzmjNjhJhywOW3M7XonHWyLavbg3u9QqnxNR0IWh//83dIB+7hjh
LUOfAE72+cv9cumMmOD8yR/GwOonZYRKehxlB1gJ85AKCLLHzCmUj7DpH8pi4dhx
s4fdy1WKkJFmC6++3sutWOWVQmgfY4aGJpff84cYYHkjqp4uLD+/CUGRrCyRJG7F
TKUUSOXrzfE/TbzPk5pJ/kmoW8d8njCWLUE99PkQwKKuOcuVMOZKeUTlG6WNOeoi
6yvEtXXc77pZBv0gX5WbsY4DNsEOcx2vkP3Aa4tb94nd+eSvcaYriOAZm8bumb7f
xYHJDLd/9aZ45PHVHeHNFfJ8bMSWIwro8tP5RjGfFpDNTI1DDQ09JNU3FwRsXRK7
3T9N66qoU+dcAN4CN09LZYbEWB5f5FYSpGLN8L/jOxzSVe+7+inYuw02nCSatclN
Sr0vjWs/uxSvbJ6F71cTx4fV2KoYtnt+r8N6j17qNdYzHDmRSKUa1zxQoHDKub+H
qnVmCsysMLitJoxQ5Ws8mtHrilUNVRqmDpC5CYbIV51/w81UeDMxnbDdrIUWVEcS
rT4hWJsqO7e8AtgnHXFgupfXsr2G/zMPxXH7YGaGhT7oSULspHVjExb8JA0Ecn18
tjrcbKIwSPsqSdg3jYd9nDUxaSABsFnjDfTs0v8m4zeNIIdL3I2P3CSX7NlSWmAP
8zT8FcYfcSK10KuWU1kSN9Veai9MV5ESLsh2TZSrhfS9GuJaBaQF8Io5QtKTKvXR
Qqvp/qHgQl08kb+JzhNwhsnyVL9AR/tNtu9qy0SOZI6ePKvAoaMrGuuQzBRRMRBX
aYJWbGdDfU21eYNZcLLcO663gHVlB3plBV9KTBD2/gzXeqdcasKZ1rEVezknoGTr
wND7Jzd/Sxvk2NOiDlXBx1UIm+rgw57l+hh9cMN0942+dA/TyQtIfHRPWeSN3fuf
xVasep0vSNgAGjXgiGyOhWDNjlhUq/rwmfqBVYGw4LCuEGdyEASCHTOyNl7cklJ9
Rak2ys0W/k5R3jXjtx50/Gm8O3qqer1CRJk1bIXAV3019hoZk93tkky0rjJqNwvt
0hv5S5xp38QN23LHeATZp3scpw8tZpfhoJPV+1jlJwYxLdmmurb1l/3e/MX8r0kC
K8hDPX/Mz6h3n+sQb1BBTYISJ1DHRkRDAQJx0RhIOKYE9UOdyo8SNcKVuM3HXxkD
aJ5kd8eVxv4x6KIZ1uKK3A7KIjLlSwFkRsV3bfpO/TgIYE5kI3L0PsZZmb6ed68v
gCPHbYbaI2NVsfUjyEmWh0yC/sdCjK6iIthuiXk6O7Uk2qqMQ8An3UybJzXqmj38
pDEPisvQGnsz7kIfvN4r4er3MGkkGSc0zpxBxQ549l1UNheHRg+gI2bsgH374Z0D
QMKtM4X5EN4gfmMce4rYfdgULILtX9Bt2+7J0uJWiW8jg/a/EYMvPpMOnUr+rxjk
DrJH0lShM8CykbLhx1c4eAMQrz2cQE8BnY3Z8JvpsE3hZar6cehXE4pks8UcJw9A
S5xbYEZeE0vVfIRNZrcKNX2A8BrrySUKbUfbG6JwaUDyZB/tUnEJ/oELDpEnuEtM
Ufx9cr3mzOCQyq2Hk28CA/SE6L5BtsrUKC+f/ElF/TTyzjKQ0caksRHwHgPXoSFy
KAjI9pHuVpV18kTcc24/B8tlrWHG83Lj47fe0WvlODof6kd9SrdJo3QjPnZKGYqG
oNBxs0G6zLV+Cql7QUCp4zfhFeXFJHmjK0ruCkMvgSvgbRGTcqYfWP99wgUV3Ac5
JiKMcpFYdon2Okc8Qq7frwPeAiaIVlC44rwQaSmlscP5xI4kHrEQamzZkVcAaHd8
TQ+w/Y0yojVm+TRysKMZmL3fqNm5eeK6crClHzKkUjMVTfPlOCHQsTbouB7D7Yq3
ZEkKCifp1S6b8O+5dgHo0pK1VzCgTUl/JzdU0IygpgxwqWSP5oaUxxLZpR3MX+FV
r1/mx36Az/rTBcIYmtziRDnwPNeCmIYy7YkAb3nZMBwE4nGg1rK+xB4WQxsSvtez
JoGLyZ8NdgftHUTstZJAwv/38aKOqgfxLx/MfpFy2lPT0a951/wJWcda6wCvloSA
IFLu9yYrZNaVBgyc7hDdc5MAAiwGtFUnR3jr6C/WomAlCMPuWCTFc11QWWuRA4Lq
7PcpjceegW+jq0qAK+z/mD0eTlESdUUAJ1Al4UdnxWnyo8PeGm1o6BGOv3shxT6j
xClwg4uKDb1pfYV2FjXH6kFExvx+RIUKCs7x1oXW7uSRCUF6RSGz/3qH8vHqiNdk
N+uYEzLMNuQhhTd9Zwra3XWEB7+PneXemdII74HhgKVQpwmfdQSiKKP+dHUqMzwF
5QiCbNUTgFYVuzEGUCSNIc4a7xXRlqjwpmIvwdPhk7iJqlTGKgmTgf6l1FeXCqKW
`protect END_PROTECTED
