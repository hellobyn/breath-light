`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7KgAo42wq5CexqVaOwM0I+NwcrZoy62Ef4HsmpI2N+bCK6TKOeDgLDqo6+X5ie4
l05XQukpxfmB1C9ayih/YEFa0zWuUvKLxecsx2HCvVqicrUxvXRnhYSDiv7wxAPI
RpuH2tHg6DLewRWwsnzIhf4TlEJ46ZPUnd/2SyRwqXg/NEV4zQtl/83iUu8xbdS3
k+B4ydUebTMOVXgHOkoLVdQTnrVQfMLXj+V9ZTFH4O6bRuGpE3ANXgSs93PE350w
2LnTv4CvZFrmOcSakeUVGQn2UFDypCEhNtPQ25QcxaVq7XKCx9kUDfvKHtU4zLiS
+SzOOA2EXZr3C+aG315qH615zGGX3ZQOcpZr8pql3KQuSlJ1zl5L4QhnTWquQ8Zz
b7M9DS09YVLATE9GcrBGyecW9YXi3Iyo8d3wqhfBna+jhk2rlk+dpMj4p0YtQVzq
MPB2Z3Jhq8qQ3U4FvRCZ1c4EgtwfPPAB+DAXXJLppX88I2Rw1oia9JXTroTQK8BS
JcjyllSae9XW3FosCEb7fOubFaUfOVRnDSItEI7hAXE9Q7Y1j7HR+7mjydQ1jxir
1ry0FjaSF3bvzYQ5RNBb3+8zWGrta9aLq3TV88rnXvk8V5X0kMen75NNjIOLO3LH
AGrTaOfLAffMQnnAAzJB9xQIa2YVJ5aboqt4K9dNgGPQLXgQ+ZJQJYdWbu1x3gXx
UyAL1b4djRNL3xP7/Fwb3fcg75g/WdEjzj3wRajh88iA9Ocp/whF684ss/ucgIRD
0lEJN5rAIbm+9NPs/Twq/tR2lGa9dUHefq6F+GOXZK6tPH9fNKw6K5AwcjS34FTu
mBM5FtkBWfzyy1nVKbyo7Gap2IBTyN0Zs6KDTqewbJ8uBPPTbp21EKvhWxsO3bbs
aE1nVO/qQTfy/pRNexD51sq+139g9ilZuO9/wOiWqmg0+PNGq8QFXhKl97Ro7Z0R
3wWhUfnZ7FeD+/KTZsQdgRF50abtcT1IOp8Lzb5K14289WNSAGh6VGzm37LjeKYy
w1r9xlfAq5Gg6TVPKh8JF4U9ViqwNvn9+SFrb81zEY7bghLlkxOAB7aDkGMGKf/X
36aPAt2aCUl0Ox3I9kV9Olxqygolib3sGdV56GCqNpFCakYrp2TEOBlcapWOkJOQ
oo2vDuLx1/j6IvxrlyOxObbc2YIM71uNHGoFYMqvHinYrrmBWCAuqmpZeM/2HEnH
G2rop1HzU8daFX+AlZztFv6R+1Y3F40zaoBZUVnYlli/4ft+hM5iMOFMr7CqjgLT
CsQIDR2sfaXiofZM4Sw2EROi8WMOb+w2uCwZa5NRa/hG6UIWTYhkJWNquV4CrVnw
YSZxUDL3WEpZOZ0P0uv1T8ITEtQwkuVZZjnD321K9ULnp4o72oyTX24wJ+AtrKAb
8rPO0JbCHTv9u6+Q+/8MuuSPUV7457BfMo1G9IJajl16vTTKNJ35hBUtUsZwKKll
4oIZxe04USD5RP7Jgd0BUVigjzwIfOc2JGWL0nA5yzg5WW+DqdetV7EvEVWBfshZ
M2BBu8n3qtq2S5exH7tuHRNlucOYAfuq61Yr0Qy1gmLn0NPdeDYaBdp96E8pnU5a
9N0OCFxSzXaGrTnK+Gx5aRKAItUHSkdtXZjRZukhlSdXkvF7MuvuqyoOxRcTqEZm
73SkFsowGj+hQC64cfbW0+GmvlGeIAvKkjrZuG+VmOuvnM8UrIJZ2yU4Gc2ou3UN
OSqTjfTSJmV5ndBlcFwUQ5qvd9M0T/GLVwv5/hyo+8T4ePv7EezKlApD0V/5mD/c
XkBteAsAlZMuWKVE97HvPtUlxU2CBh9bqEkwkgWe3PGKYATn742z6iIrLAeuH75s
ZaXowsp4sP9vZna96dUNv5gX+TIVCsN0zI1ZqqJOb/0+R8OSZ/vKKeCuVLMPAqKv
N8UqWD9PM7qNevv0dntbFp1qFI5Gpu8c+V25n9WrqwFAM6Kt5KTjz2/J/v+slFoM
`protect END_PROTECTED
