`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wEUcJw3YqrB+9j+ctKoeRfITaggbQMd2ZzkZH87a8SJtEUgBv1r8Zhs99tYCauNC
h9UZK+zDbJMaUpjAiFmynfuo3ZVaQW3c9HXlrFCRFVggIJ4+B7NtWBGy8/Y0X/mK
k/jpNuGIOT6sk+f5y7J9yi2UKg/U+Is1krZlUVg+bKniAYIG0QV1VND6o85aXHsJ
KhPsxwSaZXlXZeTdml5ylYATmbOupC9M8WwjVzR2Sm71MZtR0jw5AVN7OGQ0r58N
00LSAtfASZ5ZVVKvKcEJ5TlWIbGfPz4RxAh5ZUr9EoZivYaS0RptcSvgL3f1VqQ+
nessAvV59f5wu9BWsrOM/2QfbCwO0jeELwBS1Se5R9N/pHBAfhsAxKDFSGbtU15C
atbRsS17lGZra0nW+ZDWvCw8qgtApiAoz7uWn50HbC5G/8isChwMk9vFHkhJlELj
eL8IQbi8tNIkS6LVrVPyMpKeuuhluEovPsWK8S7XoC2SSW9MBYeBeM2CQL0d0CjP
5ixA4qSeRlHJ/egGtdPfDGlfVvxi9gHl2pOBedjNSgdmwiTM24OGXL83DUwiIaUo
DyXWqyO2cpgzrXlq6N0+j6iBEEhk47ZsPZDArMNtAeiqFrH+aAfhaQN6LMXh+I+q
RebsufY3WeZZvr4upyTMp9mSLYLaesUP3mkjMgZ56PzbBxy8YLwc+41+llFQ61I2
OtKgXj3viNkkXy2rZJP29r6+mCcLJ6aYEcGJt76bkpWU2GwIJ5Nbe2L8PYcEDf6n
jhJmx/d9VCP8NtI3JKnGwBR7P9tFp82DRGt794Q78FtLL+L2lIdsPIk3gEsZLpB+
18TEuPZAzZZptclRKva2CSukCKeySPoS5FFFpMHvCotOB5niI0QRWgqcuo4IzWHr
qWFcwhp69RCmL2hl9VrtPYXOLoTV/BJ6MTSDRHxB2Cgnm2DGzOeWqy9MOKuKcmmh
mmJ7IcKWWfFb5ugpSFXQcaEUshg1ieJ/QiQLccrOqbJ9GMuKck3pmflmFIyE+1G0
essMgqLK8OICcJX+hOqnCpApspgVYHMAx/rkfclTr2QWwEMmxPoKih5zjCUtKRs0
AUYDuZn9pJd9FqLF+0Eky7sU7ycFB0FClM30JyXYNJYbodeHvPFbXoTM5r3qwdSB
MVpmnPLJZfIT37FULeY0j/YL7i4Y/IVNB2RX2215f6yD+sL7OqzCFDp3XoCh9BD/
HbafK9z45QC9Sjg7Yd4k71V4PJRhAYfLK2dh7KBQuudtNcC6mLpgXzVsTkm0jXf9
OfAvJpkZJA+FsLkDhb1giI3eD8V8lKEODHRK/xR28EHFgTVHzeMUXz4ZGCkOWbSc
B71GteV2R+xRvkgxjQb8OA==
`protect END_PROTECTED
