`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nM/esBVcdue4cwUlZowvaopEZ74MViqGbJoJ2WnVUnYspEWKurwyT4LlWAixEb+p
chzHFrCox4wLljq9VORAAuaczuLX7IM0KDaJWQwTwjC1pPiV0dUSYxr0Ky6udu7K
IJ/KwOPoGYahlSOtnw1VUD058vbDaomNC5xw+5AJ6UTtERzPqx5Tc5lkpvpPRuPh
IRBm4F+fizhSQZT/4fBEjOW3v6zs30hB8mDkI608Hjuu4xKLl9eSMAUY/yxo/DJP
1BEk8IuLmTm7HAsUX7pECbuEeLHT3y6AQVVgI0DuGxYdjmLE/0nihFyLqgiZaI1O
+z69KH4197W7TEZR7Pd6QarAonrSs7JMxGysFOyDYZyBx225Y8gP9Eqq/THckw35
KeynaRrT1do8yxqvYUMl4HNCjJorDJpzSURumC0msabY0CgIOA6wq/vemfbGoMKD
WFyv9PIW7jOV1y9ncAsbnQxgfLEkLo/PgLqqbphxVEOmQmqzDN030P0PyatOcTXX
9QSfbbJuj8Qf1MKvmwgJJS2f6UYFUiB/uZFMY9fElNTit66RfXc3zPjMlYf6HKVe
EA1Cc0vI5G7A92i8cpp5CSHQFlz/y/cnWFX9IyBu8FuKhryh4mxwLJMAznnyPfCY
YNcClQnpZBakt/8ogR/ICR5RuMMjOJZ/W0VYGDHELRCgtXUgMxeygta8zg6qWWDh
qimr4O0BsGhXlJUm55/kTV5mwNKZ+pqncvqYta4SUhdKUI9duCa5IEChRykrC1UH
3NVQdQGrn4Kur2yrSFRjtwcWM3iGVNvOF4xkqfbusRoF7kPxwA3lEnThQ9G8jBr5
UlGas7dvYXsIvoMgqq6Au5l5EQeRqcs6WC9TEMEQVJv0SnzJWMgu8NNj461qxZIG
4pNvtF1GKoIJ7wnkwuuD3Dv8PcaYwS45HSn6+iG82fwtQGYLPs84tPrlavBfr5Wp
Ng6p+o+yq7PW2JSM5ecVwolqvXidP2JrRhO9ERNafFUWUcWx2yHkKJYkrJq2azCW
kytM7yh8CcqBwa4V6NsJBo7HWz7pfKw7PU/JC9EjEKUBxWr59RY+DN+oE3sfzx30
f/SWL45Ov7hbJaujokE8TEi5PReDX7a5YvUC4tXcCqfNo3ZIl0QQXfy4upc3eyss
IV3RQS+nykKXcXHJmVstpHbDGlxW0DdD421WM3Uh5UklU3RfRXK8+roLhe/vLVYT
Y33yQ3ylBl9bf/gDKGWyIEw50N9oiOZPIxDbt8OnQVBJf+7pD1awpiKyjOWciaCA
CAgddLAS4tANh4C7tsmdQZyiraQ95yrenRkaCYE5mxiDaUbpJTBOvy+T/T1Tp1PS
Sfsd3UAI6+s/R41C7F8n4OsxG9EL01eBsjIHNWZU2nQWLjFOVHbIZVcHzw0Nei64
6BGT192WUTQklHGCgHYgCLrBzJkKHMnhmtMfCr/AY1/MyK/jo1jVfPEDuYe6nbe/
xAc/AD849XLHDHve8gdeJsEvO/eUEurpoaNt3CAMPf7roBfSVzTWIjeUBZcZvreD
giuXbJq1q5W7i1xuSxjBPulWH2inUl7EqE8H1AcK7BMR2ey6vfBnnu+gqPIegRAo
Y018MM93FzLJL4vC93YU7m/buUdlRRbZXNYzsmMhxUTLK9hS8fH5V47WwHTBJ1kf
qJty7ZQyoFQCMnQ/+KxbvRa9mVUF/XX///lrhb/uOzx4890Cn7AK/VPJjk4zkBbd
SXun+M6Wb36WKQZ//J9BJJzh61mzfR9/Vrbsi1+3A0D/b5+2056N+uWoclt1GnuI
LwVv6Yujmk7IuvnAgBgmaAeDh4njk6VGA27xmhl5D6LOsCQ2OOLieUe+HYYwLFCd
BjdRTgFuyN1OvXcJiRS2pjl7uvnronlgJEjt8jK4y2BID38gkXrIX/YcuNwf/a21
zkUX7kYd6lB8+t0/QP8S3GOZxAXh07tJ7RdC/J4NlTpDGFpaZ2l1r+Fbe7u41Ow2
Wu/SR796C2nvGkpY0G7UU3lA+Lt3BzRG4Q8INle4Un/ymT2h3CYLYSos9hZIMLFs
jpvwiNtiAgbI1pCjklrBk96RppuSPKBthGdewEzDmTLo2UWaetz2IdpnifiUJYCR
Ghzwf6MYyI5aUA/s14bLZUyq4oycoRgzUB8S2FsyN+TAHFsirPatIGm47CCkFChz
2Hxd1r7p2MumYedYD+lNpf6AZW8ull+38sRF4d/lP+FSieV9B1arfIaM9rQextlL
4NrQeKendmnNlan09gAJGnivUaoavaqZZNoGOikmFUFpOIHY/1XY+HkWJeKQplL9
3ctEG76hVIbTp9ldHHXnTMlqAV3SZ8+cG42Cp1IunMxGjx6JY4HKUnfZ2/zUgBSq
5azXgnWN0Om6S40WUQgp4oXxsJIEXs6TadMMDT384TfP6gpxm3+gCNaOMm7PqxN0
`protect END_PROTECTED
