`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ViN2ob6j4kDQtnBEVFYe/54i+16duZROYOdAR2n4/nErDFq/3Ze7rs87h+R08DMK
A/SRxR81QkgpIEapv9BdAWvaWHXGqOrwPURHs7YZq6Lwr5LZ2l8pQyEHGij3qe+0
veLSCgGNW78kbtNrjh5cSGr1looqE2ZB60wA5XSq6m5EE55rYXkQXxQKZNObLmr7
9VUmW2nnLIxnpt6DSFydrGlYbrRKwLF5EbhD+wB0GJm/73V6CPTdbkJrgASXpIip
RjaR+XnQk9MYF+zcmppY3kKBW39/OZ8l7XattvUk9L5C0hmSTGLR7VO3UeAROP0r
w5iTgjz1Hw75lVB5sMC8Ma8gPi6zoXdAJ9g2OXVXsn58gF+SbBh1tGX9zJr5CMma
M7LkuSzuVri1s5WNqp0p+PXGUDNolaK9wKnUak/GQBRXzwaS00SbwMNPJdMS9vsH
cDkILHIzwdHE/VUL0mDUOlSRXeehyvh41ih3Y711H2wccMhUNnedKP2Je9PpbeQh
sTjBKwFruTnnalXmKpSez6ON8xSbJHqpNU3BiZ5JGzpwng7392D3ZaqCBUA7gQOo
H+8R4boRpee44myjDqOlR0zt7kGwcq0+aCdIlG35J2YEDfvNAOo2wlaZtYr4J3pz
Ko2q2xzc1b0BujGHaUP3T3WHs48jIE5CeACASDqwqDhTZfViQiZ9ws+jeevMn2zk
c3ucFRpT40JrFleC+cuPO3IAf4Ie+KkYIPyz3uPquzrIdJnn6cRapKgY0dGtsXYN
kO5n+wPn653+VbZ0uPkFXSS525ikP5OAKyMeVLv44sJfCTwlM2ft5nNAOQCD6oct
wxd32Sx+Y+DxALtoc4VvU66o6s5ANf7lthHGHtJ9U8mH9R0LIaCbDCEgI1PQRWCy
kak3kEIo3aTiIVTc9X7ZTxYarRlJcVFtg8Fg/Xzm6zmTAvWg7GAfsQsQ8MyUFgjU
1RhVZUkZhFzmzU+nwgQUy2jD5m1VbH6BV6p7i908Zstci6+9DZfe0BSyKIAPiXGX
xkVhdywchBQuuc40PNIi/ZxZs1jZNUh7abJN4LdUgHU2BedHbkd9u+Eco78yQBY9
Es7sDh4DkWJ3UV930XztFyDNuyC5XB+hXOCpM4Pz8S2/G38nbfKMK1OQgXQ8GQAz
/TKjQP99pXIOZpJOelkzhlJfoRiPKpCVHWSZvu+269VI0UqkmEbEYkeF6zbQbRrD
99dbgHyxT8iYVW7HdhV9kFAvJU1NpP5vBf13b+O5dZxE/8IT1dfFzJnuaiM5XQNr
0SKp5K2BKPuHhrT8MtxBSnlYEUFAZw995FA2Bgyyy+FGd+sUic7iyTAGucrf9w3m
gNxgCMN38fpRrn/tMySiYV3j6LVJENLnv/DgHAFXAg8jcqGk1bxZyF/xEaBfVc6Z
/TpFb1IRTkqkogNUl9MlHtv5SHgJo6jsGE7E13ZF0saK6GSXhji7pw3qlXw2Gqkw
1KZ0ucyX9tVxKwM1glEdupUQ/l0xVVw21OWB/4wUh0EyB98Gign+5F+74jJ7bOvM
7/dQ728U/MDdvvyFeem7zEQH7DzSSnaWN42TAJ3IyNBNCzYfjt/0FisBVlQz09fh
cv9lIW35xPxhHEztQNFp9Pv0zP+W08PthdcGiCk7o/ITidrOtnOLN7ep36fszOmp
SQ+sDybbUeO0Uh8peZaP+rCQi5L5kaJ8g5JTYioZR9qZ+vZgYTjMTKxr6bEBNj2g
/W3Xh6nj5i78O4MKoYAlIl5CxtB83O/nioV2Xzma9ZLUFLlFFV4xq/mYW+zYy2E9
gHKz/KPUpinLkRXyDUGmwGyLLh7tV8KGAML9wEJgRioElO5hxXGizky5UyfPJVn9
zJ/M7OCjJnZv0T3saRfAIMTQSs8cD8mXw6GQujOGU3xkBm8sM1hO6QDPhwpAz5BT
Q6n1AWVFbD2Pppr310Bg8i8l9maZwYJbVAchFr8RxVtEKDjGtib5LjzdJEbxjXRX
TWQhBbFWdrgVf3fI+uaRz5qRDYzt7S6oS+xRLX0uPqJ9G1Pa6La2aApYaYeLeGYf
sZYQLcKN5RSakZQ+Zyk99JeQ8HCum9T2H0CsUzuaDGxRk1siwRJfoKCmkZCx+BOf
6hfkmBzdDFb0TTVAPHNX4S7n3Nf4KSTUK0he+E1eNZAATPoWkr8RoStR04BuA1vM
fCsfsutVpvfvNIW1k1aP1PWbeapoFpZKQljafmlN0LktHyXoB8CDrnKRMv2qlAHA
YqCDxJ3vdmJaQvis4CXbk+EhYpRaIwaVYNDip0oUnCttIeAEUfGb6OUCqrHUw6PF
D6DkMxHA+D2kWNrMZMpKhC27I0HGtJ0gd6tuC9wX89tk4px9ZmcBIpiTPEiGOqpP
3K8xm3un1dqaLNCJAduBz63BotpLju0CXgFJ0QBz2vpT6RP/I2mF97aB9N3FPb9e
lCtrJo4FwId06cOF+9JJkLDofn3H2fx0L9gTDy9bVvCmMf9Cq28jnpTLofXI3bl7
W55+nJ5C36D5qd43UV+9YA==
`protect END_PROTECTED
