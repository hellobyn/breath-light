`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxsmENVTKpcYdhq2hr34HtnQtNgfCaDWyjYZTkIZQ50Vlz6BugElc9x3DYh/8YVd
guiOESh+Wmy8kL/cMivkuEnCI91wPv1rwkfFdhEkRhtA2a95Jf4oMF7JLdprpxkW
2t3zIVPQnHhcW+ztqUreqWHeZJ7DiYDxdYGslHBuhubdgluG9eNgHQ+rwYIwO9dc
X3RglpF6yfF04DPTAS+2yUqK+vkduNm3RHQK08s/qHtkh5Wm9/Dkos6o9vsKNvNK
OeH3GU+nd/KdSzDXboToZTgGZGVHi3b3t3SE9QHg5N9mxuAyZaEfYj/CoguJeP1y
bok4QQpg79YfCWIm+2J7LQ4OHjf7ffC9jU9PF0yhSV+BC8btM2S1M01qTZ5UqWGE
+4oYCx6ZGWoFf0CRFPctYQDFmfQYrkm6Dg9OHkipmcA3RzNjHzx2tWxYPpbOKP6+
zLgqAh3JMjHpkGIBgbwnaFJv8F59yZzqYw7Ftfz2dnfKeXNr9d4n2/Md5fcJvQrj
uruDNnIQ46U68qB7/i7dSTD0PyWTHKhZglMEezITUIM0Z9YAWeMJl0mH1NLlpBDI
SAGUG6TCQ4U4IC4IQajVt2IlngP8WF+XbuYzBF6yU16Jo+3rrZCKCybZ1Y84ZYlM
x67VhWqNdEouR07HmONnXtH/rel4ANUJUt4Cup1h7MFcEVPe81ZO8DkgEtI9wcld
CrE8XWFf5o0Gdy0EHZcNQY8Cw5RHzgUiMCFmsH4oVQRNvuxe1W08OD4fyaXWSfkL
164F2QVKGD8mFBGqQfBSX3qGxbs5yXiKM9b7nPrH2URJn1NyJuNrDoLfPdLX9Gv9
PTlFscYOp7FsMLWbsbLUDnG59ZtXK92VjzUHNn63sfGVu2EDZDbanieBXgdWBWi5
y9ywgRucVrdlrSQy+CUbsDCRFDIJ9wzE27vtY7xGAa51adg7m8m6DXvbSer4j5qF
RTOrRfv1mnSEED7qDSIf7PBiBb2MBIVswvQ7CbjTGsGFLScswX1sK0CDwUBptsqx
iuAAW+Y1j8++/hLKy8H9JNnFHWFNBKShpnmwxU5oDN9CJbYmDceP7UmmarHgXrDb
XFbXx23Mt/SwuGzeihuYSAo6UXcn+Q/A3+c+sSpK9gIYSJcYCmqVNvSdqWmx9sFL
up3nPD6rwg4rmODbj7xnPRD0Or2ep/FLXGUJpmTIftC2X3hgRDXHALT8Q3nO+jl3
RH5iNcRC23Fubgr2gaYChmGvOLUvE/po7EWEY1ry+JAkC7waS+B7XFSj+yJSmkmo
NFsic++IFj6+QqcmW98mjWsMdU9OzjnSizx5AHv/UbDmg2oIq9UOG/REZxmVIDwG
ni+URVQzNy6f7WGpPP39iWdmIQPZhFB8TVhHSqS4+qaoe5Z1RQkyUmcrzTCLluBx
kBlluOfO80hEZQEQsAmfxTAIeCBEPMCfvDnJHWKr7Qu8azTIN/FhElEH06Z+Uyz3
Vvn6OCyOY5VC9FyaoJfK4aqmOF70FgzZwwuZs3dSGAydU97k7CF8vQIznn6hRVOv
7OGKe7LIiRLHjmtQG5Fkk3EaMa4ntY22w0WCIlziS73DTya8ddqAZI8vuwIYBuOA
ofVr9kidz+Bi9R8JVuYmtk1+bf80aefpiqNMQYTkH89X+c9lqeI1lYmDWVfZjyjs
kB136H6WC3UUCb9+CSxPA3lyE08BnjwsHf3TRNltTa3Pmb0qTiMCUy0g+kqCzIbe
cA5DaZBLJ9IndpLpeke57AX1ij4cuao+HSjO2s1UvY2lKICVzFb9a9qGgzZ/cdam
cOd8pVBq6pTnJxil0KE2XqO1aI+5HfGFNLIhZp2rxAL8kPPY9YE94xo1gcapWK16
SHQ5X/OWQsuYJRlnwQXCqrJYrORd66bZeJNpCuGL98AbuB2gTOoHG9wgOVBalcUI
Bu8VjkVgTYMZh3FP0qikkD7VOrP/rMdnyIy6zw2mradGQsPGa6dMy1wLYVbRwZR2
kgzW5vMwlkeSta1RwR6z8c7nxfloa79An+Hw6+B6zOJdD/fac7NfAH5RJ3OSV5J8
u7Ph4vYEXSGM4zlFx0+jXdhWMDFGKZeZw0uBkNsZKKkbmxkmlxkwZb3WSQOOz07l
1Yt6LfG37Hza153K/q7KS+NVi3rmvFQ52xzmx3UW0DZUatf3yqSGoijZQ8ORGXtY
MtQfOpkobYcug25fiiortoyt6Jfb9vCjdPwXN2oMQ/25NeqAcNe22FNwnUk8RwZS
WUNnwDYd3eIvYDgTHmWiw5/lJQ142LutyOe1CbFB5Y9lyZoBvCtCRGk7OLRY1S8y
Ip2izOFVT2XGRRgdddlfdZj/NECaka1lZ8t2BPbkGH6OsO2X/maH7k348EoT+1Lh
kUB1AYhDJmutK33y5I8DIgR4+IA17vDDQ2KrNrEZ2IalWKwa1xZQI4GW3JSVLwFA
CChWRjt/TxWa0f6lIYSbfAKRnpP2yiIgCb0Bc7tSc06/lw0wL07aKMJT1es59E66
gRtDWnX7P8nwO407b3W541zNMa1y69bxurWGcm0wGjhV9v5nqUSKMm2cQhjFD+hE
jeJ4+vu4b60p9LiBKqjDFnOqmRYBlUsdoTmFoxwM+MsqReOTV5S9J8Ze3isBbELX
IEpQ8llo+IaVyuhyErIWfrm2A6rdrlY1I4PhHyxpU20zxth8VUMghtmR9Unitc/d
ttp5aSOnDqsJrso20mIqVO9HB3T9oY/rtnrqDraqw9cPvC/bbHB03vR7tunmxAym
vE1m1ivxTbmuCnUZ2G1OMba29heDhQuoHFZRLwitNr+Eu+NX5fZC0f3axYcJ0GZL
mfuC3x+nhbYL9MVkJXxBCR/J0//cQ1uPVvIusPJ6ofENBHT5HG48yKYf4GEPKvd+
rtxa8TnJK/WwwErafUZGI2+V0qrAzZc6GOdkKhCsRbUmzmTZjWVZ1wFM2C0PHoqd
n1wYOSnadUPHrk65er6YKrbjOWXK0D9FPQaZhUiD3OJrZN+pcDSwGN0FWOLIz3lV
TLgnubRyY5so6mEpny3NHAAuxB9ci5c6vXZYAzUGdK4urKEe0uVnCYkdHEU/jlDu
EE32zW7HcNwtDe4MKzhhimJqNe8rBP7/Q+kkOK4d486XLA8UQ6xBXjW0GAgnzaQq
F6OZ7TQLrpdFWX1eGsVf63U4WqnkbSuHxaXHPgiYIKrexmdx0Vf3j6aDLtea5wNQ
PQgmZe2TMxZf7q30aeTR9tD8fc+Oz15Iks2kPEsytVDxZ5opkGjKY6S5P18YaFkr
1p9avbUicFrFuSAdAdk7hXhFoorbRcFgiijxCQ2VUQPvLgin1DD7EAvb+5GW/dZn
F7jKssM66UNaYjN4Z9JEm44dXN9GOU4hTtJoXV4W0zRD4/OOFxExXkeYtckv5wdM
2z0jHADH7OipFZiG68bNW/ZNz9+KpYz5Wlx39EUKLOth3OPM+MpAtV2o/LjZznOl
3Hu5T5S8Nk5ukGcFluFuCPjc0vtXKNVJpFA5PatWOEmqs23aMz0lF4CP2ThUj953
dVFOwmjKtWCgC4FbqwSBCdQ/iKHCcKe7VVhtpw0mLiubW/YdCjUbpN8uKOcolonD
xmurWs+xLgLsIWD3uGHjKcyh37efsKm/bOdXVYYJ6SB8Zv4qdMdIRZ5Rr1aLPev6
gnW/LC1gLxo3JjiW/k/CWCa6G1ho78uC4l60obmMCpSB3F1/QY18adfF00UvvJC5
9AhZ5eOMFsAWVILKf8m2Z2/A8J2rBywti44nvWmUoYxJZrG7UTXNWUD2O4jAJqr7
IJo6NGRLgT27mLyvF76Xrk4IUv/3r+myWzcA7VwrsIA3NRlpN3PSCaspBc2/34Kg
STcqWPwNAO9YI23a2K6EqQGg6vaPOppnBtLGjLppGS4x/jFEKA6hTa86sFvW2g35
cjLMEhwRQsxMJDNpHzVcY3eyaJLdbDGqQflhJV2IceP8LYuN6uyeB0eiGfMs3fAS
`protect END_PROTECTED
