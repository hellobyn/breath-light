`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNqiyf6AVsWitTnNKi3Ywu2uVjdIKqTz+Pq1P4A4c54xc8KkaIGk5YAmsrMKWKqo
LdthfGLZUgodduydykGiM0IelamwIuJ5yNSrQzb4WwyRxipIES3w2x40hnpN9TrY
7WkU9agdw7CEJnfnG3+UcM6VwkdLbnV2/zBaiiC0JLTKuBRaHy7B57B55Aj5++Zi
TmSrrHJK/xpNDW3c9+Ca76LGmw/ERT11BNwwSKY8E5ovwJE4qcjxyA37LzBEH/EL
v7C3ijVlsLSQdRQfQZ4lQOYeoBdPH1ERtufn6Ll8uMFWW5wZbPc2gfdl82pEM4IA
/giKR3Qhd6L1bxMehzDCrAhQ/7C0uIllAGtHJUM03ijl6NnILLZaMT6AxLL7xguh
9md359/YgWew+5g4MEU/jbM9RPBk3QK/R9HI4zu7XvT0aSZQawQRDzltLKf6MFWM
HIJ6FdhyA4BezLpuL+zVr7o62iqtldI15Yyb+tVgwVbL/HxgZuLMNGtikmuS8Qph
BlNtjocd87eJDL2ygMcyjQodFfkjHcO2LsZ95vuNTqs5I5DyW43dB2jqMN3vSBim
EEcyH/NgdXmRG35b7II1njhB6E6HW/6uwvmcDG1iBMqycKAJhoIXy3ndQK93p7if
ii1+oUBEMhmFy2aZueIsOuwdIkGvdOfZsV5G13f8n2YqAK+3SfikUwgPKRR0EC+M
inTMy4XVLKXR5nvViRGPJSf0BLa6HLHdhK6Gm1Iv37jwQR3fE7hBR4QBov851e9o
I1rAfBTnnto44ru5Q++4OjHi3yn0Xuj570VimTu50OqopbDghgar8HKirl/c+pI0
0hMZ3s0mt4N1uPQ2dF7qDtZ2qtA0fbB/NEDMgKm/DR3RqXsPb83gfOeAGu8kB9zf
eM0jESHITcZdkDtBtc510yGIb7uUxpQro3k6Qx47PQfsIuFt/Zxj/PIWu/L3j8uy
U9dKW7CDYiRmN3jLU2nzK4VAY+30mrP8dD4NXXb+kCaYlTOgPTTFY8Xzj4qlBvAw
fixOk8ffuwVxTGmnd87rXjoWzWnAXtrd4wQTfwmeXN+qh2yHUrcQa95J4RCGmbFA
Upxdq8Phz2Pp67Q+9s2sd8zk2uf5LwYskJGSL3P4OJ8=
`protect END_PROTECTED
