`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUbmCGPrV4UnTT2wJKR3Blcl32zXypvnUx1qEVfYlruVQEnx7dHd0+G5GxKRXrH9
VvZVzddzFGqZCq8wKMBKxUMV1a3LSNBbiw9Ckasam9cuBfo50Ln721LobCrMEKwt
8vM83TknavhjlDsNHwV6FgHa444tmeD5cASeq8sx73AsNVb0FFaWwO1xq8s1dxNg
hQxJIf4SYWVwABBVxxlstMJIr91eaNmDXkKv1AVy9xXA5AZJxtEErKQp3apttydv
5D92t6PdyOAZMrjC2vO8YmvqulZ8ccuW2FMeQFV3DdwZOSboH9bPVh1tbvcc0CEE
ANpVPvQE6JYge/ka1kzQx8NY/D9BIozqkHKng+/zMZjXuk9W9BjkEZeJYompb8ns
UpD9qZoeI4ZsOlA/fZrd7FKHneyX9vSbBWapGCEnwKy3UtK167RdSdFgxMyRzp4o
grK7DWaq+F2nKmo4R0ZqVy+OXEUiMovU1LAeBR7CsiKaNYQ0VsbRcubvdFTxdsrI
scFIRJIdtKI3qPBSJfrhI3S3H56xblpAQzF9ZmNJr7Osy/gjZZ5PTGUXlGoyMOfS
LlMokd226mKdoznITk/d9Q==
`protect END_PROTECTED
