`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76MtKxDRNo53dUjhXRICMrsVZ9V7Wck3x6qFePRLgjM6e/sLtwlvOxnxLr4BEnCH
AOxloawRopEuphAaEZhRgYiSDkEZpEIKhUDgvAS72MONTLD+yKVqy0tjdHSKQMhI
OGHCFP8sqHFxOQm3ppmwQj8jR8hTOjKhzAWaGQXYYa1ylMDsiiFWgdXvXVUNwoUj
TxiUP45Djy7zLzo2F+/ac4aMfiUtK/ksxLxw55UdFpn8ZntKtphL6YHW8dOpgIJy
MuPYbhuKzAVd+Faa26r5P4uwoya8N14a/UdqHw7wtwFspIGAFupq4FczyLqDSoBs
3GQib9wET+ecMmaBATBwZw==
`protect END_PROTECTED
