`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
leV94cl4wA4feQCF7sFh5BLzddok6HRy+yEtbs6BNrcPb+bbvI0s8LgdJHuxtw7y
8ZjYd04raEBxaGB4WPa8JWTFYFC9gpS9VrbjQCvo6Ea/kazRpP+/UtbaVRxzqXdX
vo7nBTgistyQuuKxNPVn9WQKIGdgkP+7z7VQs/ks4+keNwZPucexmz5kDk+RBdxb
uAhYHpj0n5Q8PjXkQ90tb5bWjBhGhYaiJy807i/RhYMt1fZoVzQmOSjPufbBwi8Y
fxvBGpOzG2Oy8lsolJepyVYJFmGu3fTcxIekffzeYr/Yayq5TuFGzLauJUjG8jr+
ntqLQXPjifY0fsCLOUyQGmUgpklNTROKZTeSHg3AQkUUAcPW/fvIQXQkc9zS9IGY
gQs63OE9hTqIb/oJwc/PblmYBCGg3XSSM1kKfHJN3Cz3xmOURraKzvPTBY3uRXva
aEKQH5mJa6Mb8CzUVfvUYpr1INQ19TBJjTryNu9IaJSa6slkVjSavoNPb1Ps0piR
J6V/0voSz2h4y/KvCDhN8hKZtDmaHAYkbr3RNnxeMwDb+xKWQdJsz4DFq/JoGUNa
RQk9ZGjJmSyMCu1Wck7horGOqK9R/hWN2Jwr/25wkebI1eVHg3nLJ1EhIlh9CxRR
3EJZZV4KCPIPvMlC9qYFotGgBGME+roz8QYqu+HV8xIcfnRlv14PF16g/YYW7UJL
LwujVedpSW4zZcO+ZMsRw+iAx7J1KPn2d2ARLRWTi07prgM3VF28s7ZkVNYOc4qK
dBnZ7zxZTrksDpbiYaUHPWoXZK6tQC7NSi+xduw+G2Mn2oBuk4blvh6Ne82Gz6oc
ZSxT3jnqXS4UhP6XPj8MeYVAWpwNtP4wMMsKb05L03mc2AWiGwka+mUVvtXJ13vt
RC6D4O1jXVRrTmyOIwrhXGf4e4OB+ik+0gqYxWgsBKpRTv8ILumL7NF8MK7bbkJS
z2ez7A9U/A4YTjXt4dL9GjKRgd600FtE6eYCpQebEs+v+b8DhcUpiEcV1W5aJlea
Cjfh4H5tMBN8gLYv6SywilVR0vZFqFaCJTsvPcgT//I1obU+KqYvPWESsMBl0aDp
FjcsDAhtNXxw0F3nSU/wQLSPcU8A6imQ7TQlNFrkM86bLzc3QsyV+uORsjMT8cyN
CkT+NJs8FgI13CdUHnESxQnfcLIhE+1dGLuLZ44ZS8K0ENB37XT9CtWiKu9vxdTH
xRQgzSCP/ayfnYGgSHH9CBri2GYmPuta3WV1rDp1Ax8BYlc5PoWtpyI52n9K0b8X
qRCTrKoguBHySXrnvJcBYD9uTrzNmyfLsQDsMPQPzuBHrhY5chh0bcOaxAJS+nVr
Kyq1+/t1kWdvahnY/oc8xPvBtOrK4+oiyPxcX8qOQt2DbQYZGfRcqbpRh/Iz7lZb
pRyugk4imxi9zIQzCbHXmAC7ZRXqJSclcqND/sW0NNWWtmPLLWjTbmX+Yk78Ndww
+oYGGRp+hOz+S1+4yv4bNA==
`protect END_PROTECTED
