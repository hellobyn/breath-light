`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bi+UIH3jUqk5i4YLXjjlGJsiop+U7cJK4XMHhZ9EFHa6xSHyYSqlPVX1tyPO3Rbv
9fQKOJmXMgACtEN9vwI6u9yOoptAUgXX1IwlYvpZ5NLuX0yU/D2IUdgrKSr6Daoc
GK4T9NHpvnDfwG2rGQ9xyko3S8DuBom4dBSRqy+oLPZTPLBc9egl7QqvHvCyEDkZ
QwHtPIhJkrECgz00kXY4uKr4fn2m5AsHr2C4lzcCJ/4UETXY25ASLHHgnw9diZLA
Mrs2JaR2wr2aCHjEtuSlVCY110yMZk/32KAhk9b3ifapRKXjgJJWA6XRBWVkY8FT
m1oNDw3NzQTrokJC2k2+QDvsLNyq0D8wQ4MoX1AFJ40Rn6Kr55O9EZuctsQ8/WyI
Z/JTSat+EQzasnT1946hVEXuSLIcTBVVgvPN8lErKrs5ek1rOOnGZDJOJKLUzqT5
p/ssxxTxbPkKcVPopV3uTizTP1pXg34f3BSmMXregeW9b+ajR9MNJ77mwwIQStVh
rLzoHcC28McwmSJCK6ACoODKzAwpcPMplIRIkfn1giKlOYdrrZa02f7r6Yygp1v+
slvz82dFKUjRlcqivxVNOScSl1T1A6qSyZYnuHTyUrsoHa9IgA/0LJUAGbUz1/nE
mLW5T/jJopqfdifUZ3B4nBqh8CYQzGxtrXq1BJM4wf34qWY9ZoG89BC/r8UzFETK
VgcC9qk4d0vWPevLGpRwK6pyYqYRMHw1QprNXo3N9ebJ0Miq+hkRKbLTqoNd5JrW
I2vPf/oxTdqRZUi/UgmaD8jn2PaavcZ4pquPVhmTlPrU89x+XF7rTVFMQPgmUhlG
H9At/hwItqfvcZuGWxZnDbfnMs5NB7rPe02a2Qb57p0yvU30qfa8Lxbrh4NhARMY
zMkSbOUj/eIKHgwwUhSSctlpjkB/dy/LMWsNk6qcqRy0RhxQi2SGpp/+HvDWL5PL
+FsPXqr46vH42hhqDehFvkhXvpoNI4T+WNEVgRhyKl0sDq+KxCBi4n0Pxw1MzRFS
mKtyMMQKMwcd+6bYW3OlEiQxa7P56hnCMfsKRPm9SPooAGby5Vdb9UvS/C1UpMCI
kSkOTdy26pvnymM91l7Uar1EePTH+U9wXGbCn//uNSHeAjaAVgZIXjSmkKf6aIln
rjvHWfWnf0eMNngjSpi7UozMF7Q81DzT11+fXPFHwR0jUW3Nt9x/HQ7nzhL8WAb3
AP/7nz/aGI6mV5MNn2j0REOt5V9jE2XrvE9gPbGZgGPZ8uU5lxvzCy5KTa0BQWgW
nc+tt6NpNlGwhMxc+JXBci5SlaZxN6SH9Jiu8xH/fdcY3ehC73RyXmboBvNhmCjP
cAKpKjCWowfuhg/ZSJUygphymbNA3SdKuCZGMWFlAlVqH8ttQVWrm+gBL28K29EH
R9Csw861SDLokzUBL66bcBQ+b+nXWWk76VTm/xKa7lAZOho2/tJ/+qUlVtHC9uYP
G4EJtTBIjNxDCztquoIkRNOLCO8P4gwE8buZdi6HfKr3/3aN+HJm8E/Oncn0RhJ6
9NJPSvzetO50H+1N5P+UYQ==
`protect END_PROTECTED
