`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3AdRSTM60/NVITr0lDSCw3dpdzbMK6uGkQVg9mMAn2dhieWhK/iNlxwdE420Hwc
OMYvb0EBeHeuRWb0D9lnkf9wrNFaGrT3Hqca5iUwmAksOYkyrRLSsSs3Ls/ip5VM
WbOJCQ5WAIcq2lxCIQnA7Y4TY4gmCZf6fETZIq/ZwdBXHvHEJ2+rPIzl3KhGjK5g
xnp5kYrqxtYB8I4DQ1G5SuyY9jnezPl8D8jJOIR2mphf9atP6oZChi2tOsZinSAi
Omo8Tej5ssGYNzE3lOk7LaAOrrqftvZGzrmGNqj4BKT2Nlh8GAbzxwURtnGAOhkF
XDG+cnZFlClZtm9skBpBS/s8YE6D25G0YxUe2U5k6+JnFtd3VBLZxB4GXroGg6xv
iGX9e+zGE4cOnNJwPo/sFE6OrjbUwHjD5yEFVdZybqScBs9r9Czwa+Y8k7Q5nZhS
V/BTmySCoygaGdFq8npHX4DAzW8sxMOV+8R3QV1kkNx6fp/TC/yWjEARbJGMgM7A
7/kywrWLC+XuR0UcdyYymXja8cuQApAJtTuSIVJylt0sjK9TOlKBVgY9DgtJKNKz
g+8aaT8e3/zelh2SC8HkXMSNFo9FaFvAjVd63QEpmjkHnG7VCyt3t+javoHf8fhM
kBXlAKVJHCamIIoAMkeQC3pbKkkTmvK1YPTY5ay0VMQ6aiv+8JlYR7fKUPDNTG5t
P4R2pfdGf5yM23Lan45GVk3/ihHpN69+G8DvTEV5hgRy6q5KbTCuKUbQHAy9oezL
PHOn4JFH9GS4CR7b2wi8FBv9xpYpa//uSpFgXsUx21nl4vbjAMfhQDq94rDNt1hb
7y4qdeY3ZP9ToaFARYSF8A==
`protect END_PROTECTED
