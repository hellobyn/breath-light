`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxzFj888I3GUclU5SOG0abBp6Ep+r6G8zw2HWfNYCQQXrW94MnaNx8O08NEDuXWt
ZmS0+hhLIU1hrXPfg/FVb0Rx6QmmLOL1dDUUfgjytVIXv1ZxfdR8A76h5/57r2b+
MNjs0uosg6NzwVm5Jb9shlGJSGOFnNqMZ7O1VgGeQ269j+vFelutzyx4ZXuqtLI8
SAZ1KmmHUnq48XiYt+ZiYqSL+BpN1oEV8k0URAo+ivK4LIQ1BYoRFNREMx+UGQAr
uVc4rBrGL3S1ngrRq+X9Vn0A4ShlSVVe+5RXfXQCvvL4fby2bohvxsgQNOqQKEst
WfCCytXVbU8bQcOhzQmdL1YepaCHVF/4pOs8GQtpXW5cgMN3D32cQc7sE0aNTMFT
XNJqmxexOzZ2U1n4XkUSRui+SDRWU+IZxelO1eTW/sXO4k7dxQOLsx8PfsW6klir
n9TnavloYFrlNVAPPUMKE4RymnPjdIdvkZw1NNQjIvYAqFwOkk1DKYBX+E2BDhTH
G+vJ+NLcaFeO+wUPl9CMT1BLELHLe2FcZRaA+maXV5oGFDnMFPaZjbO0lJD18+u3
OCxhwQpTEqOIG8OnpIq04a/TCAT6MJiCoUV274sXPSKOmvTMiKYV7/EilufhU6oM
iWf6Ckmn0BRnODY/WuILiWouU78HvBhwOAfQrW6JMaGyWYoGnv6ItTTFTqXRVRmH
Ss9FxvR4te/ynl2vo/owGvuvECbHJN+pOOujKTA8NCfw0CqIqMo/8+mlZesDcScw
DBQ/xW3Qdwv/OysBN99MFg5yExw5NgfeYXhb7DoyRwLckVSwh41Jap/cj12XGPpO
dOy3vWI9Qu78fvK68oqQa9OAVLpIJ0O+0DAbQW0ZcX+DFB0Sn6u/7Qan2HuSz6Ty
/TKxxj752A7gewHqIE/40HADkL1iV5OBu2V2wbpnzZb9Jp6l6eTo/btgwJtGPPd1
OLfSa/veIC4NJJEsoilYG//iMHNQjEGF7LI2pIoO9lAZBdX88v701+vg9ikqWFgR
EgBsqlNdVYfYv1ZYfJiyS3dIdHyV2CTaDIHOml6hnc1LqrqdXzHAakr1uDhv/N7g
124yu7OgJg6roIx66FVeLSw8oRV5wY0woLrHY1uoMyNMW/5iiczupyC5ej7iPUzR
HkeHqh9foZnnz0HYZOQpGs5PTFZMNpJHIWMSSz4N3esyKyg1eWPsNFAqRk5XUgeW
3I8Tt1PNnNPuDh6dTKfanUaVOMIZ05eml8T+g70/bnAIAbt0KUYU56mLNqKecgkc
meWyt4yTOJ/B3tUVZuFZ5A==
`protect END_PROTECTED
