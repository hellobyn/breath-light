`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sv85WfljkkyK72a3mPHegDmPEw5GX1GXy8FEbfVqSVUOL8FOOR9qYenvbdUkJw7
yjrq1qdDrawbxCawZY90EgWM2LRUEcqcCxVR5b8br20JS6gLCZQ/zw8EOVcQU1Uo
yr8vH4Yd4ebeJrclb7zcx+d7FAOuAden0ZhDtJ8y/jIxfYavvbV3yc6TqIPcRBdh
HolOlkIT8JAZxBr6wKEnh5+Dkbecx7TltNk6TQBS1Bd/co4bK6Bh8fEflDWzP7dJ
3M9t1AhclJFFNThdwmB7wz/f34lJ30QEGHSK6F1VsjHZ5PyjUlssWzQXAwuHD8BY
b4bmsBF2uzI1/qBqCADv0wyIjrKXkyYuxEaUS6xy5XvGol47x7e9Ly0ZkTNB2LCe
yrjAtDPCS0P5KmWXPUrm91mhOjBGZPt0Ey2vDcPiaj6w8lZrJevg+kJnK+AJ8KHL
W/D1VMM1r3suqAZMF+woOsXd7C3WPO+neiqEjIqdBLzQVYPks/XUq5vB+XOmCs6V
Hw95fXZWaFShwBCCIY4bd2RwA8c9NMrmM9pGAXDymwmwk9UkgSnZMlwu35z6baOn
fmEBYwzfo5IrHPZF2EGfYZ3MIWGHrXxHXXZ3ko2Jw8xchw6Je65WV6lbT0DvpLCw
amxlN8hdrY8rWv7LDa0XvSqOXAH/hryi4ykO62UOdb6xTwx2P0KtGlFxWKVQwmix
qKjoPyfmD6ZU3g3hAYdN4eLMGIoVkEzUp09WswitpIkNe9QlAIH1nGmVYmDKNugO
uumYkBlOHLRPlMG9cZk6EV5qcp29YCnz0APboaRp8Nev1jSe46INq8NJiqyKEW1a
B0UZLx1WDspXOR6+Jdz/yhnXlJ0qrGOoYzUH8o7KIQV0DIJ7UaR3CyUaoQcHKILe
1E4rdfjwsa9uEtVTTV0UuTnsi1RUmkoJI2B121kupg8OG57wrKEE0M8LoKN6kQ+P
qI6ekWYcmSfpv1RGqgS2npl2Rq91OmyHGnmQdwcg2wKNBkjiqcWJPwZFiwzPQXXe
ypRw4pTgTp/0665Hm4uru/k3S+/Ac8sMAofBEwaz7c/XG171XbfpVVlv7XfVcs9h
cRNESvgUx/moCFyMPYZYItezPl4658fZ+GYOH5pTiP9rA6v7enZ64c6R9WjCs2dh
Pp5+FFtXxg2ehPr7xbGJ1+gRWDWVMtOB6nru962gSu6xGRg1xuSQMC3YYN697OXl
Xta/uo3hgS5E2qlqJzkntkWLSUWqH9Ptkr9uhKCJoD4rAuVQrtP068+XQTdmTb/k
STZM3M4e6O/tBd0osFW1+8BCy+MAs9w6FSgkvcajdoae2NOD+ZCSwyUoTJIWPy69
FCldVnlxQwZRgod/j4xgzwpfL88Ri/jLIVNraiaxBc/713z5d2fYiDCq7wGbY3jg
HqjP2EVduTcQZeLTfN9yH95/oTM8ZQarW3C4osDHu+OpSI1mbCsHTvxZjiJYug9x
2QFioDqnIlSDC9CvHI8vnskRo3VtSzV8AdrZl+f2T8+rTUZDADuxXzdO2sNIyEyI
CMV7Y6KA98w/nVzo+LcwBDRJjaUKRvMdpLSc6z6VDpXLcwk1UTFJfdRzmj4YXstx
dxa3VieVb/xNkJ7zA8SMIyoY8WOAeC/EPLZK7AEMzxmwJTSPE6yerlL98mGLk0tx
VSfdnltCg0AtMZzDdyCYp6QVlwpLY4etzh9YKrAqPYsb3wkm2ROEgAzTddgZihGc
U82lVYFef7wqxZkSfvVsA5i1UotIdrug3hFuafRyFTPFIv9FiU8OKWz/Cew9eZ2c
jRrk74+rsdd23yRBJNRK5nTxRKxhATScMeqN1PaWCAEEAxUhIlhzVsU/Kk/EJDJO
8TTkr6ffcsWJQdsLcsl0rr6tkAbjaxf0El0sGPvH4SCt+mNIYqTxv6fipEyiNfoo
KwbYnPOXKW7nnd4vvzzBxC2qULVP+JWCLhh6FoGjPvJoyI3ctR5PsKQFubYmaecq
tZT+BgRfg+eyWAEKyr070Q5M8puDuAbh6pSRs0vKtlH8dwKU5qhXz8bK2DJZMy5H
o3Icl2XTFfFeGmKmFHrmEe+AyzCK6S+wpply/JGDxm55CLK21LK+Hfdf+WX/vZ/D
qPSx4jSpxIyTwVHHFx7JA8SDhxao08xwJImA75H1mW3RXsZsLqevDBEJglQz3oX9
XBzoujQTBR3BXPuKnizGcSitz7FaGI3IHOOIBPduad1iRFRhnLf7vu20BOzmDv9u
KpkMAAIhNdpmWKyjgm4K0Esf4XKLuoQMfFEYe7WcPpaLQBCX8GnbLYDkJ1ZYuoXQ
QtidhRV6Dk1b+hA4z9gAERYNR5l54G2TVkTGmaiCXfysrIPyELT4D6nkiCH1dui4
ieYyjNOVTI2ty2s88YXFHLUTUkGivmprSfRpHjEDIA2BhQrEMJmDiRdG0+f30Tgy
cDrC1Kj1cP8oy+eAFKU0/z6pS9zvHI/wpvBfbDBFTRj14z+je/3rPJmCXcX/gfqx
7XmVuhCSbxyKGl2hUL9wErseOOPFJHj4svkHN2oDsW7sW0TumWGqHeMP17nF98mc
OPv224IlntNKNugIvtZyh1z9ExAaTxzI3x0nq3KIWECsBHHO6BWzHshOrWHqIppM
wW+UZY6xJ5iv0pFLNpfOVf3OrpWBvxhiaixK/x/ueFAcbq/Cv8NGXUPZbmw78Weu
SQqY1WheVR7D9X8iJSRCuN9d+hhWjydUK8T2AwGqL6aZkyo7H062eFBEgvMnwHcX
4rqYxuTETe/dgZG7sGBf5+xGkq/9QEIr9J0uz3YSmRLzzJpjsatoQ8JUK/AwSO1T
MneKqPBeu6bp5/6C8dmv6ZKDwxSZj4MwlAHtYAT3MhIbmss6k7tXFPxLcAmlhiJL
ffX/kbMaFeHMAr1n2jjTd8ytcr7HmzpRWZrimGE55G3pvLASg959k+RGxhGCXdU6
oWsRlvjBXmWcUmFCOQUpSi9Lw7eIOrF77JsLPy/+9tWnHH2OC1q+kSzEbOdNjB6o
jPunPYTxXwTXSahS+rVPV7OviQdsY9ahcX9P16VR1BlUFXwOHzprMvkM9VEBmlZh
mQ9CXfSuC6W9NndZCNGWgGBrHo0giAR1XlLXeRhaDa/sls+6dsenISHbf1fuBLkf
84KK15hU/kA/yFMXznLKhNMQU4KF9KMOSW0h3QdIXmvKB7Yqs9KEa+2Cm7R8E0cl
I6Ua12ISP/Y49Le4owFBauAd1vH0wc6ME7u8oH7Pf7EvV/42IpcTcQClCsUhE501
ImTdWTt3G1itWzkfHj3phdqBfP0rDHlOzGRg0tmn9KmzIa9tO7Yb6KTbNcyN/3Qh
WPY8gIfmqBsIuyESjTd9ashetrQ7iB8DMlF98kEAc+FQQ4Iys3+86EysZVGlWcIj
HHtqDl/5/FA0nmuTMoeTVdzvGNoUHp9+/X9cSs3T9tZKeeK+mg790WMlrrI3eGZ9
JBs64TuRLONxUfj/4Y0nQxx5RVLApHWaDHd+u1C5C3XOfPKKhUtJduqKh8qlKOdQ
kUamR8Eso7ud511sWVK4DrOQvAzGrKl8pkjn891PWEP4gf4v243OGF41nE07sFvC
yssVIACZHiLi5cJZlInlgnBhGsLjQu67jotl9D9eCeErJ5SBkHqIYjHMHQIAiQya
FlHOdABPOdE+prR/vBkf9754xXahqJlSMNnZmeFvQjtN+fjMt3rhAnvhPhtZ/1qN
uaGTNYNMEiPwk++EEg9gKT5Bz/Kig/oBbnU2pGumiMm27w6Ue9N0SGhJIUvWVS4u
P0GWYX0GO4EQY9qV2m3F8IG5FpTaSApfCl5x2EA5D9ld8FzZVqJywHIstrjdWkG9
TPQj2YD1aE4RxDczcRqN888tyLb/7lp9CRVYpw+R17JSbHJs0SAPPfSHdnRFuWFf
rPnEwgw50KLjN7Jlsu1wsMzw5tp6D9kWGwzyVSXMLXhkdWPB62UI0NozU1yRQoPd
IhVMf+uPzrHHJJHKA1r/CLRWxKMu0N9b8heq4vh4XxWl0wrQdFAwl5lCYdBYnv/x
hJYg4Yq0KXzfOjZVzxv8vQo1IOFVhMCYvyb5FGDO5dOcUjn4FOiD5nXiejX/2q+F
g/WtPgAOvlzihFdkjnCpfDvueoZjiTfnOeDkLIjSY97jOFFi0w/UUzUeW422L1sY
6FyTnCrTXV39Ubha0gsmEFovyIHWB33JDp0Cl+Z2mqb8N3FatDWL0CZ9+glbm9K+
zIW3dSvHV9/FXmkLlp/NlfYX6vP19kKypoZ2i+w/KmxsfAlO7f5kBq0vPetAXqHA
ZD9KQbmxWOGJz+wHnQwTgNwZbnA+xyiN7WXuQ+2EGigD+v7hfXn2M4cHy3CroKWJ
eWjKjkZj1DPZV4Yy63+wH0MzE8nkoySAhquaT+qNcgBQBsXjrVJ2LmieJll9umGR
Q84BDRvplLuBXwzcVPFgo3O+RmpTVrtRNcTVM2KcED/0ybP31D9pwZlU+s3tdpkO
9SWi2HXrUdEPSPVwSitYkatntMIduLIIDymPfjREKy96mjlnK8ZMQQrMcOAfPcuV
4p8k3gMqw6wxFwaQJP5vwpvN21tL/oD2V9F6kqKkdujG7FhDTOQnf89ceZxa6DEc
ey+6nJHyxo2CF0YTi9XFwokM969ugU6p/p6AyGzBVZHHS7wRLTriWzNqJCAceOV/
xMPOX7b8SIWlUUc/N4FwSoq7jSqwGqfQDrRJuMS+V9ab54ZeFQD+sCsrxScwDNWq
qHN+Tit3tVY3p8MABkXrp+AJkhZy9STVoiCE+vKlY8QWQ5+6I4glE3lWyg0YsTf4
BlSZXoOSplXleShKoC11aiZ59exf5R6O2hdSMmi+dPpBpmBWONODZAnDO12H4KRp
Uy5CDxwMaTb3/Do7suK8nfWZ2SkvXAo97vzp3rWmvMzKaT0yQrZz3ZevvfFWHGH3
VOhfcSFOdAQBVNO1hkrCu5sOneUzE6Pw/TIcG+quAX2xfPg7qcxGH77e9MSm2Oq0
nJaPGxeigsoZzJ91V//hoFnpZhlWj7DAGViIQqtEY/hqGJO7jK1Fz0+oMSjNEEzD
S57izreXUXIeJJSjPcpyI1I8Cedd5n5SXU44LQEA12vw2EBygG1BhfoQbzu5VufG
87yIlNBqz9h7bLUU80wsoBI4Dcb7/vrRRd4E2CTZEkf76aPvK1KI7LekqdKem/0k
EGfoQjQ3pxfmohfKmaAHjGxYaQxlkyJ+HMcOre/T7FEBx9aJUN0BemArVJtBi/fD
lyAfdnu5ub1XAsHMxjOmGgcJVgaB+okoLxe2zwLnLJCv3tpi/EGALbD9gennbcch
1zdAH8q49bsFoLyXDG4h/0q2tZ57LvRsUOTS++0mplaKfnsy9I4ITCm1U0Fbt6HY
EsBDcw7+7zJQFHjs9fUYmNSxuCqI36se+Zi/kJKNUVyg+Omv8pOLez7eyh5F4mDs
5JadAr4LDRBLUYGiD112Q1lIuWF5euZbwI87gSnp7HgYN+9xNoO0MXF/kTyal7ek
vPbWbGeJd/tMiIiNvwQPtsJtts6l46wgb9xPM8kx/jJmP4aXpP6FmZRfI5/qh0Yt
LrHaz9IW2HrWXV+c87Kwq4JQDuIL4wACu10lFZdVP+I763iqOfzTJw5++26NzFWa
ui+MBS238trOpaX0ZQseG86r5YVpLkDuxD1cJCpaMNZBzbS9CEcvRCl8pSGzB2gZ
BOubzqEWD0WmajZpswB9iTNyTiPkpV+G/bHta7lVyk6tYfl0BTuvEZ/MkGoooDpl
HfcQiuC4FmXt24Vq7PhO9UEkbvCbbeAcH1QTN02dT+5O4uxCw4VJj1ZsKuxdK3yh
zLfFwL/OQ4+DgvmNNgCi0vs3wySfZcGWhbHzX6maaQn2vw8Myq2v/3Sz3lv3u/tN
6a+GcJW9rZdWBM1fLDBrGb4cW13uhDEawKKemfL/esgzid4zYRZ26tpX6SuSyhPK
rleceTDN561OX+X/fzkGlZ5WUaAAeSIjrra3aknn1DyKpmfZR4/uAtefQP0K+zTK
0bz4ah1U0q5rQV+g1/l9hp+mJvmWLvv8arlMb7cdDvy2rialJQOhNI+10ET75r9F
Bhtt+TiSJ0gW2U98VsQYysG6CoAsrXa7ViBWvRAWefwT8WHMSEue15Fq6b7XWf4l
BaoBLSWOS14gPmZqXIykteYZRCmhFLcSpIuKtTFplDa3y2HZPTwu+p6kFZYM7cly
l9fujvQFemJFykPQrpr398ik/ISVs1xwZgahlsuCe2sJI9QZpLoPYAWCNC5+PBxl
h38m42uAHKEHmruHfeW6bjDdwqToAwsAlauRcpRaT3vnwfTwroxtTLUJ2YC1XEbW
HJ5SZX85m3P7Q7oNN0ufB7ogYKrZJRP/B0uMGL5rd56mm+dCkq+xhKr8qPOjqzAH
7s7qpKydie3WfcPkSza1zQ3mXla4Wo6zfM2HsIkA9ZyY8h6JRreYOLubl14Eg2St
BeNUl+RLuezvT9PtIt973Iqz21JdS6SZMvjmcxDsabC/wDUQgn42uB3Y/rhm3zcf
D0GiACMps71Es4a7qfegvxRvWC+stX77tw7WB28i3IcpObHD0kEVBENnVtwEFJ/n
nw8/TAz1rCMUqkMZDleosGGOz/+a31wzAfMKl7l3LIm1m+8BPJTsABKwR4nJpbgb
NiyRiKycK7OOW4Xt0Iyitmv0+99mY29yIZGhnHrgBcwzF0insZGOYa6DAjw5O6td
U1u0YCp9/KMNpG9tZd/4pta98ZphFv9xo2Dpe9/p8CQtMJqZYu3nLE1XnKrTC3gY
cHLGGdiubC8AyQJOZIirCFlhy1W0vG52rTrgZNO58oKd81EPwetOuJirQ6h6fGDB
b5kkHVQ/5HgtqP2gNUn1h278NIZF1LNK7V4TIf0eub0wFuqLyNwe9cBdz+zSXNsS
zi7FutNtMB/sX33S0/o/yNrgjmBm7usQrGx6lw7fATAqwTtj0YuHxX4wqPpf7No2
l6fziO5V5ON5Dsb5iAM+UdQ1mCP4HTPO8++ZKLUSe34U5iOi8C8spoWNRlF9BrNK
bnwCM7hzYYXhj1IRc4AQYujmBh3Bv5Z2BErxVT4oKUDvu2SNmS8PmU+wd4KrkMyQ
cnjHmNgImZhNEN4IHj+2nlJhgZg31tjKovGjaRjum6ksGIP1nYEeuzwyZsZdf6wn
YW6oe9HHg8EgoOF97IiECcwb9vfL/ZVObXumdjJ/Ct3sJ8EqsLlN73BIgMkiGfJQ
c4X5h2NWjJwk+H1J4D4xHJkXSNCDsVY6/jWPgq1kjp6vaqc596cDNpNqI+BsD0ai
NzHWb1z6bfFev7/T4mf5g29lFGLYGPgjC9RS1G8OI7eJOGEgxBgDQbQ6XVD9mUml
rrup8r4UBLQ3j1mY6FNd0WBGtWSF1U8fld2EIcDuMr+yGiMWbFQDKdPE1b/Wo1qn
EA4DY61Lil43VWo3YJP4UqJfm550zc9KD0Kt24WVfzNcCfydQBqyonvGxTE9PzeZ
3ze9VrzsxqPQWO/JYpS9684lsKPNeju1L35zO4MkqHyn3Is5rUNbawt2s2C+Gz4F
tUzN9Wfv7z4R5x2lisFL0KYTkJvlYEEJpbwkrl2qbBWkSgtq3JSsxZSZGRJdCgCv
BuT6tBS47YSAw5eCK/Q3yNYvK0N39UwrJVrRkjDk9HEhBCx5lAOYf+I+yEp65wHZ
HC78rQoycwp0+0PMtZZeMYQZX6192JEuG5TZFnqMdjTIgk2e7M9sfKIKhyDRWPzv
G9urS1K9UmKrkk+3W2gTRIEKEY69cQeABbLXwBPskZOJ9yWlhdWzassB09cs5l7d
Z2jPAQI5tRrpMzJRITET1Cz/27ZasOTII9RByInHp3jjaKFozumAekF+VLTheMHT
j7vOzjV7C6BIQ3umpOS8UoU2DiT5p/9IJqZuLYDxh1K/smcYhhIm0E6u7ou/4Uyg
l3avI3Sw9fEg/k0tW0wXb7qnygTGTm/kiQSLtKgBZwe30NCvp5KhLDZ6DT3rxZuE
8luFpzAfqf/6qRB3bphPErs3j10S1omb4F2cDFXiTsAb+TAtzh3VzyAxydj88cJj
zDX1B+U/WqFm522ODje9R3QIkksaKnRb3k6G4L8EyJmafNntsJnSTtzVM7dqPXZw
ktMc5WNkVXwjiabrBm+Nv/lOT+osueWqnZtWECyQOvpQWJBqwfFoXOf1N4hEkuO/
03KWOSIyB2jR2uwupGfOGn1FYGKR7ZRPPBNd8751ubFPUcqizVAN0MMDZ9q2onAG
CRoJut5PyGfBLEVz0bZa48e03YvFOm1P9qHhAhzKFvealZ4kZM5WRLy9nd+x6BXI
KXaBFxo52OqaezgLlEYgptoOhuK9SbBasa+e1ky2ENw2Sx13XbSBmbirVtBU3VT6
hgx3EtWRwf3NcCeSHqNduJ5s014W0TCmlN0sX7kwcmJCUZIwm12zjPuL3QtqFzA6
0noDK7zVSbd/bOMcfEByjP+Bwr0MTyFZbl9aBYZ6uJnCcbmr6IPAHLjxCRy9jmMn
mZ9CgmSMZ2c4PtWfyhSj2N3nLjYGRO7ptOcFN52KPOvGHUI79ZThz3FZsxFstSea
n7dbUOZw/QOxCcwW1y2oxmQWq/RULSkrmVuzlOlqY3rmMtbmm7HRr+cTQq3ywHTA
8ldIXbPvf4e+6hs6qOHQfe4YeVwUWx49InVswno4mk35CDBUP0lGwqHtxiCIKuwE
lAf6tFD5SRpRpYKqgxwk3soH1sXOwKqTKpdTEiED7o4hHWlCoe0HIg9783FAeuyg
4JIU+XPGAQN/OPTDAgBuTL0uTFHkAyktUngDJlIOqgeOYIjQl3L56wFSbC/VxDTz
BXjUPNJzFS7GQMtkVcO2l0D+l/I2jbj471kFm2HH5mDIU5ArwCNohS75Uosox1jB
UkJiUENIbZbg+QJatuEWu+PIL6czPWooDxN2cZS1n+C0ywHEsaATVsBpgCprVdLj
inrigO6Dwv1dammNLVZ1L3YZeZVgn8UYVcPaj9bk78LxzbH9BfeJJv6LQTTonFi2
ogj0RcT1f23pCp8x/ndd5syv3islqMzv3+nddC7wXbQFypI1UttEVT+STjsdZYcA
TZ5DqQk34JH/c8bWwugzL+QM2/9aSIu1FSFZwQ8hC2w8kze+jZ0XLTD+NTSTN07+
SgjNBM5/t4Bl52Grz+9uu+GtOyodZl8+7KF15WUm9Dkqq6wC2wmCnX4JzM5zhcx0
c9Ht8LyLMlxJsNg9Npj1/k/fJokNV6mRZJ430UkFqYI67AcyM3/daEubEFTe1CJV
jwORn1P30ZrmyhEA+aRpN+PYccVTlwVXH+uRMyByTtJdwA9tdlXznotyUfWVO06L
fA2cdUTaxfTWt76bahtPUocgkVPSZaj9iFRb8eJ+mD1s0inp6SbLzfvDiOKkt30H
7ZlXzxYRMSDEq7l33s4+bxaw0KnYXVShZgx5MyALNr0JKCixPZLrmY3O6KF9iMEM
VuO/m2jm+AVIK64Ej4EphouWpl4tcnWoB0JVT4ZI4uGfwmo7vxSJ8o8mmyaEGGkR
oMKh7scndp56ULBfzqpu91qB4zvNouS/Kzo60htIEerCfGb0gsPY8CCI/Lf+WQMa
vq5r1MtJfc46durXDWrgbWjjKg6KvDRnJyrNzv/xQjFI4zQRMhzx92jmJrvvp/ee
diyYQrYS94eiNKkzJBRhLQH3kvLYsKS/7L5cfYFncTm45nK1f6xjtevRWCJVTyZI
6cCFCFyuEkjAKnR8zSVo26cY/yHhp51kEkqbKCAyRrkkBPatXLIgHuCjjzcJ9Q4j
ZmvoI2pzai/5vTi+NJjF0+I1fTW1RpwsBsQ53POdI+iscsU0YUBG2+LqPWUTL3zs
fKdgyftcYmFa/XGv05KhTARhllrEu0lDkhzzkKeXir+xHET2hljJL644Np+dFOVS
BlyOllqQGWpqNAvWgqgHhyxslX9BwmV90ks6vEf9q7TWQq5pJrl5giHBSgibTwS4
Q9H2wX0gOt+s5RJZIcRg6L32p8YegWu02Dl9dL1xbmSAsLuPjCraWA0yJF0Ga25Q
MQYINBelBr5Ev1LhHBwAnEvBVaZABBhsEvN7LZiJ3kUf4wA2Th0Jq2ukBoeHDQ6I
xwnSM0Fm5LHKvooalqF2aRCQTyOC+Z+455BXQ6GbUzQ9WlJ+kmKFfnRR76VmIw6D
teNtzOyK9AQyFo9LdUN7EJbdCSMZdffVDTBML7erzMCFeQNx9xaObCpbLeN+dLDT
dFAy2fyUTGnjk1biB9X7t12bhJ8Ry5vbYmO6MEvXu+zI8beNnMusvAG2siHZL0dP
vNrtmbBpX+2YPiz7dFY380ICLTYkkHUaNGGVFhXVED73ipXBo7O7SvKrGQwTvA1U
/LQwiCYItossQ0OOScEbjMTQuOquTYNy0jDDQSUqRSj98m8gLKEu8MmplMKH0IfD
RX7yBMR3ZZ8c4qxsk6NLTKoERDKd0czLVg2hihALAd55jh/Ehlsm4rOzYJtYn2JM
O1eqZ21cbNRtAURFBjrnnOWvyPyfEe/qRn4XhiPDcP769tA9Bq7ZGaItIJsWno4A
6BebNnvvo9ucBjLhg+klP1wMV2C8IMzN/N3BdBXcAwhGV407Fv//c2vJ27422VCT
F4bBWsf3RydMzsN+WvD5CVekCvgLS8s8sIAQiZ6gck+14Ey9Qnlo8xiMQeuKEAyr
xSNifxyCgTo0IDOXF5udURHPdUljurAZlarSZyZPxClqh+8f14ohpR6nLvSJ1sy8
gOtEF9TcpLqGk6++5KQX/lHSF/2g8rtJZ4iGkS5b4Z8Vpt/eEd3cpBw54uQ3xYtL
gZQYOo0E1YQJgJK50MMaimc0d+pLpElADH3U/5zOkYPwgwX9ri+B290Cwm+d7pLI
MVf/gRQHpk6Il6zzXUJANKGfmwagrO2ZRnv1+oF8rQ23Ncv5KsdlIHfYW0ovLeLy
Y9FU2E4ao1sQgJvDm4AAwf4AS/+O2c2RB2Emjfh+HHhyQSR13g7OsgEy9MtYLeDS
yjTMKuxaFa6aBJgu5c3KCBamLzu4oMBliZQOFalu4WmUEl6JhvWCewIAbS9LHoLl
/ALk2Qw5itsrqqYm90xyyLd9LltdBIG7koN1oBUwD4ow8eGhGAuw9/Yocs7lzx6W
T26FJMuVCIrs4m5j6+X/0o0xL5K1deBSkqtwzBfsyYgfDZoMFR8mHZs+Di6ZcgcK
HvRvPhDueX0lnRewKpTZhw73x1zTvCinxQc5Uvhfn7qbeGzwB4RxpobBUSHAvtOz
XHsdf4lSz3ouFpqomKhDeIvKGpBqJ7MAj9XTyCOzQ5NkcICBZgI1ZQ6yO3Na486+
3vaBqW+iKghc30cCE8ov6WhKfPdREGevI+se0HVXmIlMzbiPGYWHb7b76V7+S2TQ
/7EwvoFEfSy57k3ULNQokJcabOgnkexK4e/NLCIUCuR3f8WWBxg2nIxFYkZccUR+
KYKg0QdC6TN4buNZw795j/FdnC6IwRbrHFe5+h7LBEzjT7e6yVNFHSgFBgD19Qw4
RCo7m79POZf9dLD3B9ePTh35c2QfYv1aKbV2PVNw3WtuQpLa8SwyuXqLgWznBFa5
eWDkjc9I+DCpwgoMQY22c9vp1ItLDkcHRURlXSmXgUiELCUgHI8Qk/ukzElXmli6
03lT7KUxcOL3Y6zU/+PqzkMpcry5B6Y7qPprCKcWgJgwa8attuyeId1TeIG30SBp
Q7julDLMsH2G2oPbewsxvJ6LnsWy8Kbr2t+tsBTBLe2Jx6yzuNGBIvMlFvS1Jk+4
yS9q677OG0rkfBksvVcAZIoz7wNOUbTEjtgbMIqDReBf7CyDNuUJGVRELVjV5FfC
PlRMK2w+JN6O5LxYYJ4ysuyyIFCHBtO/BW2ChudYCLWAOPIdDPjgSkiGSXrNMVmi
L23Gq7/UnxccExEXb8zQeinNL3DZIc2rUIs+cH8eO5FyRyLv4oS5PMrm6EgC1g4C
TCh9Yc5GKnkMxFYp2bnj6q81SBD8mwpN7c7SjwX7uPus49zk8t8dly6OkYFKb1Lk
2YnfbbipiaDuLeJv6Yl7py2kxyLZJX/qf8o8SJW/uaJy8X4xP/8ZwfX8YCqXY/o4
nTvo7XzxgHhfD1c7UKEWWAP+yCtp8piuOMjS0+d+t188GoHLzbtXtm16J+h4/0g0
f3+E1CbC2/GwHi7mV2NsxrvPI4oLd2935fHEhJ/xIKsqwE55d22nZPdLU5QQRjcT
BLiNe1+wt5oyeWi6ce0sLTqJkAM43ld+Wql06jJ5su+O2mLn205ixcCkUXQ3PReO
s74BnDaM6Kaeh2xgXusJ3W7FkIzLgV87mWY0Ny8oPsMqM25nxdx4ZhoA1I3ENc3M
yMU2lwdpJ4dKsE8WR73RnMGWrBQ7oqNUvZUUF0NAVC1A414ti04rlP2uxcELQh6t
fYjR21WSEAvllpbATY3936VTmRleIoegZVTe2nATis5rVH+WxqluKqoM4l6XSfWL
9Tig95aO5lKUG0ht3aY3i5Bpml70ow1eQNhoKIwGSzL8wBreHMpoYd5qcjaYVZVw
XPqIf8FwYEoYQqcmRWxVhjYFFy0jlbgF5Cu4rxlInWp3hqTahhq1MOv+aiW0kgN+
PueAFKZm+0qC4imGxchLmZhJDYbyAJS+xkmMb91QUwfjczZvSgEhP/pbyrFtH87r
7EhJrWG8Br0r2gq8WbgSkW15wmMNTXrcGmLdR1m6FKskeZfwL4PA3u0LYVD4q2Ah
1/gjrwWWKuEkjV/e8AD19q0s2T8vZ+81YXxIXWP9AC684l1Yfud+xAKbgPrkQUZA
waupwzKVReD7C/0Y0Lsrl0QTDzg4iF+BhUkrHJBoyRWdsz27d6bNdpgGy3ImV3o2
L2fjGhSVL6ptNss170m+BkIvVnXqcqLI88GnFphd4sAaFI4NKmkVy95r44wK8iHd
Twlho2wHrSqdZhoUBxq7fTcjw9Rq37Pu5MpUmxGwMp9AIcMbFfidbleWLBeH4Gmq
1VvTpz3cS0C9O3NsgcI1cQqoV9pH1/1FypAlXXPg+guccaJeAh94P9F/yqpFYOqb
S2nZ8nww7Ieos/BEDezfuTk1wFgDrGJIElJ7dxObu6mSX8AkM2aeu6s57v9AOQip
7wCDRWIPwalSGbUZbh241F9ftppI5vJAGxOEG5EslkEMXxaiwV5lY6bwui9X3STV
V6DdpYslBa0NRDa8ggzGj4hI9+r9Zz4+10wMGd7r0Lxzfrd/jWxkOapIYN81MBmS
SqhPf6CFt6iF0qRARPH9IHrMwdpFnJH1ih+LxO39uNFwZuqpgyLMDw6p7ZrYv9ei
DLXgY9NGuhWBLTOokx5HIHPmvfmDfWTJlPGwo+P3PaIKKcuNhwsLoUnaKJxJGIhM
QkXXRUTgo7UAee9/oUk3p1Z1n1vsrFYx5jCsDf5n+ipSiCUNE+sxwNLZU1t1/XiX
BXJOFd4TKEwcKFkn4cu4ishPsgIZZ8flEbVy6Mf2dVD2kd7T2ud6Lsiznb1IU7YH
QN36brncBnDxp928B8J2xFDqI1MYHfb+KKf3EVwn3lzCIzytIfe6/vTZYaOAjXhJ
1RKApFzolOEWDv/MVXY80YmUz+ua4Bfez+RrTLFQGuIm2tjk0x295Pt6lqN32QZf
Np3D/pr5Xs8M5ogB3lTwQcte5aaYM0vmIdY7hMzPnYPCkmpSrGsImcm+w6PO+Rxp
GFWYMWT8VIOKOPYI0nYdQGUsNuDq3W01lPyKa14d9QNwgYbqN6yK4Pa2i4RK/SGX
5PeqZ36ZGfa+SoTfvz3wsywmY7u4CqB+Wm8DafueKmcSLd+MwWRCzhhNgNDt/VII
c+ym6jB0UE8CnB6KIuBT0A==
`protect END_PROTECTED
