`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FL8/48Nhy7nYnDBuzcYppDeJh4xA72Avrhk82xv6CNm1US0fQTzIPh5b8oZCtqHz
GyB0Zmy5rFUaXA2flPTPgf5qbFR1kAAf+TCxi/8H6igV2uvFxKqzm0oBbR/UNMut
8BjmWFPPBLlNUNlxByu84EqTi98NWF1vft9DUK/E04AEy6pJRKP/C0Iay4YknhYx
0jv+vE7AN8Aql0dG3LFUqcaSAR5x4/zRz676wJ2BnZFXkMuTI6UZuR8+mC9mYtHb
Nxqud2USopjJdagFoAOJwz+KIFOAS3TZzTI9+/uVo7OvnjHCQgFagYaHEwlORfJx
10/C7Ze816wBlBJ0fqoeEKpvpwIhmEZIy8F9R7VePKHpdG9r6AfGW/0SMg6FOqPy
UFtjqCJmDiEYhbMRWw6NSmB61H4CqjNHYKaeTu1G303PlpF6oN90APJFLkHQDR98
5thy7cbykdbv2zLrmDk5Zg1va5CuKGsPvfuBM2vVT7sp3cbC4SZSBZ7y75iRn4il
GUs3j2gs/wjLKWuWAc8baz0gxt2Q+rHYUY3ASSSn16njbkvJ895Ed8zfTUt7FiPm
mHgVS91lmJ2oXQOlgYSEyEFey/Ie4SKkg3Uv2vtkVVbjrmlYaVNNBYgIPqHWnbPy
wd8Zv9st0TzwE8BuGRRG102DBEDrxgLfQt8sk9RkB9tecjwi9fcU4KuY0NZ1Q2Vg
pOZlt+zRLYW+FB/840FyWSuMrnMnnZim9ef1eCAFspPQNuEUkroFJYA2cM/AHlHH
CputrtJrPvm5pAVSI8GEtl+RGo7UNWkl20hgwUT2/8Pzm623OIpMuVejq2r2Qc1h
S3Tog0opnuhVckqTtcbzWuSLTkra0oSW2JK+lhwUbk7hq4dfjiWN5HSQYx4Y5wdS
xIdaTdyedDGT1jqv7NwSkuKYAUOX0u5LxXA+qXATig9ZGKPzDywty8/N8e7KkpN+
wYAPNXAqgXXjon4OScTbQKuS0Gh/bBACtj7XUy9+oGbSNBi5oYPLx+89oXNqV3DV
xrQf+XWjoWclUIrft+XF9K4WQ6IdJeSsOvHLNP4+i1E5qYY2/UAt/FgRCFAOmlgP
Sc/AhbQuIZJ6i01Kb3BIh3o0ag87JxACEv3E3aMwgsq26aCZcY5axO5bxmeT9Tm9
v42UOapPgABmnyMPEqJOEw==
`protect END_PROTECTED
