`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PRBmHrPefgYQZzn8lLHZybNSA3zM9yhlErHLYGPf4hxGWJmKQ7ZvsiIjZHQlmi6o
6KXuWpB2pQqgsGPl0/XMgA1t6MYT8iOilfHH5D15S5G5qUpCR97eICtwZG0diuAs
+Kl7MGNKLNeiRMuYWsxM28TJClP7CBB4wMe9tnCoBT8icUJYDlhMekTM6Jn7rwG7
2TWwwfRqxHsReLVlt/hN7DZqpD7tQLDFKnlhVDxWxAUPocmWPK2NYT0irRiHUf7y
i+5tkoPaqHTibGhRq0cxSgaxBvl4R3+h6WCcBqWn5AEfE5YraqRFfHk1Me/DruA3
mDuDu/ZeJ4zHRv8OwYUk1RGFrz4/YA1yxpPw/45UuQz2N4x593US3HMdtwg4H5xE
qW1FqvVLH6r2Tpf8HtBmQHNCJzxJUfy6pONhstDH0yr2lW6QkQ370MRICk1czsvI
M92wqt6lt/yAAaSujY1ma/QuTLc267uaGQGYQDQqB4zkTPdhZUmq9zV3X0dIhU5n
BwoZDadLJ3KS3nLoLVR8coJzGbtaapURwAc+gXopu2Abq8AmxMOP5dnVWEwLjAJI
NY0EDTsHVCN1t3w7k/OvBgHenoWOaHTMroDR+kRb0f/5a0P/3MECjVhRr8kuwQpM
2RacZUtRPdtCejFLel2XDViHvrIM3IZs4mPHlScSttckRiChBvbjvhGla9N4gEwk
c6OzaKasy2KNv9/k7AJPW9CVtN0KhI5sKn+KFfEUZTrBo1F6gjrLx6uJBFi0SJGn
UhPOauKUH2TO4Vwqa0Iz6CCuFiXW+Gn2xc49GoDudYHHUU6mKVTl23bJSgSboAV4
2/CSOqV1n3pSViG8XEd1PEWO6aWXB4L9o8kz/YNVGQ88i11veVzr+OU7RFUWAfdo
uvGd1L8+pY0z9T3HgrW8HTkfd6Cq3qLEjnksX8N1lXz7Gbf3FCV6ZATEhIWFIjF/
nKh25zVOs7U/dSXP9nDHt5MjGw39WJeNLVZlKK9K/QrrrbeOwO9YwJhXKd8VJEge
+0KSU1Zpsk0ZqbLCd2EUBwXBQEZFcWbEuW2XeENcAeX1UwGaSKF9dGK7DlU4nFGr
nBj/67n8s0Wtj4hUmu7cHff8JIAlzBUgupeOE/GkrAPGtMlDRgKnzbzeqg479Mlm
bRmOPT+/AkYAmAEBPXqranG7CT/59O01uARiYPCeKRC1uWVcQONuK1NfZletKVBr
iH8J7dW2yNN8l7GQO6RHhZpY/ogR2H+LiwoPhBUD8YWYzUJTQ8ZkrvAqWcoO37Ha
ppSSQYNJCW5EtoNeYdMRmF47GIuahr5/zQ3Z3xaIpVeQguYrijSWggMMxtFnjjUy
3qB8ZjpqbmRrOz3VNHKNHwQdSVDUoegb9Izp7QUDkRWjdHE1MSs451lWgMY3b591
NZRSBhWwRH/94F/CeqbDsGK/yg5ZfsbT0DKsBvNA8Y8ZrsblQ9biCqbaV8bwdD1Z
BDaILJyUYM0W5P82U4ysXIltng2vtRIqdrRryauD+UFmbzas+Y2sVO3bX4J4s1kC
5IRhVQldicBuxSawhb34DUJGgBUdhamYziXiBpnJeU24FQnZtFYB2SYh7yPt5KmF
LNxTHNOSwl6EaE2mFCLoIAwQSGt2ui3ew3Gv+sXvVaFjawpzzu1tdYOD9NGU78pV
Tz/6zO2mzfPxV6s/IFGXu7XUk1v9q3tJhfZ/Oed7wrg5U1tABaIfkcK5USerCc65
GdQG9sV/3poZPrVxD4ijACqouX7g/BXtE1TXLpMXUzrEDNiHFXKnnKMgEev2EIG/
2WDd98WsjVKapAwFZ5Uahn+FdCjCmwbmT3FMqimkyZfW8sSvUuCRb9It9fVAIwbg
WjYvoLRDILA+ClMTrspRBn9UnsOdzGg2yyyye+Z9I8CoRjpiT3xWZr/NWMvM/FOY
IfEIh6t46jq7l3DExULU6Rhe7j04F9c5R7j9OyGmuF2zCiHRcnhmkngNGBGRzrN+
obfqZH76og8Zler1lQ20kweQ7gQTaN8DmQgIxkY9cwREjYPjlRXtU4uAEKwQHz8j
S1tR38kLhWA6xocJGE/ny7R1Wq5TB+tG+85DaqujcE4AOVDFoSd+BtVR5Lv8uyH0
uhT/Wu3hPuLmFpgiDM5VP8snEkYKQJfu9C4OgHE1PSRuLkbuaxzhXIpTH6gfRbE8
392TpZfvLHWge1N8V/PppxnOAPXqMH92/h6opWw+EupyVO+5IlX2ho8ldUpWkkLc
vVdT2oKrrpMTe0LkfHoMgTPEC/5AzksoPDSOPrjIWBJd/P3kmRLexrQDb8/EIgY5
oSUVptwKdM/Ow2L21rvZiMB03R/47njfowWHdH7ZxdyYHIiAGtE0D+ThF+3UtNhE
UWU3qM0mg0N76QmxDMGmHIBJhLWvX84Hlp0TnmX+k/zQrIFMeOCuA5873BWiHTfx
EKBQxZYhiwujZ8NSL7/cywdJMxDdihlF59CgJNakzXbi7Y7zDI4KMtFn80u0pxMQ
O3s+ziFa6rfZUQqObFOPayL0CIwIvLLHmXsG5vnJtZb1VgEjAhn/7GMj06LzCXFy
vMJXMNCv28UrjWKy2Cv9blcO7uISHm7CFEBUn9gysJG2gIaBnvVaZgYmD2mINXsB
uWPtXeh3x+0oUd2AlAUyzi97lumpTj1sPTSZZ8mfuV3uonq2tmq+CzChuYv46JzH
FW4S36xSrVisU1ph5rJzJ3c/P9hn/c4vw9TNunJRuUy+TFf35q8qRLDJnB73xYDk
lEeX5TTCgesx56+iYrE5YyGZAfEbcM0IDU5O93g5WdRO5HQmTVYhqCt4lHT0rgRH
uGocwN3vAOus/vpi/+jPiN9AIdnrLvlA8o6alIG1R6ySN2AqYfe08peFXD4mHoCM
qDnraxOvG1ux5HsAFhcXzgOYaT/P5JtMIsSSWJsbdl8IutBo0AVcXlFoLmfXGmtx
EQuzo5l+DpQ+iOJTIUmdgRpcClf3RfWpGNTZ1XEOlybFYDDgmV9lZrEHcy3wZaps
4mArg8p860Es+Crj+W5gbGSJL62sLOKarDzCIv74685NFn7eL6DVnycH24UQvV0w
0dEzxeGljs/B5lMY6AQq9PVmxuQkkYt4YF6+VwVNHmZNPWy50GFOjxg/R77G1UGh
XvTItbPec+3p4wtPryRwWnBvqCzWtGps8+/BOEYp15lKz/Sv1nlp2j/MFsD66ORk
rbwHlFKJT8iy64YyMzxenGRJ+TV0daZ49HyJBaae1SmfDQSI4FEO8D02vudFmPZE
f1DMbrX9DfTcbYjC9oFDhOLwca1mIBIKIYzzt6aGhiI6pEwTnz2iNzXKceE5Sjtq
CUs04FlKcUx2kN8Xto7kFMzUldDhCQXetDGTnZRRz8pg3KaxhinRaXohoA+ilIuJ
x4Z4SjrIWdlYGPxkj3izadUZvM5FHK1ZP6QVeR8TncIqZcm6WStrvLQPP5pbV9AA
GJNaV5Tg9a827sQ3ZgNTQZ1bfEEBh4pWKvhdZd2PEtNDIDvrNARLpLCz3+8Mg6E8
IYirgm8llq1dEeci3ISy0zijPdlpnVnRT185FIh9J2z5COzqNBGgvwNTBRngWP/d
ze0zTsN1exGeQC9QG4yJ14BaHpSbPbbRw3HnxjX2FJasuMExCbBIBQ7DEg2dLIhS
vkEzuttcHpMLnTb5KShojZ4/pOzHwm/jGaF/O8dgI4NBijkU/LnvAuLi27ZjkTYu
LmMtDLlV/cwDEDl1V7wMxwL/N/NhgLEo4ZW2n4+4+oohCY5Vj2OwU5wIK7tSTmyq
lXCqzInRvDYh0+oFPXGTsCMJmSYd+DC8uOAr19vjZi3b/5y0fIqnYip9QPpeVeO7
l1Oun99X0Zohqh8O36F58DOMAjyAq/0Fzx5cgSjOlQ9HQTfd9ObFbAypQR/orHjp
eBNnuRVQeucsnF+E8gDi+5xQZHz0NdJp3RcCnLv/FpavsILMGTBuEJi+Q6Z1OONH
2nNtSX45mNf0mZA4CypHbJQt6haEzCFa7UflmzSXidnwyLT3j/4JnJ8htz0x2Qif
5UsKzx0L7fEfZaEFfuc+vpl/KvKJQ9y40uPPL5B4bwrvYoP7kJF5ygiDd53sKMaH
v5F2U524P1l+93KzoCJp4VUbriLaxzL5B8PWQdjS/T3H4jOgG0I+7tmvulgt64KT
rrrNKkSkNsbmFlWbDFhs6v1w/TflxyyJIoD9yat6xwAnJ0zTor6khK78atKUUedD
IpsqEuQ0ng9fV1yJ1IQFgL2BERRELIhVduv+kuiXRY4pLBLmP5VWh/YHlZI0eSoK
vj8HOZpWgllWmRETNd4dS9mkQ04XQJdTrhthCrHmy77u5JiHF+x9y37I3e+0WTaP
lozm/XSyzir5mfhEfTp5J/wB7txtyj2fz1LGDBZkfGwn8YcAmqgCbYwhAtBvAA8Q
BvaUTVNZlIiS8OgPFZ9DaT6nRYuEAEKo72AkGJG4okQrKU4SqcaEFIUSM9hGEDU+
hkVsB1+P43h4TgDC1OMIsIauMNBtb9w5DUdnke/gt40p58hMbgyKDhRcYuvMKPZe
w2ABLbyrxU6RfBG9/WXYIYQG+OwWy1YvWY5XpHMzTlr+AsUIk5rkGF63qvSvWaZP
B5SqEWQa+uAtSowknE5CXpT3Q66veuUdQg43EzX4fkkc7ydhibuip4B5TBx4ERc3
MqTW/eJP42w4etOEHQdloEW52yYGxgZ1gnmyT4DeinIEKFZElvCAWWLrHnz3xHe9
PLdNsIifBhTVBjd4a9n+0nZpI0XpdFchVVHGIFyGox5FWTcEB5suzQJ3B3Ecn4Cy
yvTveJgtdKCSVyjAGcU+sQKi/GNr6NfKSDFrB+kROpAS2ciPTa5YFn9ljZgf5k0H
KDtXi8j4DfEWgqzmqXPArQf7CZ5MX78/BYQ2asg+PO1rhNG0YWgiS9PaY4Uq/BuG
OLQPkShH8eKqNpJMgn0JFt5JREtMLGYY+JyIBR0oKNrzP9Vupcc1wBglqtlS9QcC
62XcQqO7yL/xE87oBu9ahhpAzSNVsTjQTQrp9HoPVwCjNmz4PewkAEvoX1iKokJN
gCgVxY5qnItpqYWDN2xcZjP7YzYbjswRKz0E9FkEN5ho5GVrUpgw3fzh5MRf8mu8
HIfY1/2yDq3wp9AZ/oTV9ee2Q6y2Fgjfd2GUi6bDNu444oWvDPNDEskSf4YWxcEU
F3DSAq/ZoBdhZDLx/1Ch77jSSkZTeKvGnVJjT2/Q1utHJ46CgqGvkYg7oHAtGSNd
FMlqCu6PxAGZyOSnPVO16vJhFaDQvjsWnH59U6H1BcOsHS3ZEv/BlMzCLoRBVVWg
GKBnHojqFE3KXr38XRnJpTNSajfxtP8XHwrd7wzmI3/CiEAnvL84JWxL6yHF8QN4
/9ZJPLSaaam8H7qRktiyxYj5xp4QmJqblfdQhQVP8jeHzgFg+y7T/YPmqDzy0p7I
lsfG3nmYeQiRjyRRF7nt2FiIQPo7zEUj/BfKA5BJjaCqVhBC2nuLj6dDmWkjUMeg
iH2BR8Xa/vksxjq06mesivPmmLLi0t6VAPX7sVovX8zVnoGGnH8QwZZejhlIduXM
3xvNXStgvQ8iqFHnhn8TkuNlo/yAvz7PgvWtkb7WiTU9Ig/B0ril4vj0gQ9IlYuZ
87NfXJVgCKvc+cpAAukxXy9uahpv9+Y0acvrWrh6p4rbXJoIf2idyZ5auKyyRQ/c
BOq5kivJt58JV/4EBTGyT1yF0kdr6ySBkLqThX95BYKBeLwVZdwGPPAqbcBVUq0R
L8K26fI1AMdEp4458efbeG5IqZ67bswEtWrXassgTdcxzDmEMcJ7cqL1Z1aGY+lH
Rsdo0uYEIfDCwX1uGQXLOFiWigQ7gFHERvyGdgD6ViN7Mb/GrYxRPtBxzVWDBucV
Of42SfcXd3nHyXqQRQ3sC7GxGqiVCZrOdOG0UX4f8KRuX17LiRAVkVAle5YNrhZG
Vu+N7HKCjCW13+SGGvHPIvKFBxc+WlN6iFazfdwtO3aD1wHGh6rCVetq2ZCIEmHT
A04FaGG06iKwLVpIQex2o043hYmfaf1uFBTjnGcHR0WETd1DuEeqwwbory25tObo
VT4qT6pf2py20akAyr/3SSwz9B116mazeBg56Tq0nKQ1JDNbvT3TjLUwngnnojA2
Nyz9nHfKnjGBSWMA0Qa2/aQt+dg2kV9d/v9vOx3EYK7W6Al589oCyrDnbpW7wVRk
BUZKbXA5x9dgUE1v3FFEHAqq6SwzkhcfVVjgH6siTrNXrgezlCnNxUG7qRLnff7h
ZdPl8kwlZhNxrTFTS5sUFwtWZs7bTLXPP58HAVuGBbqPdakGL1yee5N1+vlFoovS
nkob67pzYK9Uv37McM4yOCHchnUcUQfXU4mw/3WDYXKd5RoW2Hp1JXs6kjSbQhkE
kzlnVGPmB/D7XumKmTH2DP1PnFF6IROLLZPH/SI4xDnreYvThaKeqYe3BmP6PDpO
O/wR/X8cOoCQ5OpVJr395a52uQ8/xgnfeifVwyaNmAVuGIHoYXwDJNLEVa5/FFiq
F+NgMM6LpVIGn/6scszHPlF7Eqwp5xtfhEnbtwa0ngecBfO38ZOdOjXwp61lxG1x
Lxu9u9B4zMlGfVBowPgR3TtmzJYkBh8Fwq8qlPVrRHOyCwuUY/lTvVvOI2JzKIuX
KjCZbY2vP6bqfZ6bM8oGpBkuqBm3EaLLXmPlr2AmT/z9nMAJ6zpCXKvg+DRlWcK4
DR1TPZ1rYqiBiqAMBGDk4vxAT5SrUg8ZCRXPUI4fwrZnPYoA1V1ZLRu7Hc98MySy
8gpJJ97dvQWCucLU5Fr0DmYDnzpJPJJbqrF1asUuIGI+L0AJbwxKsr1juHvbDlGs
pVVZ4h6WzYGVvyvoLpsMbI6KYmVey4XkgHqRWHgbDfTsiS7PgaoYnsVkO0k2Zh2j
2wyXv5ewfdpebIfZoElSrlIntWotIf056XwcAN4AcNEW7Wigx3D02UacP/mHw5TM
YFpcy/UjIghkCfrSEwdwIhsyCLRu0xeYlrHZHB4Exe46PXBCEgRGfxK8rOeFOaum
cEhggxGac1Ya9lClp1nRFL5aV0t/7LdQ+KmMB3yqC1WFfuj9n30NLHNdWUlhwtYX
UFrNNLMVMAeVouYC6pM2/LBWJ7s3kyqPMeETka9TxkwzJN2WlSI8l4dk06MndhRj
M0GeZOTLIANRfcHzMEPVq58iwYL92LVkp0lJzO0dvP0U5rtxpgK9CaL9CN/6LwXv
GoqRtZn1HzrI9c9qTITmLdF4N9LcbFf7cOwCHMh8MfIccd4m242JjQos1k2Evy6W
zAI0elVTkhEEoaV/MhzGZ3pMiPyHlj2Op40zkPl0raevlz0bjggfAa0a4s+Ki5Vm
6rQZp9x8Mw5eoSBzwjWfbb6FO3IvAKGiWlcTb4MZ+LVIw2NWmxQu6hm3GrJy9NQr
BZ3Jze4bcKP6nKOTtdwvZqR77raplsuLAz4AQDwV1pXN7Co9FZ3xH9JnG5+tYZsP
r5/T7CXhAZuyFv3uvoX3tCH8X74jNEWHQvUZMbTmPdAMsuh2HR89RSKebi24CQZD
fJuh1X0wAOAIV9/Z1QcwUs9lVM0YQwXuKDr4h1t9ob/P5ToSAnbM0snyz3I2W4Od
PUSs5eNS081TAFRInSWrCGSD0UHDBOIe86pkfNWJ6v8kKENrV0FaPKXhNREEfqgy
SsiKKzdZ4HjBUUjJJZyVhj2pQTgE6sjBUUy86sM240Rm1oDIx+2cN0tcNOXlgm/y
Zv96+Rp/vW7ZLdlsUT+wmC8CZYkl7U98VXnNf46KcMk=
`protect END_PROTECTED
