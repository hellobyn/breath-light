`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1dgnrUOtWxuFBwbQbMtsyHl4nKPFHZMQCJNZx1zi/XduDifDUgGC5LfoHurnhhX
9kxhRzf1Vo8Q7wyPyAcR7UioXLO9oFoLjm6J4imGPpCuDryJR3H4ni0U71Jqcq8i
OgxHylzDoFdo54no/gvtM2RgJSK7Oy/AFLuBc8EVrBlNjP9XsBChDhC5+94Ii7V7
PJ7+dZ1qF5CZzoPcNBDtNb1JxV+0Cp0iwacVweoCu4WTJWhvOZWGIjDOeYFchoUL
QV6OSouiuoAL7DVNzdOD9oOGJBjkG8yG77eshB7dK/OwRczsshP+KqcpnJP0WMF1
usg3vkEh4CjHv/JcgWeBB915Xp1J7LE2jvH7V1WkcFjADzxXnwwXyo6LttN5aTLd
OD/LdqEoXOZblNEukjjCPUTKlDLPWM+Vp2OYDFDI0egUrar+U2lAyJQbsCfOVC/F
aFSC6Gdor5bcME7ktsPkZgLo9lz8u5aZCknOIOv0jaIS34f/Ekni4foU6ZbtHlyK
RP+D5TsBm8gEnTmX5f7WaAjBTa05vHXWwd7d2LyoOgWgvmgLzgrDiW3B84okD3zV
ZNC9H7C7UusRyMSWTsKBIfObSG2DipO7v/268GfBI67E06Oj7AS6ijEjy6G0rsls
mvp9nvq/urc4uO1Oky87qWA/GPjtIFCRcxJ7VIKoLRxooU3D9r1CglwtFvQOC+6s
dubbQWzGlAo6EiMpQsiQOGDB0k2glrAiI5viVEiVhAwMC6IPThcNw+IQ3WoA7wCh
G8xWQAx+qksS+aGIV8F3KORwLGr31tCQ2SQE4B1LoLnLAYURYPjxrbnmWieLTc+T
zIJTrgVS75FT/jIQAJAwsx9CNAy+1xkP1uPvnkbIR6iI3/BcZ2v6fyDuru8zp/rb
k9kuB2aEfzR/NpxS5+mpvz01EDACxwgFjAQS1KclZl5/V+/YyTQmwaSNBz7quGew
sq7vGtfPyoH4GJnIPBtX8WqV7jICOTqUr/QWxvh2h6VuUy2wwQtsMdPjeXJ1Kn3G
VbO7fKWISNhWAczP/UCCZN9vTuj1GRAX4zEZpBc1rPA7681Y3fUFefQCOfuFBJ7o
2jazJJvWprQY0y2RSOyR6KUqywPXJzoMDnJ94lMCmnUL/djD45rEqxcT30HKg4xD
SUqoD0Ux+9mGoNamJH06KsoHzduXcgb+kgYqahKW7qI3wFTL/TSFj/GynxReDF8I
ggRjkTVudmiy7S9mlGPIJz6r4ZIumjJscYnUdZi4MeeVrLCdx2ccLBV2K4VGLOxQ
zbuWxD5l2ZMnl24cZGCJuL6Q+s5mUjc7A91mvw5n+YJijYQcHy8oHdLf9ME0LC4/
XBPavjgT2525JqX6SPN7GtltlRih5d6TdIy56bvro82HwtA8ELCvG2yDojOh8SlD
H7vtDS704uCE4/g/aiyXIbXe3YUz+u4uZry7iy+H4n+Zea/a1GC92RWY+q9cjKKe
B936rMLFKGNSuDaHjG2inkL5W+DBGO9+tOxi2+up1JMlqckZGJXc6PSXe86kF7WF
6Yl93ufDAu6maO43ho7KctpisZ3NUdrs81NSE07pwP8pzzWxFQDvfuGPk0FbTrZn
9TXvkByIhUu6Tr1ZrSnWf6ZQK2lrOD4Ng8afxpE8dIRR6neAbnbqActtu6Mgtioz
KkUQDS/VwUz+zWsF6jlkxyYWPw9ISsIdGPYY31ZeoklYc7oXnF5VXOOt/MxpdCQO
K+sQjtHa6uOz+vFm6ypID1wRLe8sQxX5FcWCqSlCXkLPJZDiCDpbZ2yiMvfLA0L5
z2+Joj9BDOZDAiaIKFk4lH6kWtfJdt4XX7sV61YJhSSeTOyNaFTj/KO52xWoSWa4
gGHqSqNd9SbBUiH5B3/nWvm9hi/X1VIaff4p2cwv92Fu0wouLoBLUp5XfzAyPfWl
EYQko3z7SpUn7aRYS4vCmDGUr2yjsShrtFqnTLvK+SHzPsxD5+1yac4IUrGFz6AR
1ypyJzgng6PhedQkjZRkkxA3MajnpcpKe+l+RLbN0pc7q2zSNWhANu7kj+hynZ3B
pq69meLhNA/dp2+953lipoandoBIySHh8zy5GhgLhH4xiMuNsQd549rEWl1/c8o3
LnVCegKB/MyoejRUC1i5p3BiaFC51TTTpjKkp1pJAmUq5jjCQjoPLlHF6D+ba0lV
d0Ty7i01jWJRiSO5Z6es5DSliaa81dk3nO9T0y/gDtjqyVnhrs+DL6QEns9g7n2B
t8dNqM0UX/6lNVEEBF9S0qqzSt41hCXus5OdzpKqBZrh9n47vuV1dFnrWvWvarOy
zk4dNL/HnEqkS7DhcIp3lGwPRiaJfG8QIW9yyYFljQAnJwDQAti9aq54rFS93hn+
HiMiX3RY2PapPDWMHuWDCWEFA/RiCz3RQmuWOIfCAU67n0qg/yTycyfrSJVQkTRp
14h8m5cwT+YojSpSOSjMk1NX90uWZJqoRpW053MCWxK3W52yDf4pLU5kRhWYs5Rp
/l7yzxTJ93PnHHGL/S0Hlecj6IOUW8tfYV6UX24KCoYnaG2K8kCdYbUCs7s1E8XP
bbf+UmUVWIoBW+NygKjiLeqSC6+uOBtZEuYruBisH6fSpLWwsw0vkMsbLnWySLRl
XSrbb/lmhqcxp2qBk3EfHmrmz4d8ripUgYzPGp1R6bkhnsRIFTuiSgJKXlsc8oKw
koa2O8yPLhkztmn08Ep1uPEWRNo2LjEZ5oiPF7YBmG7XbSnzsI3QwITKUcLg5Yze
Zdf2Ec8hu8p2liscntLdtrZVznoeJMmfrZvjbnXXsW+P3O4pzf0MTiHZrApGBX95
zffP3S2laQklzOucAahLcHWj/kltE5cWK2GvMwCQ9tDw4fta73JH5HXCYXRMoiAW
gl/G9dYOyDRTwI0IIEJE08NlzxNpOfoM9z7KtQRgmgc/B3yYWOC9YzitzKrJHBmo
xsbdooKQeMY7yo8EoDweqX4+Ie0D350W1dflSlv+2PM76OA2eUhtcA7Vw/eo1+D9
wSQ7GuELAjw/G6hM003XrolwwMcu3j8Sh46CYL0MgKIQ46deUdLWCJtDWpcxiu/c
AqzvCtUwP/t1xyXBR+KUIV3EZe5QuamS7vByR1fozos1Dk6+bYeN8X1TgLfXrFwY
DIMcacGubnE2Y0RfVywWxmGsEGb+8WmJjxpAYGZX2Xep9K1nb9MEGFwbV4S4/XRo
UT/tuVZ5dRIguo/Lvf/ROxCKXF9/VLIzfH6zmhVwPWsiVUIuLnhYBGaElV/SwS3I
7n6+fOyJWzFpyedpDHaSfV7spT3vVLDMIGxh3wuwgVh7a0SVUK69NDUZjBe6S6El
U9yCfQ0OG45+/WBttpKYaanKNDAFHqeJ4US3Mu9NhWZDGrC04N4wvqtscBdMdwRt
ljYIUZR1zLeey+0RkEH0t1yRLqtvYFfttjcsigAy3R95jB0vJvrdzryj6wPey3Bm
xJdg2XEiuNJKBDRPJHa6ENo7T3/Y1Hsl/JKhswD7tB2LfiuZDxwkYOMqMqWYKqFR
YLPtu2MGO+p2FK4gad4XaFGcwVVsiOa8EP72NObrflfGvXUJy1CwDkcbjS/uLCz2
a186Sb6/NXwxenqqQbOr8qL31q2m1QHKTjJ0IAapceZB2Np/qe5d9ZWIvePuzdm/
GWYMZBHPF+hmfBw0JsoPZz44OBmoh3ulHnnquCrmOoDDGWqQi6yKGzapWCQKnv6v
LvCrmU5eGhh0S4FA6tRawey3VijOrHnWgaK6Y5PUiQ7NwBORwFBI1awGpLLR9Qh8
BB4sagdrVVdNgLiX05sb4YMQlBx4NOgameIj8eYvn4ptxRJ0bCr5467EIijNLdOX
kRvbc5K0u0nYI4gcA/tO3KaejwxEtv6IB17LBL1r2c44OTPZk2pujFBdwGIw8bnn
Ty55YZlhCKfNNapmkHpSEVVOEkWcMXyXGNQaibSfkx66up1yNzs1WUpcTRtvO4N5
M7dBwfEsxqp30nANwOZ1LC0q2C3Uo2tAF1oyHkG30JepIvJESfgzm5OUbiqcs0V6
iu6oeSsF4uU9YFjjloto7/inZQSv2hAnZF4i79bP/+MYZyVE+6ZdfQr+Z7QPf/Kd
jFmu+m/ImIMHiBQ8/BjwUQu1mZF1p31XWtau+/+V5WGeV/6guOy3m7lmr40NX9fn
+cC3GcWCw4K2iOjsq+m5OGNS8RLXGgB99Sn1Q/UdGX6h8Voj7VpOAb3IoTK/egDc
qKT/8ttlrdHskOH9E0p4Uh2KQEkK79dsCgNXMRzmXjzAyeRuY4W+KAbe/L26Uin7
eOcRzpAAIEkfi+6/xBhoxcfqlMCg18XW+UMQ668sd9by/o8YEK2fe5gZ9vxrafyW
aD3lVtzvHfbyY09Fx/ScB3k29Y6vAl1q0FEyK717H293NGQikJw8oD+p82fVpYNG
zsAVivX/TS9eDegwOWMCFv9YenCAT19q/1mC3b+RWoaCoTdYKD2IdE7Fd23Ji89K
u3fvP6Y/4j0kmUUr+5WZ8R8aLbhMSL4vUgACsd5tKBuEPW7fZmlHE7PZPQRfAqcH
7tNH226GQ0UxUMtiYuqxXqG9Wr0cfT6yHTdMWv/hJjbkieVFUmVzpFR7kwIY+SAJ
/x2s/adhlppPyTQHa3CWyeZJjyNo3h3EWEsHgR+YV+Ux9GrIqFLZ6PNgOD3qZyBy
TMtIX163e8ywO3kS6OH4HopmJFZvn3MhYhb6dSXXp950Co8mTUy5FpLP4cFCRLep
PjbO+XHsJvCYgQoXf7Y4sUFu7y8swKLI1W2r+vFFnSEBtLnLTzGB3dbSKO5+9KzE
P1UQFgBRnwzu2S1dBLp8beZesdB0JMYeGUpbdXyiTCGN2bT3hdSFoeOCOW5P+HFj
J97yj/6k7IsPdWLtzqcMRo9DmsaZO9gChlV91MrW4/cIYLTLXefAe8LcsK8yntMG
mdjMY1wasea5RHQJdhPgyz5QIJeMhdgpnTq/tMrD4EU3lYIVN2SBsiKTzErBRn+s
XZXBKUCFGTg+cEf8o8aQY/zLVUf+yd7x+dsVUs+tuCnWGH+o6k1bL6qrWxbits9t
fKKV/uF/StoOTkkd8KCIwVZcxEoVfHDgsU1/0VHtxAoZRJN8y4aG0ZOVH4GfB487
nK+9BPy+CLtxjF2BEQZ3yOhQ5CvUZ+/LIeY798BakuBjjOHVg16dgMlH8rHR6fT6
r834VdVIkw5OVnzhQjiujXWxbXyNkYfo4I//4NGAwi23GwrztIYdFNVvNcWxfRgw
jngrhMSO5h/BI8mleV6UqOMCnN38bVyLOrcaZF0FCndoMCAX8JG/wsw/s4Jxhn0e
24O3fXrKQ+IjK4LMvdoqkBPLGN0TXTJh+GgxOrwrt9XANDsw02c8cIWybz0vcLGl
ZEB4lfRp4QlOzzPS/yDHYoQtAY1ozmJg24IEFkb3bnlE9j9tTD0+Pt/6TMgGH+TD
fuKAhc26x3OTYDHANV3yvFdWqDUCbeynQ5NonlHToBQrfF5ieF/OI67Ef2K0P3HY
2rXVKvAj85qs1pqPywxf4sCu00492w7s2pkKmotR19ycSY9QC9+lfGeMr3SPtK1K
DEZ6SFaxkhlSTD+eb+y/Xov/swDbpL1oxbebhjyGCctW6m+HIA3y9mAXpejSDg9Z
uS+2gxdaiHuBMBaaIxG8QtqNX/WAvJ/xLCuMvCP3R60JhJ6wZMhE31l2orkAMTDM
93cal4xBPNwj01IQjM6noCzfDRPFR+XbwjOwON0Q66GeCQQ9wNyf/B3P9bK2iqqv
edi0K+/68zMWLOd8MiCkLti8iFVRstJaEWdgROUEHK+L9E47dsgij6ASrs98SOWn
g99aOgszKDhA1BGRKc1Awb6yFRh+o4N0NzNp9F6n6ym0P5Rx1R6RtfL/7fvtqw0O
fFtbFfG83EDOzUyH3lEv5obfxGlPUrufcIu5yGHp2uFpSo+HrvFqvCgH5X7EHdnX
BG5fES7rpC9irPNtWAiFgWLgdXuHH370hNGeeH9sAnhIOMnvxSF/wlt1zJXyUzmG
WcevxxfiOtB8MJiPDkjttG3BdOnmbsU5zz2z5kVAmdh3xjIV6QBOc56b1t0DwOFw
Htn9GVshhcT1W4jdj4isdq7QDODZHyi4KjwHvkT1vpAEu9JwdmqeUisF2q/e1gY6
CGBdoAuvsI/N8Yc7UkZ7bk5MRVdEbZ3t1ryWLmg2ijGcKHOeIFqwmsR18wZViQNQ
EA+CvA1VNNoPrziLXShNaR5wD7N8TEyUN3H/W5LGaX61BMAdg6OjmMNd5T7Hz75W
o8/v/2r0taewbSTFRxF2Ni846B48A6FHni61bm5QNSWB++5NTfMwEnt81ymibjas
s193vDLhta+XhtnkDKxg8kTtVGzJu+BURxD+R7Kv9n+GB6eT2WVRbfoU+RiLBQjA
wimBjzXcTO5Ih+2nFynp6QIV5/0rP4iDztDSJ36i2qAQ4X4+A4tq49XuWvV+vKFd
EtgnCKzXdPuZseFODW1g2jEbyTky72+ZVtSVcKn4F293hmc6W3Eu2N7jFMt4LyHQ
Sys0Padl5FmEAPT7vLIMQfF7WTWSjm7G6M8WIY6I/0YaghD5Mn4aPnPDnAhRGJPi
afntH50UfE0/32547doytntebmSTyjoERhqU3MWt72jPNjcFeGKNoZ+lLOpUgBae
EJN7iAu5uquJha7bkCR8NEb2/AWsVxU7KTmfT7Mr4JuSMjhrEFByAzqnfBuS2M2C
skx7vbUEtLIf+T2XcEPSYXCxXEJtLlu1Sv4o/8B7TVLnW5xPi8gmUgikUo057YJr
f4G8Ua/SCMJ/EMxk1FigkZOMJnMJfISlgo8Ko1yjwllyKJxa1DIkkH3pCVcIpZ5U
4G8v59IrCsjYSm6NKWK9CmwBIR/aVVaB6EfVSO4EWV8ziIgOpjyxl37WhONTlMub
Fk+3OQ29vlWtI3ieZP7VHcM4XUUBOGjPUVqbazJI74zZPM3sZiXyShCECQVgFMdF
XfKJBuifcLEn42Wk4UXQhMBj/HmKXMDPFVrqLIxvfrk831sjkX0loGaYqJD3PwcY
0D0mm5nnaT6kbhU51eMuT1HEHzGQ/TB5wCygheeX4pH3/xSlV3rLBM/aL6XS+ZuK
qw8haK6Ke9pT2tlQ3osKQffRP3VuLDgQARALsMH/gukz9FWNu/7T1CG6Gw1QnjYG
vvyXzE1segxFEqKYpfZGFubaSHsWx2MRgmvbhKpa8NKnN5JrulWZw5CxpxFyX+53
+kY/0+Aqq8Tt6Mg5ZxoUAuFNALJlv375wJxdaaRlJ15QtK3P55soE7Gy6DLzlk3Q
82ba0/7T+iFDOOKbg/r1V8p8aephQ8XLkkzy55kuy95FCdkRN0KY7yaQYwS/7fXz
U2W1h4uDTrI2ZaO5068Z2KBYcznC0LTWWgvvdO1lhuNAuZ0X1leIph49CnzdO2aA
ijgAivqMtyHkm2KG2/dEVA6bun0dWdCFRll49iWgCcf6dUdP4buPSyF9eJOM6M3R
zfNEjN4JPd2Uitopl0w8yZ/2oMrsObDpx9PQlMaENX/AwtkedL4u6XwLyrjNNlzf
K/ktsX7Sl6BMyfW5Yt2ffGbPvO7L4+QK6zr/IxTraJqXcPHAaeBU8TWiqEVXpm+V
W3yafmkS3TGqnHP8KNmV/4Rs6KXpENYvl6Fvm1NMEHJnJJPth75JIQjBM97S/qeU
/31IVVYx39m5glHJZddZKEBG7lqCZnbI+vV6lpLfQuy6DErJjws5AczkBWJ22bpv
6+EKYL2SYRgPbOqCFT8cVD2peIGt/dz2dNlY6VMe8EPh0To0Igo3To6362VAx8jO
QGp43iNcuYAupUC2iGKWm69FvoDdHL8YNXtJ1U0zCf6+3utJmOODFAK/Tt7AcTW7
Lb8p8wE8WYmYACrB7+Pmd377dC+s/28M0N7D3r3BrnMuZ1kBV/VQvbcgBOAF8akF
pvGKmaGeHEgfq8RLKml9DTBaaOPAXMJw4FJ/ul8oRBHcfISeM7d0cxOsnyWWaldh
ityMojKMlgrnw42GnjyUSYPPuqWn4NLC8TC4kuC0qGu7chwGxFb+Gf7j3gR5UDGS
TChMq5mYQRaeKpV6AkYBNuOa8eaM7qz0TYFLuFuIrVd/Qq8FKdYbNi7aVWBccEz1
UxtUctXENlrZI1ED/FDikd5X4IpvJpMEujJeFSHVOCXCrXRLfeXr6JKtvw1qCKpa
n6u19DtNjsQEBDGjnI7LtZrmvIbLqWBU3tv4ZZUtSM986Tntp4gEfm4vT3J+P9BL
kaSoxXUx2sp+rsxq79oErfFtGHnps0wCtgxw+B7v2CjjrxOFXiwBns2t+1dr7hvi
NTk0GTfeRQ24fiAc+FyYrF+BCJ7qCbodVSWYJp4CbQjFAYFVQ4aldKHPGIfMSrL2
i5w/jbnrNipZbSjLUvO09zcvpxGHKzq/VUSRRIAdWqy9JX0+O57OcbrTVS74tkye
pGlx85M/AxKkAWi+tSbpmEfinmTjSxZgqw3vSO2I80m8YfFkb9g/i75DyuL8phdj
GNTycJ7gnJSbA+BdnjhoIWMa3LQ2xGpDBnNwB3TNAszxt64MepM0gEr5FYesIiEg
heMF+qS9JO24eqneKRDm6zsFVRGd+0syF6DXs9Ekw8RZbWRCtJbuD61ZXKXNJuQ+
KDaUSMW7kXSkjtENHz3BfhiW91p7f8z2niiyND4aZISIlxUUs6RTnBnoSirTHdMh
v5sOik5snf/NnWQD38IRpNfDePQN+/4pF+8tWTOjA1VYY4rhFNCpvHydKruQSJhA
IpkeL/O2d3MRvbwb9N4H06aTb6DrL0bB/ZUb4V2mkrqlCAliGKev9d7AN22lkqXh
bmgHPl31Wa/wfqViTbhrWCHqJDzYnvEmoJ97aXCVTnUpk0BK08BqdVxa8EMQ1zzY
JxITueKLjhTVEc0hZIY1N9Y5Q8OrDKUV1pRqCtSgjrGEwdtTMG7FI4sbnLXYMMQh
b/tDKOEJicL8soIwENS+GuApaC+IRILdoIX+iW8BkbrWuTvFly/MGNrAslmuWpgO
CZpZaBovxIdSMPj+jls3t0PJiXCKFnDX0GiRYvgrZ775p+b8zkBc+hLSXdBqFT0E
NzncLx5RAWSyUeo8Xu18mOYsUkH72tRrrLfepMLoiLJ7DFTT01GWD+ot8j6q+I0w
xjSkHA8vN4lUG/y2Ybi5Fnl5S37JCeZB8u1K9dt7FNz3knoxOkvGOy5w5bJKptbv
uKXFdskWMkwfMWhsHB9WwDXKN2EwFJQn5/WQaQXGxJGF9d3sB/V3x9RCkoyT6I0M
Vi4aDC+AO8IF13Ro463rBmEkyKfyhrTs8Ka6ZeloNDPt+OSfd9dgZRaqeQ6nLfIU
SqWj6zOs9jIEVBXlQvoVq+S4ZwQHbOm5MFJ1dUkiVtpbKGliZicKHH1walq+5C+a
fpZXruo24YAUwkxFeXzg5xlmUVcNROc46GadGrrv4tSg+B1NtXjz8mti96xYocU0
ABtX10KyZv4mPz1CXYpDOMmPrPVfUnnoLu6sckn3Gh0ppEnZuAvHc+479pSzKj2a
TinzJMfijiC5WEyIWkgRS1WPJcnSsYxVPEQVEx8P7Fmori9cRWgCkeRuabe371Fv
4Dqlu2ija7ul8zocfY8J0LmoS/znqVUAZFVxqzzKk19m1Q+VQo6OYlp6HLnp1jKP
6i/qvUU8Nk0J6n7OiLG22bZMgVPkadtA7Qx9x4bLyI7PooXlb2ooNslb/ke2h4/3
hqzEL/bdBrkBVyxT2hStQM4+PQUHBeyifw6LrIKmbuCJVQoC25C+Qc8tyf+AiqSe
oZrQhpktDGroBZO4WTm9csKBOdVfqZAHiShlK6GsGrcCi6bozRQK9Frnonsoh1Fo
d/Xx28MwQU15O4qIkVEup0xWHMNZKQo7sTvISAw+a3eKKgAyzGqW4TEd5iPO53PZ
VW57MQZTB/Bpp1/tyeM9ZtK28Rs5X2meRsLkvqqsn5hQvAp60TWm+75+RvtNk/OL
9sg4FcMxjJiJKhgpM884AG5oaz3F1QmY5991fGnF9sbxbsSbBpqdjJBe58xN7/sl
WkwHQbEFRnT3404f/n/eqrB9wtiA7SvqoKn1t6BUzz/a0Mrk3oJETVDBF/ZWfNK4
UHTm7sIOuEhHwlcPIWQfWRHRVmrXtgEzZvVDMyl5/jnHGZwlDCgOQqufugtftqid
/1SLaMUon/wC+wgeQ6kivWSs3cW5cu7R74ANkRLX7Mcuakof1qMLTgH9WRW7pKFB
M2hV5kB5SJ8B6oEygsJHJWuKbv3s3cjpZSSsnew+fC0Zt4xV7rNw/fElzTKh3L2a
gVsawv5W0Li1jpwC59+LHQDH+PDHrT9IpQ5q0B8enJwqYdGRF9DCVue4bsdrt/Wa
lxKNZLejdDsoEu496pVj7qXmJcyallnwzbOrO3Gbc1uPLy8Xoca0F43zCKPJStRg
Z1w3dec+3iU75joCHy38zvK9aSSjYl5iz6fXRaAN2hzbF4ri19UrnEItp9eVbpS4
2Ie2P3yrjlE9eFJE5lzWjbJ0j22hmXAWDQuwGjT8riLH4hl9UxWyyPbKIbNA2Ka1
pw03Wtc55FYs7uKQSR8NkyvFBRxo6xcU7hOvoqZS0hfbpobM5WaglMZMwv9PEj5J
6GjEgaP+AjC2KYiEAfcgGjZALmc+/sG8GjradBpW9hqDTEhepPVxuv5bsIfE890d
gI+3f2mug7pTo2EaVpORN+j+rh+/CxmYkVHRCU/1f7f2/rlW6pgqI4hb9x11GhkK
baMjoL5uvnZJZ5KnXy2L3INZ0LUj03etvgTKFKoO9OqUlVhXuvMSZn+TgdLmh7YR
sofBgtTrwGlBgdPJlz961BRzYTxChmhYArBQRr3egJPicyvQ7iNOUNZYkvJEDZk8
RmVF7nuBujMO/heqWIYX9Mb7PsCf+9s8Wri8nJenYRr8LAA1cogD97y28fmN+dAt
i7PM4Y20jo0IZWxTigNujy7YGb/bN+evf+xnAxDYhhBR/Hs1XDXpp4tShvrmQAvx
s8tnXgcwKXy/nWLWN/O1/IHXI6MCc0m9OQQWaPagTrYtBqGg4EsvBtfurewp/5zv
gbSw+lZ+uPTFqaXsmnxs7vRKMHOqTmfA45jCwlEvKzAd9jFwykQ7F0qaAQ068F/F
a/HwCLSQpXT1yP4glqlzdVnRP76dI9iwEZr5PjvzlArUnqrR/DN6AXlAugzBbyl4
w462ULYn4ZkJALR0EcJWbt9mu1oYH1o4D1FgCBKzhlS1Eomc0B2smQ+ayY213vsM
/5ZoPFTyHJDgP68r+x2PqNcB0b2BU4GHh5MSnjIVj5tR3dub5+4Cex0cUXPQk/lz
zSZc/zrQ9FlXj8QYW/KnWgWsM88voW7oCFUjOd5o+6Z+pGSZevh2YI/GLAoOPNbE
/PmtojZsE0RUSljCK58GEah4MhCeXGTLrsEmcwTWBxORN+AGuCfDRhAYjzaFEKtC
X8X0WgvPZXEp+rKGcSCUm43IPDmS5DcG7VPo5rjrA7xsi0KWPvl1rqJko/WGi6kN
YxsE4Q0dBKyKd5wWT5Np42gdt6E9I6zT7l5I7qfnEqx1yj3epbXTRWuheFa6WEMS
Tblf2ygc0LDquQyzd6X6S2z63lBxQPwlctrgcQtnCR5TkGssfePE7R0Cd9rB2ZOb
N5bFRyrKsL+uQFsgp+Hhy/qI/B86YN3HOIWzp6YrdLz47Fki35wcgA9TKqS6pd9l
4bAs0+dzlArHHBbQZaZ0AG7Lvuy9M8PI+4Nxtlo3mr2A1rOPrNEKm2jTnipeJtxY
o2dFRVXJRJMk9rz8StlN+DqGjzG+nkXMYsSG6dGXI5+ztZmQDS04kqacUySn4Ses
AMcBRPQQ7WwTvZ5EFp+9cpHJ8N25sP9JncWt37zeJtFFuOup5zdmQS/2CROghqSz
ZrXWi0qTbrKLPs8LWVDAwcIK3IVM0j+rtTV/J6qCe2SlzBChFqmoPrj/ehn4HLFR
aqEeaMeI7eJR3oR0hs/WXVEWlc/gU3k8pvtv31mSfKS30dwIbjTbmDcbK2hs0ZJd
GqUbc5D5Irr6J/EL5qSBFyPg/EieFUGnLog1DQs06sPN/5ulno63cUaEsH7EbMSe
YsCgdw2b/oYcPHkUPpevyURcI/Uw/IMzYTRxRv74Gl1zVcP8FVR8vtz15s/WLGmO
AhTFBvKacHisqZY/ymVBCQ6yvVyHjpA70O+fiObjIqLdsdzGyCEpjMJh/G+sVFg3
rzy79JMhhcmeQvM0tNGPXXWiE2LrLUhczotgEIDfVW8rzum33X2DK10c0mFZxi/n
XSgNM/RaVoGS3kmZwUJCiMGyeoF2O4ZIFqakTLSJIL5jLpurZJzvKUNt2XyW3Fx3
97Al9DRTGKAtzpNJB/bR8Q3g5DWC2JIUYwhy/PZy0/0f0aU9iFzr+pZdWaHtmIzp
BwPsfZhbudicziI+TjwN1XD548KjiHMB6ZVlZaQwWGXVSjp/UPiI1DlXyX6Hi6cg
ptaY6gyamonBCgu5UXvkaR6FBor7S2SHIteQUoLxPsLfWNVb0nntTzyplOdjdOQQ
JZw3w9GJqV28YWHaGcdFrzsLAk/TRbF4Rdq4C+iEvlgx77bQG8HoZnIFVI3tseqy
pDjGNKpxoBdJZyxXRvleNfRi59odUN4+xCQGpHhZyeuJUUUu8vQMRBCtAcORGXJF
3mMg4Q4AWvAwpn5Oi3/qG1UFNT2RM9TmvtZVMM2mof6kXECpK8Sai1jlrWSv0bSh
SXRgD5h0qBgSSBtxRFYkezes1+LLW1/GxWmQslSw46hDYvDP2iDv5wPPnade+iXT
ktbJQYa1gqG7GeM6HcKxzM/iy7p7VogbBt2F9ZcwUwVRVzIXa7y8CaYwSczCQXln
1zk7J0W3msKxWjwK96tSi3DORscHUU6uZ4eCOUjPd4ey/iexEEnmKEi+ZHTmUpzp
3m8GCB16Dy2QxhTAYzqwFObPSFnLohazceTMJPyITG2TUATJVjq5dJp649+9+k0A
TPOxHOuzRdU1D8MPsoXTQuHj2XPU26hOWhY1JbwMiVsFsVO1q+DIAGna+UvGORsQ
xvKuaYAVIQoL5zk3xtWTye22j4momar+TUq4KpWVysLeMJvBamonbtQ0WzlXDoqm
TuJK++9kz/IlNPi5l3n9ql9kGVBgMR8zRC75dSkGxy/EcSQff/+8hGmKwaZ+HQsP
bR/v/TL41F/20ExWYBd913hQu4yIvRoSu3Zz4NaBWUGrGSvz49phVHuz4cqWBAnl
3gPHWygL82i4VZqWYAWt9o5AKVsueVcwva4M9ooQPK1aNdsIg1q1cr/LO5FCtAJO
Ji908odi/S8d58Jhr6vEH2NQbQPutjPk0ZaBkVlh2UR3Nxto3tFzT6Yr6xqM6aW2
aWtdcNVwQBV0FuIJlNM0Br5ir/W/ewelyCvDt3Gxm/bUulnNhdsiTKUUazZnQ+MZ
nsHLPGUiBvFPdu3F0z3440At8CyC9qKMff/ctB8EW/58C99PwIq8wMSp5RPxkrDE
PMtjs27FX1EKRYrMK3Ur/JxyHpng6+wVi39Kz8WOOupT7vNPG8rCGuXN6O72+aUG
Kmkx9LaHxQTMqbAkEXL/UcqMMxnUAoixrMkZjMkRqM57d1kDzrjnvc2oCNsJjTWg
fos/meALbkkwkoJGTYkSINe6sYSpJbiQxUN/pHlvjtD/6TZKA3HaCtNLXOe13C24
ZHZTylJoiZqOxpQ/JuZ14nJlD711UOof/rGnzc/itmd/32Cx/CUVhuG+U8ajxP21
bzU1Bu2GWXcCJgp2/HAzStIwKAnNFLC741YVWssWLSO9IRqJLgh+WAUk6+IWH00X
ln05hQCQRAglRKm6E3Q55/tTF4YVXqavKjiZ/TaBWqaCLEZuqqZrocM9UJ50jg4l
yZbbqmnuswIZWfEQ60umhRnW+6i6bfzOlqmpglBFk+L/cZ2xhhfUwnlunmls2ZuV
cW+CZpYW1g7w4+808fQ8jwXBlYws8pC8LVhT5EC6x7jNV25PfUgiUAIielHGmYJV
A+2oZgPby5ENyH9QJl021mElZsCV0k25mQYi7HO/QkX7tzY7k4OQMBYVXWixUSVF
gXEBHPAXTH/bGyPPsbAc4fSlt6Rt/amQj9/2+0tCTfrymwz1Vbv1Ngcgy3xqncQ5
UpAorvpH33/VtRQnqJaCRCzZqI3e4l4+tLa11TPpeRLAV4TzDymcqnONT7kjNORc
67EPJ8Q+IFmi0+gODNT1Z+DP4TyN+58tmw02LYye11Ie9HLRhrStjmjRyHVMvR9h
u/evrSrMZIWhPwHcyMU67llSwpKmxEyosO37SGk6HC5dcN4cZDL4+UhlFeV1m7KS
q1S2B0PlmYIlPXRTSeD2MwuswCveRqenFz0jbZvlh3hlJ+IaM8T45LLnZW1yFSdv
4wpwoyq+4A2aWiYUzLw6VOL+kKKfYKiXkFQdB0JVE6ww/HqoYFGtKCC+sJ2ULSTZ
fRN/jK6TuAvsBvtCayvMGbjRPON1kAZgBB+qS2kWJ2UlTQekSmPZMyUpf4h8YvFu
dY3L2cIhDDwLJjvstuwQUyTVH5Ny7kxkieg45mTFMXQ03aAsEhUXoceWJ0rYryhG
YApMN0EfRD2fHoLuRHCRAIVHptQnsBi02USWyvP4eeqxtGSJFzWML09xoThV4iO/
4+LZFriXrfA3L4eNVR6vYnbRNBFyK7li+8Udl78s+9Pjq2py/7s1onjJOmxqYxb9
yKFe7gUWnCYMcf6B0v2VWf/rzyIfYKblc0+xmIL8R7Jz9Q7hIczJcIIxACeRkDpl
XjvFa03vT5wHmj4Ix4bBia9nEaCdQDEA4zUwft5MFxTLv4p3+iRoiR1X1kmSe19M
ivZLEoXqrxDfcZtwBHboKc9UtTlsZafHtJmsGcqjS6VcC+C0qX4cVFISMz8rOp8k
EXwvcjaqfogrRl89psMrRnyjRfgX2lKcsJHsbfJf5SibIYQtasuMrgN8gKM4h3Jw
wVbHAlBrj0hF2PgBZ8DVpPOICiqk8IoZ+A5JlQiHtiLMrsTQteYF9x+CUIziir5k
vk6Xx6WkehGKFKIIBpr5LMe6f4A9GwLICvkV5uNZ7gpFTOGOf4vzpW71s2tRatf0
LHmvbKAo8CMZdTA8oPJZ61WrEu0ItFkVVZ1DwG4qSlpLbBJDHC18MKQqO3u919qU
86Zp+XqPQ0NqUJvDq+nSsKTzJ5W3hdPWhWqSF8J/WbHbL5moHmeo0772r5ZN5uzw
Y65cbR9ulJ/ZTq3gY1e1WqBHj1cg7sufQWkJn1C5PKC/ejF8hyBp2OtCJ5O9Y0nZ
soLmgoK5xIpBsJKJZ/dE8Fy+PdESa374OA9Wec04mJy3joUEp7AvSJ2rQ9WgcOkV
PdARs73U/ttFHwciridypTWJMPB4l4YB9ukFY9cYfsZ19lv/HtQcsR0xl00CRUzE
j59tke/u3MGWAMZ+2GZPuQaeSruuwVS18MYAH5ccN1RzO0kg3VY7/g8aZeIsEBIu
eQpQDpqRsSRnLb/uGDO+1zb5kp24Kx4QPvZ07FwYuVY=
`protect END_PROTECTED
