`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d12TWCBRobeC5g7sKTyKrXaBX8YLOgm2MF9UhzooAatlL4X3sQrKTR5cXcOuolaS
/7XrEepfV2whXorOU+JrzTgJyWINuhVmO7K5nZi3akqBDmP8d+JwUnYfjsceW7FM
f1Z6n1iYoea5emwjWhiSTQnzfjM2ElZa3x4lCE04iS7wpc3JFKPl9IJ8vw0PsVWe
UH6ErfhPFCPAGuG+sZhAKdb10b8pqJnKcUrK1pv7/pl8HrOcpArcxiifnMSXQEki
lq1LH6bO2tqCmJXEHv1S+lPfkxs6kRe4cbPMZd+v3oVLxm8uMmlaVUI4p8jWdzXY
aT8bheI6TuGaOk85Qtc1ClKRSzhXyM+yElSgoykL86R4ei1GoRhq6aktc+cTXCrx
O51HUKBwGMuqwkvTEUScwRblZ4tIAKMxTn0ptfWPq0Q5K3Qo5yLOWlBHsh4zmkAB
BqsrOjFzgsi2pR22pDOPl3DbBwPTtUsxGNwa7I7d0uH1r9SFP/v7Bi4/k6AdIQ6Y
tgGR3K1SWPCbcX7zoUZ1X8FYoHrogo6JJJAh+VbLR/M=
`protect END_PROTECTED
