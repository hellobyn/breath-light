`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJDW03gmeKEHrJRToL+UNqJ/AkZBtJExEz3qn1f4CXirGsg6Ik2IHlE0RnyQ/Jq0
kXAWerC7uA7nmr3RB/7P9vwBlIj0HyH9g+mrHjNTTltItSvsjlT0fRzt6bl2Imug
IXgTdJO4pMLL/9pdMHWcK6D4E849E/FLMuq8Zfz8CQMQ+PiXNCawmxkz2fC0Uieo
m0WzXgy67hBN5+3mmPwBxAmdDDBor8i6kXQdUlaVeXWG3PVAFWiRqokxZecFZoOv
a1JpUhiN83wHMt6voRZs5nvrkKGdBDr/xz1eQa7qWGkoblRtsN0o7Do2aJiZRhE5
25LcXiU6nG9jLs+6gAG9MM+Fx7SlqoS7PlDQCLxnVvQSLBuoCVhLevoRt/6QCJE8
hHgYXzRNdA4X8StqkejCTQ==
`protect END_PROTECTED
