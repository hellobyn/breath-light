`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjWQhOJiQPPZ6pWo1qb43HkC1quAwlxLVansD7ic2M7AgmGcN/3OxBGahTybI8sg
gdCEunruBcQqoUZy8HUKouxdyDSvi+7+PuNlMuc/g9UW90WzbV54O/tD3fvX5aby
aKrGgvJKMo79yhCthwHHf+SZ8AknAs/gDAazvCXDsBqXSoEkF3Kq2OH/8mH9yLtk
4VjaD136RwImyPui2fESaOjI4/DEc1fsFEf1EL7YE5DmN1YpBUBTqnV06H3eHsbO
l3NpkoX6emn2qQMLTnqIeKcvXi6cYE1WMZ7frvATjzDDgQ64dcvKJ0fImzJ/YxH8
xI5XWPVGl6z9pb4HW9zfoswOT6CMUej+tryK92SnFwaHJV4qDnK21+KJMBCxVdss
WfWLArZ+FFeASpdR7ZjNpWN44BZNL430OmidXa8tfBWigK0fIzpEp92of/9VDA6t
ukPJt4J3/f/owGXHL+K1F4MOBC3U5VTe6lMYHhccYgYr/eq/H8zOiIlVbyezCiuf
DOixLixZvS3IXc1kS6E1mVnbM9j49O2ULvfE/lkc2JIyA/LRYPQu0pMWkyHMtKjt
MzEFNY84ZVg/a8sB4Ps/WPatulRdE8YWC8kCScnm0fc2GaL0hA9m3tnMKg0oD44B
dIUBD7ZXdtl9ykYeMS+Qhz5KCy7NzBLQekpS1ct34t62OSRnxauPIlzjAfiYrW23
JlpuGWjNxBYZIJ0Bj95Tkx+zIxTucTmUWwpx2BlVYBxSxi2Go85eZ+7hObJI92U6
RFe1zUJGjxhDMPMweO/BaSKD3jI8D06eGnaFQR6Oy/M/xzSJXo8GQFvqecrlnhRy
OOBiRJzPtZBec42Qj0L7EPW0crqSBZ5z/cuTxjLssbYSC757836PBqe+F9w+t3sK
OWNVeE2fedym41l8+D2ici9upTs4bgfktcBfvU+WDRs/zmihK7L69gno1mjfN2OG
7eQuOdFTJMGqkphB0qfLflPW6CHrBk43uS/V9L3ZOGJScRpLV9aWwIrtD7cG6jm+
nFUL1GPIREAzMH1nBOGRoPZm/kgxxO/bAUlixdWtYUP4BT7mFwBmNmbVR5ENSlV5
+oiQhHMEGhCHNOZfBOgdFFhkWqAKH/cCAtVUmXGHiAg/y5TY+Hfwmw3UoqXRsGyV
pDuXBqhcc8jIDTsTzFmi4Q+5VIKCuW+mxcXmH9PaeKbwxHYvvXzzj9rey0cY93JE
mNoOBjv9x573EfZ3Y0+ObGJ76ZZV4L9uZy9sAO3f5J1mpx2+7nL9yO0F2m+g8CTn
/YvE3K+81edS7Efmkk8h6CVF/RugWC7KI5tgcXDvVOhG5QCAEcKfLlqZ4rpXV8e/
NCMk3slvBKTatj+oc9bJfopAQHN3RZfghPWET+g7o98ZZUDruu7bEZEkInE6Ft5f
wCy3vzqxo8pvY79sVHAta94XIDoDb4Na+kizyQcLqYmkLisi+YNotjQK99InppfI
2aLHQIq0jazSvGAOqqe+BUogoQ73mmTHQDLAjACrxL/UKak1RsUxTK/KIq+PhEwm
EqiZfMc41GEzuT7xMsbHTyr9wUBJ8tr3g1i/7H3teI2jWevLZ/+HuaFkZ2z2j3YF
obYBhVuCaByEXOgbJ4bKYact4+7/7oG6xN4kloIBTn7kvHYrf8NDsRxh+xxP48UT
bx75T21cXaYK6Z74USVsxu2U49ui+B4AuEsRuR31K6xkTUjooepQXrABwdhjrZ/Q
FDo5DvsLJ/3Bo7SqKuGrSCfKL3zxR5EeTE5gNMKqdyjZNQOxKDIvgOkbTrcOqbaQ
4dFT3wwQ2WPw8CtixdCEbypHADjVqeLJP0VVOtWeaum0QGX6LLPpBU4QU+0Bvkcd
DEzTPh+FZFwKIQMUPJoVLLtnP0BxZb0xhTpfS70Om56uuNAKVYzOeYmzHgS6AYzk
ypXIf132xk78XvE/lBERPfuv30VcSiM9C8hMME+ROTnE/ugPwDy1xu2pfiY27LUw
ecmvTZWCxA+G0geCFXi5kcT3Uk83k2xBUVqcdbhT0mw=
`protect END_PROTECTED
