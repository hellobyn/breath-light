`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqYLw7C8LU7xsRTPvCBOPjuXngYO3V8JGsmSiTSzKG6eyhddBr0UjDnoEslrRdlz
lbmgQCUErCWQnUf/ixV0Hgp0ha2RKBu7Au55xC8D1raJ/QdgAijRJpBm9BDRwzCX
CS8DqIZe3VWDimRiArcamB/LwBOz5tYJHUg8fioRbl+BI63I+Mxz+utZNuDUcq/A
CuEzZDgu7jQWp9ctRqjJDU9aQpDJBZ3sJUS+bvnGaQu2vVjKczrfGGgXe6mwn/+A
Xa1YAwR72WdU0axAy5pfuy0RzxiSSRpdXtKkgxyd20PgX6rzglJcYX+WdIaH+Cxg
cg/GpWq57IjvxBCoNJA8/4MeHDgO92uWhgWTy7PLmqooJFt03ezxqS1c3cQ4SuEN
j87pjzUBJtJq/30gF8Q3/mZKtEqRrhCo6i6AoOHWEBPONvfHDzM7ZRJVQ0vIcC4a
uKcn7ikGN6FVVwla9Ater0G8zWFUiqFeuiZNLXgQ/Zz9/qM4mkEBXGzgLUTqL4eK
VR+x9ByqMB9epfP4ufaaTMnOeVoXmK2DPgtPGSN0slG/out1zJkmgIm8WMFhzHM+
9obSDAenU3Ht8yiLp/xUbq+0J5Il6BjRBW9nMVX1wPgcFoQLdMOx3U2IRnQ4a9vx
lq9SyvkgeEPay9243SxrCk2jiPrHPDqEdaf+66z+KV43McpVid4VWvwN8eGsBXsp
tznwJ2NHhsYjjEQ+bWIBDDpAQP4NGigUQzC85/NqCv9OJMtHraT9/exMBj3Z0rDV
7ZmtHYvTgQuVRl8Ytfo4PuigjAekmtZggRMPUjyZmZ+OENOUivkeL7vI7DvfWhSr
pT0lou2hBWaUvvrByJQZyJsWHh+SJU7S3H39He0hzTar0Oqn8zmuhA90GgACPWSm
10AU6HAWZxhVCtN+sEnn+XNNCCjaXLhO8W2cHDQ8PvsQ0OMm6AOuKkax8SZfFESX
LK7WkLDY3fOsGQHyRs5ShJsjLHnWEhhQNj3bjGoJ0yxO9NBjol/ZWlQMrIZzfdOg
Bm4PmzxpMvIjoCXC6p4AjtaSwW/7He9d/mtkUZ3KxA1byRqujKduBj9P/LhXT1LA
RFqkbq7FkTwAK/dhYenQDIu0JODY+MgBSF3YWCZR2zOkW8ZrcTPSClvi/vb7yCf0
+Hnetbbd48LFPgXd8nawkhuaC/JLYxAOZmA8R527a+3dxE20FntYGA8m5CZse7uV
YncFEziXWFyR55AugcID8LlrJFI25J8SYt/3pUC+qcSXUmXL/CCsAbHGjHzg/4pp
LRTqv0EtCnjkALxdvlAUJNcvcaCWoCblkyrd1zq8hoxAn2y81l8cre6MLHQbQEFy
MlDbu/5GxIoXvkpXzisdp196aE3nmlBQ0xAJhK2E3pv5DmX7lGOHdvJAJZm+FrP4
oxZwK+firQerK6GI/1bovohZ2vSKm7r3eLEzdTcbuDes5jVvEpoLM3hHXxNDLj+/
eLQEfxuctAwHFU+Nb/sfer34EfxkEU/cQZNG3b+VuFhZ1h5Otau3AzySOsZATAAJ
0GPQUOGVORrfdlcMDC6GYcBNzb4YuNNjcxhs2WmK5uVAon+kd+ETJkoog8PgnQiM
ffuiquhTr02/c5FWsbA2GooDwmbS84Q4xqDzfVGgUlbL/Sv/7MtIpefzVeXsYSHE
xqBNZBgQqZiHNdPt5oM1N/Fz28ycyAE3kvyH8CDYi/JAPHrXS7xmuJNR6Xl/uDYY
Hfm+T7nsdWlPmbrQxk8Io0RH8a1G1BOSoKm/ZJayqQWzBCMwBjUcGPNoWLhUNUrg
2Z2giTrKKQfF2ijnA+DZiFvjlDC8A4QsL6ht3udPKPib5SYyvpCmRnOCPl1JytGO
hCFUJjd1xOXY92yrWTZj8F+SMRqHh2LNQCsSaSQfKAVGi6qmVonfoKaQeP6F8F1V
+a1lpXuFsW2YNEWgRvGmqqQMvwfbXlrhJ1ZJ4bEKkrzoN8OpbZTy3BCFq03E0u3U
O9hk4iFnrBoeEIpvJ0LzWwEvGm5yq/Iy6x0vE6S9MxH0sc6YlBGcC95I7UQjpOmd
XDh4x1O80KoK6YUaGGIvD82dtdHQJeS977bWb8pukfU3NAIaYq4dg0YAjqctOyIh
oqbLkkDCMrzaHcLkMK95R8eZ0SzRYqqtSnDl489wQIjJpzei5ULUgqa5efURo6PE
TOxeqDU9+HoCIIxjkdhMzb+OrGKUS86fRoDAyLS5eOQ2yjiQPGzsVb15Gh6TqiJf
Hw1GIhGlbs/IbrDTtt8pXtBNhyelBaG1QagfbzgkUDMbBCMrOF9qOvtMiezpL2q3
+95jNHVNQ2yiwrq/xVQj+4qzc8WodiAUBXU0YcG0odRN3LcXOrHFESbAAvhqMVLR
/M9PWGGiEDRsSmZRJ7/nuLxSxf8NRYAFFgnvtysvCBSsQsE+6bx7fuxiELqXNgQl
I8gVBN/Ls5yAaNseUgn+elJeUcW+MWPs1Pe7LRdZN0eaduEF3hg2g+MRw9QEgPgx
p3HwMI0m6AH3bzgyhliCmYE1SgN9GrfNo35I4eRtigqaZqPOCenJlqFPSr8IqR5j
IyDPjhABdW0z3habm8WY/btSK64taIl0XZtCgHkMhq95x5Bz6njhW7wQW7xCsV1/
92rIF8stTWvfxJGO55Hrxzv1qTDWMeXud2gzsCCFY6HFXpW74CuTVl/5o7VaoTGs
Vn1Gm+E5yWzF5BAkNI1lr3hGCD5MyXrEdaO422Gm0mEbuZXo3W8X7Gv/pSC85RAn
zdP56+HsrnCpNG6fGWsGDA7eS/nRcNTSpvmP/1HRMXDC31XMIni99xfueSxv78p1
zKHCRV4jivlseZkKofr5RkJtxWszJVjqCVRrE0xwfGuynHq+4pvabQ+qn/Q9dQfz
kI9Ls+1hPnvucpTOXHRMcjsz5NJCRFFc13Ff6nPFJZ9lBj8Jn9ZsLcAHeleZV7vJ
vZ4XEZzUyWRl7hDW5PjzO6OAM0Z8kIxR2U+LwXbUTz6r5zrF2WopRpBj/izhxwCZ
UyaUtA+PnhgMxalFCkaUyS6VCPX2Xh2RKXpnpAaJQV5Wte3lKbNUO7hBjS3Eo8EY
+JXcff1aggnTMiJelkQmTd1Wi4+GbFFDZxhkCoUqjyVQfUgyvOvXwB0El4Or+RrH
TELJ8xCFs1foKNKkc2ZgDVkTQ8YDTjY6LGTmWKLfSEMYMgYK92rEGKJI7vSfuGC/
S+ELxBOujMokqoUPvpMV/ilcpJ+j9FYKImZ3Wj9dkNbDjX/UMIByPgT6KJtWSmpp
PlrLxlja37lQftsi201/s/Iw7KBiSmFW2RD4DVvtU7Tx19X/PfhRg+YR9sHiurJj
3uIaXQqEbfVP3Z6yllp+DZk/eUMyq4DODb9HjTnybwcjLBtHU8A1vW1ooOBfSAyT
t+W4FQwugpZy4wD56pGmFIZWfKpmmrmtQqK+rKfMhkIFj/7kCjucWUxzqoWbnyV3
SzZ8609hEACgr0xGbCIcCJtgUu1kzrpyhoRD/1vGNOHbWOa6ygiuICggyXvBD8X7
gtUF8NPHDrWDZIPERF2WDXoa25DtbnT7EblZvO2FTjLa5La39VWlcZitj+MKHaYs
IR8s/4tC3zGihCKRC1NGXTyYFBOFCvd8c91uWq5HJIKsV8wdxlKARFO4PZMg9w1W
t4xlZGMoYkOe4iayONYoR4/0yapv9ieP9NcwwzF3PMTiiHrGarXhYFqRelkzKitE
PdGrpMgLIkztfaSu1MfPpUYGrYv4/hucDvXLxmSgdIPT3PCXj/IQidBFpeZNpNOF
SfDVznGOYmPqsnpFzRCo7UIpN+nbQmxiiKndR6PKQ0lmKlQ8bgOxSlD95JLNzIIY
g5SOlrqrW5yHRgiP2+dUBHDgaOKwR4dNsx4miuZ+TMiFOfh9Gr9s9R7OC8pDTiuK
jXOHZTjqgJreXH4LHvg2GQQjvbPzj9Kn64CFYqhzg0R+jn3tDO/pupoLoLWUsxXq
Idc+FvD336mnfdqOCvPw5/sYK0cTeA4wqufePZtHafKP9UIxGhYOv5r9NZSb5ei8
+cimswylZLl6MoWmZE99kladK0fonruHN5cC6XJ1SESVXCQMgPxf/ycJir9nA3q8
V86Ei3x9Lp5NGrHVDC6KOq8c7LC4NEwf57qBCd+iMfaT9lJ8scRF5AV26/9UiDE6
2uZ8gy7tEyqOQodJeqn7KcbGW0ytP0qLV1L+ax6uW6OYEUAyQ/aOU54URgPbSCkm
t46yvt3vXvSMMXNhQFgVs5QGXep5SiUjs7aglO51IVTdWWzcZQkMFKOpUhIitDHu
R3Sz9rse57YmNQ4hTQufwNdX8QytPuBZ2qFxDU0V1jm5evM/F5WWSZ2rOn/igzPl
jhjvpApQ4hNRrAYZNz3M8ilhIXG7H19iD5lihyGMSAIZxBcV286q7q3JMH51imj5
HwXig4Sy+Fr5ujrlHH8fTGiZK3m1/MbcefVbvSjat2In8YOJ0qJmTrbN4SlkSDAO
XjSBLqTYb8nv37rZa1lhT524VuEKtsGMCUzk7PMnDxDNuIYJgFehJdlkaPQcWkMn
v/kIUPFdmV2JhuxSzze/wuz9ILFvhP5O9IBuX7wTQOrXSDiWL0u/THsW0zFAu4Sg
czjnZKnkHtUtqsGNWJT/u5VSMPo84EHBgFHRn/pnWLw27eGT+e8eCTUIvpTiNlwY
9AeaLpK3sXWLKQelf1kIPRZThtggVCAugeMCv9dzvzqLKhtfFs80NsajvdrOabXS
3/H9Km1v3xOhY0AyglacYOL5/WIFxFrNFzWu+XpluF1a4I8/nC3ou+yCxRQlbVpZ
O5a/OUFLFP87lUnUg1TTdZ+QMPT5G6pT/04bAhRDW2ayESDYdrJXtPy0XRJCzkZe
QgOBqky2QM0dwchW8yPcJoDRAWlww285TpPqriyfvv5NR0rxa8+BRZMeEKoUIBdu
fIW9qkNwgId71epOBkPjiYPGA/ZhyfdmBvv5V57esYn7SYjHQasFJ2LVIYH+PIsv
QrWB/5+ADymIg3mgXQCl42zj/gHOhJQK6Cwr3oUjcE6G/MUAUIjHIvKWDgLLkB5Y
Zx86MaPVQz4dQggcrEcRhnBvbpXzVzcvTs0Xbp+qEHXHdjU2lA50jDzuQuamPzYa
plTUFnVPQg1cEWX97D4jgk2hby75oE5p3mlvBn9Jj4bDfkkgqpXPT38XrkKixckK
kN+/fm5SlsCF8nu/VuBS661bCVl/xJ8PiMKU2XSJWXr1ZRGN/H28rt48mCNnItRm
gxOkZFMGEQH8AnN7FYo+VOEdovwFH0sEeYzZANeUiaT/GGYUxvHXe0J/s18z7TsH
KGrQIhiqt7eNvHvYgHssrI1LhFxG3kW8+Z25BKUKxJ/e4wgsdSryH1XCH/FpYGAo
2QiIgY+VYSJZCmeo6whYjceMw+GA0J4t1rUN0rM24AiSRwVUC3yutp970ihcI+JI
Rp+BcZTfYxpslD3a3rUnkqrh41Nz6kCNy0qGe/cCNEs6dYM80Dzdtom8gOYGAeKA
IZv50eg4hqpxW3+wlG+78fvrgJU7OHqjhTi4YY+eljD9zYafITdWenT0AH+Uo8WU
89kH+OvUrM/LQqtTI4kDkLrN0J5Sj7SvAgvge3cTx4V0paYhx8xTETy8LOsxzCKQ
KU6gVcfl3kfKUHN0jTaseQFlA1lHfwBuTjVSUwj5KGiZnhJVNqxl2dX/G+pDUivu
xyGKyp73RXnBy3bRP2163h9KFLCyU3jBKfBl6nxxJN3ccXU1jS0sbawKp2JgGsDH
H1hlLDNG8ORuNmGeY29maZ9hlhbHPJ97T2LDI5Euzsq3ZwoH6ouIpmyBjj1FU+wm
iPD+zkhGkag3YYoNSvbT0GIKyXq8TPds84mOPvg4D6Jz+K9HqnLkZtJd+JRegFne
jAOfBMF0F+aTYmfJVNyovsnorzJ96xowk9+V9FI8rC4wTkE5a3pSoiZ/2dBtXyCR
ddivCqHtKI5Yeq0Fdnfca2pNQOAMigUMsDWNm7plkpUw5Ufj9QxTSFX8aDNf0sRH
RY1C1ACICUqOp2y5pjyhUD3nAj062nS273dM2FrAh+EP3+moc3nte//ssNpFDRCq
cmzMXnSfzID5XYfv9ROtrkNKkWFdV4JcLP7DS9pEEVbcDZVbqFAVcB5NWtbKwUbj
H0lOm52DffbEGshyJixilXWAxBRL1ys7MCaRNX41VzXl6S583NFkd9p4wt9Ul/uY
Bv+9QpRn7SUf/UlaappbRNvCkDertFqsGe9m5exZpItcC8BevM3QtPxZO7f55YFF
5l3JyAiom5p1oRwsOEUXHSHOJU2rFKvFDrbOp/BEht2iR3X9RYjZPJihj3v5p+sD
jSEbOnZAP5bTZdURPhjzBUm4BSAgDvappf4PS70dcjlHnj/py3Zzks7+LBcw3eCm
036pmJf23l0Wf2+6OPZ+RjPP1rh/0dFkB8DD1I/zJzjQxLTL8tyP2kYhY/e76p4T
xOiH2d4T4vkaKXmNaTkCCrhnG4SBkWmoaFWkwVKShbuy4jKwCQGQ2xTb4QI2ZEsG
uMCeH+izq7YtBkUVC/g+Pxi72F0uUS17Hjh4FENHUgYoqzbg1yBlYczUNyKs/INZ
EVE2Ze4NweWqRYZqLZBGkgblPSeC4g+SlI5702bHecAgkGk7Ypy1qrlnyLJQ0h6e
bEeacgeu9E1zc8JcN2jlcajJDA20nuXymohCa2PePIFP/+o9Z5+MGFIdkKFJnKm5
gN8QffinhXmSPnaXELXfYBBi1V/kerTHhy2LnUg67CM=
`protect END_PROTECTED
