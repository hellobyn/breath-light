`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y54qEDYOO8KKC2I8DFcYmWbJaNXMCdqD4mMyEMDcKwJYIDp18FBuFQ3Bvky6xyzk
PQcCs3rNIeYdbb2KtbfDAtmG6KupmHBykEfz9fV5OgqDpFV367wGiOD6ms11oCcc
iyEWsCsb3DIvAmAgp7pi+pZUi/6QcS/Yy2wf55XRiO6kXfVzrdZFJ29N7fXwVh6F
FPVv2kyfpuGvtemjYucMGffn/mlqN6Fvs/GuASbJxphYyYgaMbqrY7PGOAwWR/Hr
+stvYQavyx0ev+HoeL2xbHaYPQZIkA7BismZrequsCCzGPNBW0jE/XOiOwSUQPq+
9lX3+3IqhApLRcoF4bXUE0m1A78fRIWjFyMixLaAQnwPKPZI13324iJEuzQgKq04
hDSR5xnEnt2uGXJflop9BbelLx9eG8Hi1Av5GInnd4C6mvVqe7/fEQIoIGKZx8ns
tmLqaZckKxrGPqFv0Ai/ZqFarhqsb1njmNseM1PvGYGeCh+h7IExbk9UwqGM2r8d
JTFBLESZNNSlQ97LhpwvHqS+G8atZpaYKwE8OzDoVoHHEBq/53KyLlKl0seqfQNZ
oXylEanp0p6XOIinG7FyLoi0sz1kSoiuw5KRdweNKAhpDSaULZlvKCRZj3YRXn0z
Vb1Pz5UNYER2zrbGaIO4iktMdetLnrFNfMfyEC1uwDIlwOuYfkIhA+pyMzShVwOg
rvsS9uIUKlKuP0AeJKo4mjUSWs65sYvkd2SmDulDX5lisPX49QfEjreY3jpbH/Le
54KdhZf82tGlThdynET6S9C9DZDZ5a23qlGJT23d+5Xc299HhgdhYDLTEGFK5arh
YiLRZNlquEiAq481MJlC+zNkuO8Yc7EeMbPEtuEnkdLRxOboQZTUYYsLTEeMBeKU
7hHCnyx7PO7+wvD09gK0UkRTet1W7qUluLvRAx4ob/ZATfBV6qmrSGefDgI2x3o0
PC5k0cz/U03n/3oBsNYPyOmB67w525VCaoFjRtE/8w+NRsIAQfgttuD7QmhdGs7o
KwyN6cbZjuULnrPHWALvtm75ZbT5ri+TWt6apUlyDKbmy8JauMeUwbkEWsxqFMTp
4831RGxxwZ1VGzAzP/O/i0jDUNASZXcyOy/+EnFIDrl7gDlZClW59FAStHmqdDXg
DubSQhRzu5WFuDOfddEtP8jxkAUI563aTQ5PzD1yTuiBdwRpnbJEpwHyhjHxVxYV
6UGMSyYQH2GPUznAoilUadqdF1JcR52rlOd4NZIHsEvLiZTfmV+6M/zBEiJRj8aD
/Y6563zvO1tvkDeG/c0JYVqCxuF6FSDC5I7aF0CX7uAd3xhYySXVSA1Tu9G4uCKG
SBAvJNo1f0AzKif2473SHrzR96ILsOU34sOFlWBge1bH/naKw5GUTfRZ36fc9Nwo
weJhmPzaIz+nqwl71wbDwI/VoX/+vIp3l06WHAmt0lFgw+u7webF8mablkeK4Bye
F/5OMjabA1AvIjit57KCdhitVsUoEDw4ftHnk/faSPSTNy3SBxTibvrFAu41KdHN
z9fv32e5Xaj5l+hnT3o2Yx0FFpv2RH0octt8Bt6/Iz7jzq5nrVUsnXX1NF2GKAI7
/B60ltulCPvfMXSGsgdT77KSJ308enuyzl3R9BfffDD4a5EGoBoFcYIyad9repU3
98Y8I92EosrldK1RDXr5Glek2WolyjkdMKHFy+nQUHnMRHc2M7u9DfBL9CNJQoXT
ZEuiF1DC2AyCPpBfvk5PPbVNSDeZ5QeqjrxBtm9DPxhLjX1mhnAHibOp+Axjskpa
+G5ClFmVnw+DhumPPiT/pA+o5Gc9z7uOIuUUZ5AHG7HXbKvGBPThblvjiCLl16vb
SFzd72uKHjT9YS0AMLDE5ewxuS9AD1deFrxJUPXIJku3/KJCxKikKGhnYWQ5sLYP
CPhLW7zGhtM1JwAz3fG9cckk+qzw33d4AkK64LQkvn13IzLFOu5ecoOWFEf5HdRf
iB1qi/A20djqmBWl3liY++6H8iKPz9Mgfj7AMC5yDxbhsjVR9cTaZCj9AyrcDEv1
XY3Pc1/IKq49MtTynBv1dSQlYztFtQKsy66nk/v7LoeZWfio5hmFfDCjuSKU35hn
U4U9dz3Cblqf/jLOwLEb0C1WahqXgOvXSzCYEuWFu9jJkgsYiArVK/ID3DCWGfKN
0/evOB+YcLT5/qPah4RN9PYsS+zpmpSNYRApL8J+8jIemofuz/KJo1nun12PutVg
ngl6vmmTrzsvyJH5S1f8jT7xhjAEVyP/ZNXhlC1+QEIqGXDiIRNA1XYCdZqdV3pk
nLRI93rg+ubSN/czo1ne2oRQKvCRa/LmrJrU9MpnFpG0c8hU5A+nbXAZnlE+GRmf
IKGU/bAX4q1fHv+z3slzdA==
`protect END_PROTECTED
