`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgkQ8LInPEmWpY34S1OH6A9OZ5HEyAib5CFrAcfOAL6n6NMsUwr1tlMozYdDyioQ
xuToyLti4gSHK9Dnn3XrhoqcppGGwa15WFLZfegvI3OkzPqDDVgtEv0LDZglrhCi
tSz3EB8nygRmkDOf04RE+6AkD5Ps1+faGvqyAomwJ2guW6Cc8ue31qIxwrrPm8bT
cpI1mUa2P14rIJvJF/FKM8/9iFX0EwTUl1F7CL1SQLoIYQaPWNI3QDZcVo2Oy43z
0yOjADjlFsAWgKrH2rnkXSAJCIpv1yepGKWzcclWDvboAUe4rNe8+QNlKD8Magnf
M33FX7sJQJWvIc6mfq07suxVOqSTY4XMNfqR07KVgDOH3TskOZ4/Pc5mP5t26jTb
Zjff8hi3hH8+KswDPhPqEN+rMetrdZae9Mtgl7y1epO5AYLYfoLcKDw2faR6C+tf
VN/hR4PxGWJMN73i5rQ5eQ7jRE5o6WXD51S3tdSGmrIvrouc0oTzrAPjaPymaaml
Cg2c9v3lYBtDj60u5FuPMYb8qNf34A2A0J3ngT3tZnbey+l0ksrrIdZcWPsqthPR
348s7S6V0Uif4ZDUbnrEHBkLsPjz1HGbgS8RzkHCUgZSRFg9IwYgIuTWSA3UdLsr
tQqxfSzr1ieB7FUoKzJmgOFShknOpmUwAtKp3xM0v1PwW9Rf944S4GB8U4rvuk+Q
3reOKqjR81kLcs+nBfuv5dMNVJoz8y5+6OLxHKgTPZsA/Q++iFEJV/UlwoZbiig6
D30PwbE7LC0upYzgVXWPHAfvpTiP+WGetT477zJD8hQQv3rn0am7YH2cXxs/i7BT
4Nuuvi282v5JqmDldWimlYl5BreNSaPUiMEAlVSXihNHKqUtc3TpukKy861GLF8B
nF+Tx0c5a2hV5zwh1j6fq7SM1pulCcYkEyb0/ltlpICBIr8tu3IpbeAN0XGNWAmQ
/+jD53l1yzueVfwDfc902oroxNlukG+DiRwK+JDgYJytMADvJI4FBLywS8Q2V31W
FPxGkYoCGgg/kkiKFwiy7u4SWNnvGu5Mq/6RvGBin/b+Y8BEeSYBbKv5LIVD4LjF
lt1CaMn+y7Scoa0ocoxzYjELdqbM4LabWevlbLYw4fTl/oUQODvrm+3Zk3As8bZ0
zRtHZwLeHzUXBLiNX30qLg==
`protect END_PROTECTED
