`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2HvOwSoFqiU+7IgC4mmwQA/F7icvO6eTp8kai+KJLki54UUEfDjr9ssbts+YRE7
wyJYprBg1rKDaECdF1RhuAmP71jdLjO4A7pJj/Y6OMbFH8xaZR+R024KDa3C/33N
T1EWRcU/p/JQnBsbeHokeB3aFIBkiOHtdZOh694pJALJ7qukl9ztTHOm/LQ0uCVF
ulQnrhDngFpmRJvsKrY48GOp/TGVRLgq6uI8EOYsLHg0Azy5qMNpUqqZUFKy9ERW
MmYxwDq5nN9K28kQB0MeNpVUlh2Fsj4lNKTdKro3NBZUlwBNxL6uI+b6Mxk8EdqY
uBRQucKgHmskE+u4OvlJCKyaHpe6lIDtHtNXFymLQYpSHPbCUHJP4s0a0o4HMR7A
jphftwXl4QQazVzZBGWLRGXNWUOskRuvkb8eHEAJ1VNXDQHDCEtSVjtShfaBgglu
N+RXTwkCctFDt+lFRxCpvdxKupIxsplLvpdKfszFiO1EHbbYdGBwGdkD7egilsCQ
9+l2kXxaOAYflG7NfdQajgNPuM0y6gyYEDLl8brOq9fDT+Jr6ZpcAWSURMxYZpsk
aDx875wecDE+7WlVbvAz0dHDwgbIXPvBjQ4RwbzbthSrzJosp1O7y5B4VXXvbqHR
Q/5xfMfeWikxioJqruJXRkHWYYnYYUjO9HER7FVksG5ZfVVXZUK+scl3otP5KH7y
gFLwjezLoK054Ab+FMKxpJ6kVv8e+HoCo3MTQC3N0pBEjTILEYIHnCIviPQ6aDex
N2KjSr6duF88nSuf6t2J0pUi6BUVky1FdLbzrAqH6XCGlbjBcYbp7lJODi7yOD7Z
IonB7o8x6QBrhqtVI5aSQkqEJ+T46y4sBHUXbpjZMFlRBWc+Xq9qMorEXLv8O/IZ
0YG1KrAHUAUQdkxW6NS11XCJ/AqJeI7GxKD/WkMfM+y/9kIZ55MEc355VzJ4nPFK
yDhQV2UNRXg1TN/mFvAKK9xQ4e/smTGAShrUTQ8HyMTvIMKaKmOB34NCokcvGTPZ
L5/66pC8xabC4TPLzdXhs3bnLgPSB8InGB83dFOrfWmkzcofAh18i2faDupbVh1+
aiGjPTNm/dv25mCe0JR+ogwd5J4auAupaauFe0WiF8K3i6QFwIWnF8uRD99ikCpt
Yt5aXJAWHxdy3wiUk4qYOdZXln0d5saq5+h6VcfNRuU69hdsADDncglxSZxHEx7B
g1NSuM7CQInFinK/eNe5yC7isSV3sR8QDlexAKljjmnQiOO1cqxYv/J76Wd6cyvJ
sOmrKMq4lpJzOKLtTygH2ZtmmQLe8tZGEeZjWxJ2DGpEjlEUxoauUl9rhmjXJI89
obnkZlXuGhmgBYuNjTeiRJUbUK0notARfDT0BH5UNzr9I1WxK/+rGzGu4mf3M0BU
XJxkwEf4wfJfiOeAodf5EVuE5HWLP3ufsTDfyTL4tbdUdzHqaem5NMGvdLS1msCt
jg1Gwi8qPJ6ibg9xQgffRO9H5bP8l6Ed5sFxe/afzfTLzrzB/M69Xv9334o9OD3z
bC6TQugUVU2MB6iOch5+UmcHy6JaRjPGUKy5kDeH5JwiWhTxQInL33wcadH1PxcG
TMqe94g9hNQy0H+AS3f/MJ7prLdWlgEDyrFtY6b+XE/a2Q58jJDrwQMl1pHi23Be
FWGEAjUB4saN4LSduXJsoTTqIWmrorT+4SGNdYYBshkr90BJSOxEPGSpT035xK2l
nT+rqBwG3GEc4ZuNNfzRlTJmDKwOeI8hV2Lzg69HmzPL2PUh4NfNdMsEJfJgmKdZ
mVr7HqTkXRRglmimWTfA9G5XVGAdFL+MDyC1d4DpUvk6GAtSt9bGXCw0R1HbLHcH
oP6zKS2SqryAAviTGqR9sjVP5VyDAwNfJ3oR9dfJricvMDomU2/F00BSlKWKnxtD
tpnylQnycF2g+MDOMD+fc+rouTbrEibOsPMMJlGzJM7Mn9dGVV2B86YEeNhN3W6S
HDPRqAUgtHnM7Q5vCT54LuO+4mI/o76YshwaWSFMbVZ6EQ50GFPlelSczZwCWBsM
Xbnz0ecAXftCM2jMKd2okzQvej0HSVUBsfT/2ZFsW06zG0vIfvhXflBis/QXppbQ
B/01126eOwEdu4JZ05BkLNw5o1Gu28a6VXKDqikK8mrqAhZIbmnyy9txtOonnN/j
+OsqsgywjPiWMaYVTY2G+1voWttXTbxN0SuXEWx/tEdewIq3p+C2Qc4dSHatij1K
GNFHJhksBQvy45+vow2HKZfLVKcMb1reSz0xHMNLp/FqdJkJCSpQMVvRjogmAUH5
dgevMmkQPzmxfgxeiPMjRNA0XY+xCbOZhoUCE6gwxOqHU8SMDekmas8KfOoiMWb0
smKAjI3DcmtA/ROGoXIoPhIngIKwc0bHLIMf+XWA6LyH88hDRl2Q1ZJvvHBDCuj/
O1dXA3v3Aekb2BeLdmArN8ToBsaChsg3ReN72BPCW2J4I8mpKQC8JVoyRUfByuJb
X0mKBWkD7ZoLEDrVbsy2maMhsbE1jnREII+MhgVRDReTejBYWuiNTvpA9JBfodJx
bKkezyDouVY8XGKOdFP5N6Ce0QK+LXhGZEZh0CgXs3CWNLVYSYARweLxk6a/LAhk
4sZIdb9rgyZjlFIbGLKxcoeIWOpNs5WoLG2660RunlpfQP7o9x7h5yt54ZSQjGBy
3BEwHMxYzxxEeBGlj5P9hLvsX5/ebTJ9lHDr8uvVMFa5BdLvpSo5BBq1J/88Q4dy
aw/E2RWqa0m8j0yJi3wpK5ycptr1vMvfJzuumdwd7THa3Il59DPAYtrWuzX8fwbM
I8TMBgrl8PuXKdkjo6+Uxk66smHEM0s1M9uw5y+YGQnCxAbxAhCDroeaouhYzSti
3cYGNvb4tpzERPcpbR8FWR0uIyi662IkV48rOrw6yAkNoNX9w+kC9m8rxxiiDLSG
fZn2LmQy7BI5OZHqJSw+T2KKUgZI2tl/gz1yhFZGXHU=
`protect END_PROTECTED
