`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWH3pgIRNJkXMaX9CgA+hB+XUTAxhGOHvR0nQ/KrpnTpWc72Z8Ljd8+zW1h1qVYp
G+QQEqXoauzVtS4rgi/LA7Qn+yjGhr4/j6ZP+hhKPk0PSCNTkrSmkSYBAtBU/mAs
phHoDxKe2jQGMRDwu96Uts/CCEuGaPkvsnmaOCd3k98uce84UfAw3BYKkLTGmAH1
5URpea3DJRrlmZmfAZyK1ZsqfUsFvroAKdRF+1ZY2/DqDSVl/PV9As/Y10CTXsXo
P+E8FRMSgvu/IQ2N/xR5q4Yv8YnPSXgGoMEqBSW+1DIEBOAtRW0+axTuWqAeesID
mbevQwFzo1qRkbYBV+Z3qhmx+HXlP+AfaIxVfWW3P2g98AxjV1QXJLAudsrMzryn
W/7ZSl47gZ8Uwz/2aNE87KUkRCvvkF0/kAuXzlKfkGWitjKANnL1Y29pMZ+VII/X
+95SBS2BhAV6XZbzMYpXwB1EJuIBtCnF+KsBX8T0V2IJBs6qR/rMl2B9kSj717KB
gGRz6ERqVwNsDG/IVRKe9z3XD5rcY0ojsRtu4rN3jscSXRJ/bRDrK1c16fMGE8Cy
cJ996bohAl4rH0KWAjcFZmeK3l0B3oXZvQADJdLg7MwoHT9JLz37MZdm64j4FedJ
HPU0YQQAt2OMYWW934nzOaZStMGDNITN3z8E9+z7VDSbQK1zm8ITTY3nepjM7nq+
RI1D0bkcbrXg4EDIK/oNz/i/RZzvIRhaH9SloHQbF1ycomMvSXpi4YZwO0HAG698
MRyIqFCd///NSi75wblegwuyc6blgp0FWyS4N1bgHH1NvK5sVKw8gYowBRGkLliD
wInSU8caloo1p6KonyC383ZMXVOHZMajChpAhzVpHe9KKOof6PuXK47TJSbvP3Nq
kI/RASOV9x8oU8JSOE4pfxt9vDAX90aSwFeEe/RfAocc/bxHtqNSfV/+4VIDe1bh
qHmKV6gPoKOAdmC8hDSu5ZBJYhwFyTllGSrCRpO3Fj+3YpbEr0OHA+QHm9GyS+lf
dVpLHzn34i8aTYpmrTRp/u4WsXeRdwAUiLEtA4R+iNRjBEWoE6fuAFfJm7Osx9l1
SadkmU2uYlEABY+KaNFD4wliS/yl3nRolhynpinK+pdCgtiMwePCEOWTgiX+aMoE
JwXxw39B8YJ3csXkdQuxpL4cL0UMin9RMoN44KvzYg9jeuDfjUY4ruIY0FPAq1qJ
8AJXq/p8hnMO0/gQRFfAtb7Y8b/nX2/35LyOUFmxw9wVadMJtnEG33t9m5Vib5Ge
k6SvSFD+IRi7rY3beK4KC2ENbS/yFF0r0h/zae3T2tgMRdyEP636eQT46wqly2Ta
8y9rDxwx21WwOLT2md68naalPXIgtdy2CNAfGsh6Sk4C2dmI8M2EOhyx7qHSjV0f
HqnaLbFp+NZBklxPncAJ8c7yr1252dDlc4e70kaYZMQC3f8JUfWR8IcoIAJoBvo/
UBTx/UaBlH+i+knpt7NfGcGUvFgbwKplP+hqtd2vCRLWzue9wa91uNioKPFz5lJ2
iim9Nwua8GpyNuHhPLJE57NUzg6npry7PBQREPmSWNqy3LtBmtdEDvgm9KmXQlym
ap92XP6JNX0swDYAaNTXyF+E7HsAwKFDUr9mtssBoNEkctraM/jnHOsRTrJu/OuR
xeHMTdphTBMqqhWyrG3vuyMg5KQjtCm7BP2GyCKcmVbiJ1996GA7A/ZwNzFCi4ZN
6OcmVFlvLv5A6u0J1MQXIEj/nY68xZZImtpOeyMe9nD8pW744GqpbbJx3urck17P
clB8vpAtA7aidPITMwam1xMXTg+xTmQ0xzfEf0JcpfGO+VYgjJ1JHI4uoGaEmQkL
VSiJtynoO02Ys9J8Rk+XzXV2jK/R7c+0YTr/ZCFPsUQ3Dq1xIIFP5r80L5aTFTWD
3NrvvS8eruPRPHVEmO5J2/Gn+SnuTiph/0NeOIXrKmedPT9pwQNgwK0K7adXEXls
7fdQxuHQn9HikPSS8OsVVkFXeddwt7lcK9j+9at2NOmjc+XpteeUEpOsgQdlgZnG
4GE5O4232zVZEsz/qhKZY8gBVYqT3+nlJ3FnSaDPXBaO42kk+MD4bbXgAB7NqOYW
XK/mI3233XgsNcY6ee6tfQJgOtVRukFPQWrZfleILoQSJdMNXeIKbVRwhuQkdD4b
i1D3chIiNi2D92wypZL5jdcnnXi7S+oToE9O/2iJeu3PywOzVNFFr9mSiR4JmoPC
+W7uo1NOSI4ZJG4Dki6ZqAxu2ayKsBTW7/RKy7Jwbo1mhr8Bv32q0cAUDZWftrNO
uwuilGafvLoWAu6bHNdaOsmJDL0XR+5NdKqqVCijj50DihRlZXye6XLuCy8YQww6
yy6sf0RSz18IDY/nnkZ3UjQdJhi4lQsHZhvIrMmUA2kf/PMw1/4NluEeFJ/svEDL
AdM5EV++BrBtNXXgIDOHq6L/+nwdwt35MmzFD8g0CpK+xRDK5OhWzOU0jbAtaGpG
M26Q0vJd7taxFjzirOv+ogjJEQw7/pTBxFrS37xnsJi3vxo2W+NI2IlPbQIQCdn6
P8vg5vaLI3wgaiw0HV8+nM3orjLtOHSor6FfQdYcu6Ci5Pxj1A3uoIqQ9uUCrCn7
ZhCPTfD3jwJfTAUQiPX6VELVKHDfDefMdWZxQeGOPXH6yAOefbGO2sAZ5krYSR0s
UCtsJD/s3ztWoL+d6bhYs1SepH0f8/ucYbKiJH9IP2cCexh6YXbvWmoHbs8buufH
UmrM1euKVAqE1PtM37DYV+Mda7Uo+si6c2195Lt34WScb226H0HmYAi4nK45bW7O
wMLYlIwL89ODYpL5+SYAzj2S+Cq2tggWGvovioukfD7znqckLPGm/rvxe0vUbpeN
6bs7ue/MGzYQfwgIBeOlFTfKQkT+NcRouyXsqaEehuW8hVnrIJnAY/CX37rwNaR9
ZzE09PekmBs/OBPvCtqiTvTBdmn3e846ZUiM276JnotBt7UqHZSxWYsL8r19mRJo
d4Z+hi78nQDv/OCzzcUUJN7BxC42HmG2fvClULWbY8lYMbOLeFe5ZF3qcfAnJ0/B
pTPw2gKrhYUg3+XKlSqZdxtTB1cKR0YIOcM6h3suQGaHdteTWH1z34pL/WhKUqz+
1yNUa9bFWUwHKZ+ynWJJD10QAvl/+XiSWmj7EJyeFjv8BFh7SDSLLi9k9eVo3i3e
u5ou0Wc/1wEqdtuT+qn71EK60YY1i7to6uceV60JwEli71jU32maADVhIsfs0Q+Q
SuM5KxPBWiv6AwI3ekMlD5DbG3HI2tb9CWQz+e4/8nv2xxmAnv7WSvrkRCeboNih
CPw8/RUUXiLcLpNXlz3w5rgaql06XFCm48GHIkdyJ4l6GmxpYAtkkjp7OTgyGh3L
cv5LTQLhpkCbmBlUeOD0KA34HaoIpXyqHPixwtFG8G1JcQ+htZnvelbtn27rwkdQ
hrZ/vurH6xHaA87XoAulrhimafS7/rTdR9XI2ZWzI2wPfupF1JRSBaHGZweAd4TR
k/DuGxoHlnMtN1ZOXFOHNl8scQqa3YTAuk8BI6fkXO1a25pXDLNtcUDSB/1XBBqK
20RtVsN3SNYJn8tD3eCngoxSpEv6I+eYu+DZ4AQiq/VPXIGT7E18sxjlZEnxVBdW
gXuniqq63cGrDG+ptGVdBgnoo41Ek42hL2cWMsecqkl1ZpZjDu55ya3DNSoWzxB1
e+/4PWTyutJ5NgNTbyQEw5dtyCSmt8EKU7Nx4weDJ233RdZ974A+o3z2wULtv3mJ
urGmUbSodjjS+U0H4OTOQFfmgSxR16Vx1QM2bTDMMJ7aWZpbh5SgV28Bl0dZX8hu
EuUKpXyNyqibT8MlErS8ose7FIz+OQN/pJLWfQOlJXkVHfLUSju7mXPvGccXFLFN
vdKOUH9IHufwM0j5Bmd6kn8krnt5GljS3/BOzuq7KfsSy3uGWGbmStmyrkVPm+GC
hRPqSxipWtjzIN8EqF8l0mmmz90zgD7Y7WInElPwh93g+RecDmZzVAJMz0juG0Kr
UGWyNnw9NlAAtajt9G9GGLgaw80psRmnlh9M4CQK0qeSVuJLFEYk+FZ6qw+U54HT
RDjIOAy0Wb4L7+bdYWr8rD90pMsXvKgBDJwLyt9u44wuQwI/zbfjuIr5YeKLLrWJ
m8jPptUZq2rXJFXTAvb4KSbAL0LeGFljIHSkd/bRfUYvID0udMQceD8HX+WzXCMU
WDQid3ESQY633R855IiKCOuKZ5z8jmCnAAfuuvzGj8sjgm5ThevBQdYxHZbGNYDT
25qblDdN9HkyxQ6jneGwGar+b9iZETaP3WSzsd92iBFJntSaAOFrpweC8UudFwqi
j1TNv0nk58DX2+/NmluOBYDFjHlbehR/dSbbc7coDjN6aOrfkQHo8GsfsGAF9ykm
ppKkc/1Q60LfsNFDIJAcMlsfRJai9JVMyin04PpC39GX+0NY4ZCPDUvgHb1IQ3nA
S5+boC5RsBnsJZsDEme4zy5Iv3rts2Z0plq1XTyXzbeoOifD8Bh+1LjqY2XbwTla
SjdSGYsQM5ee6NQzUUHgZVSIKDMcDp7jYz2Y4wR8g7dJASlQh/UZ1d0eNF/S6psD
RzP/n2enn33c6WrG3v6iZWfi4t/QRqkO3Fg45rHLoyPpETJmY/BgpjTFgDKrk7z+
+TCLHBX84aPiTumHUxzvx6HZK91ICArSZOua4LanhtDNQgfSFTvvoCREAufzgbBK
DIRTx/NB0D2SwgtX/aogKICcf04CCdq2OUSRXzB/3TWEsB9ezcnOa5GSMs1A/+vf
2A56hhvyCEKg/rKWurolToSOAo9IfTXY4EkJyAEoe1pKE6T5l1RRHBG1RqaK33GP
kMhY4dlaJge6DQj0sCNZzJSN0cyMVUQTpLtF1gWyw6ptbIdwtso4Ztx9iNgvmt/M
KBFDz/7yujG5ChcaiPBT6CwbvvaOuBhDn2vjdO7imMjJIqqjq6wc61bebD6SMO+s
Swb7CgyMmysP1yN6RN/q9MKFnTRyqavQsVldE0JIPeexpMWDtaob6NIZxkRKOBqq
K2y8pD8oeRu3xxytv2iT9mSuyNmK+5jkxx/7Snx6wRiyTGfqv3XdCnUg8Xh1EmuO
zfSEqw6W/UkcFG7lgX7frrajZXW0Oh9fZxGGTsXgd6cLAccXHexVJ+WIxAev1LGd
mG4gqAob+xeV6dSBDlT8gPOvgJuqiz+yn/OeawWfrSxtYJvhrGNgAxRSNHHmRV/B
49KImovQ6bL6H6c4CJLc9DuWXjNIVmfx2d6eL2u9P845fsanFIKBwnwId4cLAcsK
K/2G+a/u8tfHsNTPPMb9rtb3wnbXEYZkKRGFaJq+/oAeSNI8uFNekutPldFRqEOC
X9lGfJSFCErpD+aG8IuzbEIeh0vBgNQ+FkVVkhjM2qbxRfHF3zL4Qn/efuEZsxWj
gBiENhzQCmfY8ci5eJXImYgQNINWpvwG0+ALjfs+6ZAoVRBM2uEWOYymfmsP0T0A
a1UKj+RnyPjjUnMj4Kj6YT4aYXsH9Mm4gXVr47qET0fGtGrHpNnQ1cEgbAXwCN6q
LwwzObZ5Ydu8GuIPtT4S/k0q0fj0pOWhwQKeybVF8sbe3Db99zFdF60D6yZhhPGF
wnMwtfZb/7+VEBQ8HuYvpQysqSuWudN1QU7sOABiPG3gOm4WwABS6jnJJie4eDJr
skA/Bua7zsIIAHsbd6iD2kFhcv4dth+3SddWLHaXzvAGv6RAW3UXa1/tqs8oCx58
KcyZcuJpA/1pJvyJEcKXQMdrV7yEx/LTs/rLg/9uuTSeVPUFu3heHaNc1NljzJb3
r1hwu2xTm9F8frAAN2vorUu5FygZlCOHr94vgTGi1ySJBpWpAM3mX5r4NkyLNlkV
Wcm4yzDMv4ALpazGzECAlmnDfROkk0xQYkazdI89YX275o8kDGCitcCWPEbC9I+F
WityOqnS3DyrmfdwjwQIP+7U64whhNLh+uDJox2IIbFfWAwPmALUc/Rn7TqDcnmX
tGl46i8Uzxq8za0s/QpvqhYjIXgLeUhBJcQUg1z5JgsCOWGBSqIX+xYjQgbgmIUM
UoRW7ifPhXsTIn/VFSN0CorA56/6EOrIEwPM/2QxP82a8pDO9VZhO8/NulD+yAcz
OoHP1d65fityA0oYsS6gLqOzIvaVnLWHIzvYBwNnxrFnLZIMR6XVimWg7E+DXz2n
u7TncYgHGtx+6Dtd22njejEHlO8z7ABW5ZahOVacZ9oVnWW307I7FltCE1ucmud8
CETDBMLmgE9X6uDGy5nIMffOIIh16fecxdTC4Dg0p0XjYwfn5TWDYaJ0oISgDv2D
TpTeyII8Y9nH4YcDCnlXqDQ4YOGRMnQpkSp423jy+ywguL7xdBTTiD4Qnn6nyHEp
lm4B3/qAlFc3vMiJm8Ow+shcl6+W7g/uNB5CiVvhCjx0JaW8GN5J9Kgt3umWk7tU
DjUzyKmVgEbFmmPIQa3Cn6tDcg9DhCFwSy8LecLwwy1r27cVT5+POmlRS9Xrrcql
CJkLYPN4cPHSJ7tlLwP97mGECLq2nWWydiwEX8eoP3inAJ39q7YflWCgkd7Uxo7M
FrXpuEm29Mwy/PNIDsiHD+p6RP7wgCWgrZmBVptLqHx2iQbOTjmYAJFiexYRILON
nXCIppvWO88Qssv9+bEBBMQX4JZ4/HPFg8mnJ3UK57QNsWNY7FsvtdvJPkmzky/Q
3Y11YqzOSnA38cFktZb3jAnUDIBf+/wUoyA2hZE3RmEe+pUy0sBkIhdvXsCuqeiE
BmbpWfCQJ/UCyjdAoYYK4hF4FVRuLzBzTt8iLtXGbjSTpYuawWZ7RJz0F/+jtoD0
k0+4e3i7+pSBktEBzD+XhLP43lVJbGrRfOKJ5vc6+ugNCO2PV8w1L2ByBHaQ1mdo
1JEUUrIJjupnlQuUPuPH51RQ9eWO++GsJ+n0ObXJwhLJry/g09888imXAlkMCJ91
TrvuzUv6HQhvcPnX/qqWHRMRb9j11OyqSTezv4n+iBzUERC0kk0i+Mqi87VvmK7t
TplOc9FfQy/9MXtcGWqJo1t1BA2LaPPl4PpGY04nczVOjmBqCBk7PJ+wR7wRhyEv
2h1CKMUjBIhkc+5wqHnonIQwGF0HDVVCovirwvRMwTMBJex/fD28tBdmu6GESukN
xvt9yNW7Ep+PaUuYRdVvcIWww/3KojTKBL+oDvCOS1l7L3GJviA9R2Sel7NY9n9U
FzzneIe/EiHGQpEFwNyg18EIsPhmNt8KU94lkGkb7FCHTt+jg2uuFk0r+5uJrK3P
9BLppsREOvzCGiuc0hLXQJltDTB0dT+GE4guBm5imeve9Elj21i4XuIDGK6kcoLz
fM2mPmmnugj02qYpowlOedZZftLum6ZUH+mEUJCKYXxE6r93hOHnwRGRaSm5EE+7
9jkv/BQu9IunA+dTQsawGUh59/2yaUk1212iv6sb8xOW1Tkxn544Mtg1O386YzAY
Jw2tQ/I0JS1nbSlntL3VwIiBd+hv9PQT4BeCXQ89w4XCgWmcl/w/kywZnwncGF6B
UIDcTMEHFzdOXibIbyzgJui6al97X5bD9rHweAkGO7VJ15IWeqY3kh5rpVs1nvgw
5ccmEEWgCxLSEtEqniZHgtBCrfC1XDFmxqACl+2PHNhRymy6/gA03hCXKoKfvdUp
eV4hFGXScECHleC7vKx72d43wckI+9rRJTU8D6pY0GkaLUoBE9XWA5V1o9/ePeDo
OX4u+Hn2UqJ502FeGRRuhIkq7pkc2OXPr852cG5VNUbVrQ/H6xGQrnczORQGUfN+
z11pgb9Izuw/j3C3oDn7b3zXgRu3TsVp/OtvuyAd2YL1k6ARCB9UW444O/WX7+Dh
9YlApTbMTgjL8vnB1SJNT9ND1++FGyihUzLfRROinDMWiHuBEIiuhZE3YwF14qAl
pP/1aotn4PPAnxjQloNadX+5dqkoPapf93nGKt8HSv+paeRm0ZOuOBLCzl95/E9B
9SmohmheYhH9jBVaCweowAM8YcdW5KxtZdduvhWVZHzv2THWE0zjS4ScfPWG8pdO
dEysJDRn3BxGNgDjYjgyivSv3crB0Zy7PHiD/kEMh9cTgHKYeYfAWY2k6cr1ZkwF
vhAgVUb60QMYXX1KiQPM1r7aNBtyCrZzCtBYrp4B/qyTE3DSGeWeS1blxe9hjslX
oKMiKDn/poKpcQznolYpTE5X+jgJqWHs8sHjtyDfDs+JYy7xiVJgYOj9ynjznzxa
RKH8HRSbhKltcH1vBy6onzDOFduOd3OB2a0iF619K5w3GiKdnJG1WYaQgwu8zgA5
hKgNNCGwp5fKhh6h8Jd4Wu1Rwq+ZuoLy1XkWtoxCDa9FoVQWD7D6zbiITT4yfgjA
HF3ZDOhpPaVlwPRRLT9RFS/UuI8LskwjRQWE+iqezsCXiriOuGDxBq+psp14tw8j
VyYqCVpYb9jRQqKyLxptExTVKR6rcXUMbX+GgNczZ+NZO+FulPky50OA0hDfnmC/
zDokQmhCG+7tVLe3idieh/xpRSZgyfi0uQqjjTH+1X/ErliOCaZjOzfGSHYeaauI
dhgccMQ4ewmZuxoekbZuOUwvYfhcwfNAJoVRbWjjldBdZuAjJYCmWvMNM+4zGQr9
f7SwrjdFKy0PxqJzO0WfAS83HRD/Bh0xZJoPV59Dhza+cMdMPzT3eWHTBp8KLSfe
03SL4iiK+tOHm2p42vQbrXtsUSt4UhF9jIj2D05t6wuTVYPIgaPHetuCtL9kb3h8
g9uu8CcQMopebeDK5flWTJhqYePEQ9/MmgKEsDlppxqSX9yyRuasMC/gjIklyvSw
lzJJLbyMG4s9IRN2vkNFaoLWX6fDBJFZNkoD1qyOiO1T3xz5EBGiTbTybiLKfErt
cnVLKotinfTH18Ligrirtk0/x9H9tRYUMMCWZ/9uScMNALDa8hTOKiUcJnINLLsJ
8cyE+YvfXPVy5avkFZyl6XEoJ3zhqbxtwHgp31EXjyuMPgeKRsBZGZ71cgZ826lE
2rWGWA8kCasPQiLh5ZQaNmOK/RzbbcfFbAiE/w74wpnn1aYQZYUOst0zcGSJQWcq
3+vFjkRzQQjgDk4EJZjj6Prk+FUypui55bTlr9fXN0Ve8vmk/PurwFa9OBtQxNN5
Q5aQeBXmZfYSFGv6bbBu0qwoDpdaNTObm62E9wBKo75YA+frDJW/rN/QOLNgvrEt
77nblAVFoDsgEY/f1bMAQLc5InRBNYCN1lw4fkYB1aIO5B2oA8ie3eBj1R2fzYVI
sgw34klyurffWDcZdOBmKXj832uOybOXraBh5J/B3MhYCu6+B6c1s3LnKUqBcCin
mGWV2G4bhxX0eRSRsD0Z4TqRhXyuG2gUiONy/jrh07mXiJOEh30t9QTCw6hbORzh
8mvX2GiHnTXL3okq3e+wHy2GY98p9krxwm4KFDIyfNUXVU8rzU9NCi1vj6/Vu+MZ
g/94IiLfhX7OLEwGuNPbdF+BmnBbxUE14bh0snRGJ3YehHd/1ssmG2jKgPHvlKIO
QOVpwuClBi5q6oong9+EQzsURCRt1gdq+UDXUds2FRspc7uZRKu+4PMkUeqCavRr
lO56iPNj7PXSz1B3COZC9riMx6GtudWaAihPKuxThnBqAbqfFAAQBMKu8HpFHfCL
LAyeqI8ZYYBtiEOwnPIFS7icXyvn5ykItb4Gn8MLyv5B2aYqEMymihzU6KCFxOFI
kgzzOB7PN3gfLT4R3N6PFg6vTc8iNwsQIj48NpNJFJLoDp+JRa5eV+zTZdCdEy3i
y+mbQJRYv64mugTarolDW7UenUPstJSCTRY8EBNdPtMOOgQVITjVuMiuIYbgt6rL
Lb0cfZ/FXgVMEiABAdsTv/db01rnd+lMku5NKdgkyZvXz8NvIw0f+TSTWMx4dPZG
PFxoyj26xL2TRrwvjzTb3cuL3ivAJ4ptjK7UwBC4Wy+shwPPHh7j6pf4CV0ebMCx
54sehqZyOyo15J6aas+RC2OZEy58Jpo8ZTsYyec/7oPa5xYJrhSJGAbsmgFrhllg
AukSkT+VNjCv2sgRenmI55RurBDNRYRPloKbzoz9llEUHlpCOITUSPeC73pmwmke
GyoVtQc8pLs8lGL2XmMNL6cNCyAlHmmUAAUe8cxQkdWNCUROFl4MbHK/VgEIj1YW
mKQoWlyUiGOdFntpAYZg7azWlZK3cdmLJEUfeBYABq5sLVKrtb3U0iZjY1+z3yd0
ex68Zi77sU0dZrcPAMm1fkccAoMwPiMwFoHs9IfHh31OQMOx7nrA3EezCks0uuRa
/BxowoapU2UxxztlPXPoqurFUp2t9iGwVQw0/Lhy+mAY1HaNcalKAQ1LtMQAImNr
pBxWTnnFkaGrAkG3vNz0VScl2Eh6oy8/duYj4QP2ryKnsEVBlXcsOgo0l4OFFTjC
ZPDzxieMSUJgxR2c+896wd5GlwFHeb+3FKqUXmg5M57uwuxgtdeD5ERObfQIUiBN
0KOiUFItj4WpRZShunvNRkZKMlcjGijGs9VBKdiPxgIFdXWqS5Fbf9k9/ofq2/yE
Pc7lVVKi2F6r8TOtFGJC9W0lMdcVpMJp7C9zWODSs37maihJ6LUUEfu+La/NEmb8
oSzTgoX3j+w9po9WYC2y3/cvk41YgjVdM/7dymMjzhy+G7Zh8w9WUAyMTzOAxLzw
KSiJZCFRDvCYVbY9MycBBab62Vz05f0VCFxZpGuIpxtg1J45+2/ogYFb1EEU4cPl
GAXzHZRC6tqV1dAdinrpUkSDwIaxu0njwe85uvU11LgQ28yx7EwVri5I7Izy0QpD
TCcP7w4Cgyq3qX4mJnI9MMhUz8sABDvKXJhqWMD6iCYLnItQFaqFnfifRAKozWf0
j4ATUe15HlqWEXDNC2OXXr2B7tGeXVXTU5P72TEaMESztuMYYRUGPZKMkobPQEdc
7bfLLG5OfmW/9MworLAU9TU0Ez0an+GY4FEefVFslr37yn0M/wNCQqNqmPsKcCIG
/6Sr4R02U91XEqesjizjIpTUB0oa5EIZzyxD6Vb6Y5Ny/AHMNda4/9eXry1EmCgs
LhoGpqT92rRulExm24kO4gB11b9K3OQOsfj5ew8zUl0nTnNAVWnnDe+Giu3b9/He
D92NruszNkaoLnSnuh/3oC4YQja1LdBuhihj/VD9bLkw0tmL0L9NpYLoHOHc+qUI
qXzs+jdN58t6OPuGDtO60aXiKBJUksMhzfgdpm2hj6j3LGOmrmjofm1ofKOMSqjp
Lpu6Tni4l2ihbFI1hah71MLKstFwX/u1BHC4NfD2vzEVaTho/N2+P0YrA+khMMy7
LNAd8uvx1Jqx/bYpNf+4byzheBR2GQDtiAiCAFDfDyHF2x8RBZzys1x4mI04Z3My
VXpNsZsE1f1DzTnjqNh6eoRrBD4tDmKXdXcRBu5ldSqmprCApUCRl8sgAnEHNg89
DQZfLspCRJeAnJ+DKmTKWsdvdCKk2x8mci0BGr/8EIhDiayUEq1S1eax/DP731Dx
tiw4PT3Og/i/rWJWohmKauewMi7OyWABwfYyBZlw+7gd9kpFhgRRdHgDHl9fmGa4
NFCKE/NXfgf4XerEiQNZnkHna5asNA9BSiVgLKNhZK+47bcJmRu8jsUSbdKbx7g1
ToXZKGXprgC5EayaCBJxg0uP8NAXhrLBmdcZ6RkR4YFl+N1HYl1mTVtK8uFmW6PB
fWz7d261LUBIwYOhNnNMbDed0/OXh8VNynZaMRGeRmzzPofKJ4QQa6fBRM11pauJ
LwBVR+4RY87PyIzuXqd1TF7De66eMs6L+80w61r4OMnbb0S6oD91jBZFUXRdLL9t
dRIxfdb1VDal5sr/abP+MTWyv696vVGeAwK6pjGSQvYv5yfPU088JkFBw0qKbWYa
Ewm6OJ+sYuFIiswzRNNJiPQMTprecRt4C/roEW7RL6IYQp6q31lODDw81k5A6ugk
HiQHyyClilpfGtwY5lKRP1ddBo7J5C2bbu11RAgNDSVGXHdHoYIbvzGiIndzlBHl
qycOUhcmXgkFEjp1/lJwywdnQiB4cc4kkm0uhUzMGqazA0xhtsqvozS7EVg7lGOh
cbyxf8AjcAremMBlzYT4POhSP/yZyh3gGcBJTG5+tkeKOxFfF6Au+0mwmYO41nPN
ISRsbZYeuBYrwHJabRrZTgUd11QuLkdTcxQKwyBaCaSDTga+OcPJ20GuAO+bcaql
kKLrtDIx+Zu4zsVyRbemyWd4V2cYq0VlyGWjSfau7MKag6dgvg1ba30m7cMLdNBz
MlKZ7Aal0w7ZQMuOilg5j1T5E4viCRt/S9tbrQFeHs7+mNPKt2TZCuXWQe1taEYl
fjCnT4GSPvOI5Dl+FlnUbIZvFkIZ2LTUrqdohE7iIuxuDmhmWd6LG8U0mMQBTg/y
9ILmqpkbUffqDRl8j6ZCskdu3itMMjYDY/4+I/fJY41nX06dX1eMrrPnqvrz2gmS
Mg3D2Kb+De1Mu1SCu56L6zI1vB9V7kqcFfk5AVvV6GQFpyHawEC1aNtg8N+I1GT5
1rLvsOgv7htgQNtF4Wgo9VM0V56Yr2u78lCISXrmACwIpdDe1renhV3Mhcqw/oRt
mw8GzDmLe28H8QG3jmQq3WHKw0J2UIf+dPMk6zqgo91K20aqtSYTpxCBqoTDnSgv
zuS9MlxqnU+pmmbFlogofvd09uysdpcq4dnKOogGj5HPvwyGJkZRQZxZdwJTfIyc
4b82EgCXrgN7I5t0cFFa7XUvW3Nt/Ni2hUym+7iGx02EMzmYTmNzYXTY6S7EffZ1
VCBj1S1GmRMxk109qrYYuNA+cxmjizkI0a7pD9YC54gK2vfxgtD3y/sSr8ku5mNi
16z2JW6VfvS5fqym7yJh7VCs8zG/mYBEZ8YvNjNDngANUSquUvbCauuaLt1WAYcQ
5cZNbT3z+e5dKhPdqZQCu1Zm44yWE3E3q4sGeFchkjDUVZ6nqjJChSUyk3ADdeUX
aqASkdwncnEeA6o29h2W7l6AW8VEGYD1grWVANQ1V70/lZ8HE49+RSk8APw8VS02
322Rx4qlGm/SUNkCDjpoUHD0T3SKTR0FaL2ETs/WiT7TKjaJt7BpECqDHz3/+lvu
Nx5rsWJFpB3gMHNXPnU0KmoLQQWGyo43s+VKzPjMBODuMd6MwVtRKTzT6bI8UM2i
tzFvR1XiMMeU4HyOf+C1EI2kc3ccfjwYtCG0SbVV0UTQy8EL0z6XFTH4DT+6diHO
gCHZcfjBU25P8BfwKQ6QqL3q2sACeDKtSHu3VLwjqlYrrfktg8cXBxyDWRAh7ICP
obgbW2G/FnhCtfeXDTU/nokhgOWvU6PswLyEYUbpj28YaCYjyMB/EvU6cAYP241+
aWt6LeO5VaMG0G1cVZ1zkyLi08hs88NQNIFudl8rdaIujK+pJRmDfYJVVUKWHq7k
GxKrLnZRxFY5rswsLDxBgCTAdiyJinI8iXosxTdRjvqOE5DFwCk4j1RCJlCbycxV
qO6IHmXA94zlRIlMcUZNZYI55syJztyzb05knIJ6qjTR5PHSRGcYS2Zfsr+21TGA
VuCUNuzmeIRdiW/NiIejgFWc7lB60EEnqX4BHpGV2FAJeHwzW8nB07rvS/HEILI4
CdzX38/dkprXvILSXlDKrCKlIpIVy/S0KOWub8mfLjH0tpmVPiqVxRrUIAr6lxaX
WYPD97tBSCAMn4QdumMFfoRXQ4xIqZSnMbBGyA522UjJisJVM635VXk8mLX7KdF/
nqeyRtyVSoi1h2pGUB+KxulpXbJVDEVdw8H10xaCu6lisW4049GkqCzxWSbUwOq5
Upnd9weIeB3g9hZZaiFKixjWjU8Ffoph7tqrznL8JnisYHV9JqwplHyf2ELCUMt+
BG8SCEwteJVv2Lirey4giRUEPYsxqV8BfsS4qaPshKk6NUjiBaoR8TJywryD2q4I
huAwjuglbvJQAqWcl+0cuBDh8pxKOSZ0Ctkti9OM1aTq1CbWsv9FwwqBjZXdBWWw
DYnk8VwYjWEHjzT1sMwWfSm8/6w7DLUZhC+H8ySlX4WiYFuDuI8dY8gv08jjxG1H
PfiFXChdU3e+2YDXrP9APujjSvF397in4rMgHduk7mQ1AfzbKclb4XMILsfVyr69
CXYtjdMgkAmKYb8F/1aKKYd8PIiCTT7uS8nsakMRGqjS4C4PbX0gDJnfMci5xNxH
8f3Cwna9d4kLgeNNd50QPmp9IaE1JD34AOImzBAdUy3qtimpmJr8+k4s0o5PZsVH
K6KYf/2nMQvlOExFrx0r7Ip+1ISSG8ne8AGuqUvRQ6wIH3z1azOXsnSSMBtofHlq
LsgX9EQeH9eqCu3uUtDl5P+lNv+7spNnlmvk/lB2+NwouDQuzlPtuAbIwZQIWnu1
NryaEk162JYMsDAUJZNt3alZ6yBcXEKAbz0y9wK5gMgLvoKyOm9LBIGu14ZoFVAp
4UC7inrv9FLpjEhE/lTZoWJIj6fUu0ZWt/Ty5AxT2QhedWLp9v4Qrj4b2gZ6Bo9+
m5242XX/NRlU5pCUbOCI1qdkE9oYqJVFP79Vkh7HGdhazw1nLDri5WP/t7lNizm5
J3b7KKoK+wfzaCmrFwAOeZdrYr55sIU2yIIbpR8XBfoaYPfBgum/PIMeLss0fg1w
vYEEag8cnHimNbsHrgnlMTvVxGNFbjT2r1ZL/dgK5esoKrgrs0F2e/SD+iD2Ljk9
JwyLg8l3kdnDUfHzgdJGZFhuAtDw36Shxk1DN5PfSc/Isz58uVFz2R9pV/y0NPnP
qOX7dwjJ6mskJYcXUu2/vuFSuY3cLZLE6EQlBpC/u9br9kg2pQblp9w6LqwoqDBp
UIbciEohZ7hTjx2cwUvKJilczgLiL5vDt/YxwYcosMg731gzgQqjk8OeKRsp7M2I
kCHJ1WFv61UbgdGI+QbhUjtbhTpuXkn7eWnAuUWPLHajb8Zuv++R7Ntj6mYlpBI0
hdVuJ+W4uYVMfCJt95w2M5BMCExs/hxZpIo6RsgeubC8NxCcA46xQOyK3nMeNZuI
Y+mQoYyntVqwO/zjTK+M5SKHO9B47JZy5k0/Kyo7rXNS7BbUVH6qeIXnZ2Q7TlMk
Xm5yuuf2DMZwb2UrGJKhFtWoG/RDNm1kf3IlBMtTgKBxjBH5wIxp2+naiOeL2Tuv
gQ58MvEd6RQCBGrTEYnLOs6lH90nbA2IbethOVL4DqZyLKrx2M2/FAUAVQZFaXO6
THvN7nGBhmZ5uhy2iAIgH3ibgjncLl3EhsSS41D97r0AV2tjbSDz7S6avO973jWw
EfU2EoyfISEpMP26Ce4z+PXBZiQ2UkuhrpvrvteTNki7/7Yxygv4poDg6/hpxDoy
I2rMpfGh8nQZBFZGB/LLyJD7ZegfvDCG/hG5syY8PdcReSVMjFS7joc7FpfkHMeI
/Fuj9G9Ml9C2uHbkzFbFD+Ngyg2jXkjmG8TVl3J/3/c+E1UTba74v/RNCiXw54Z3
Z0pcLFaqNjSZ4MSz5ZbPIVlAGn9fLDnzMLJpSP0Ei9SmvAWLx1CABTMdjd4rbB/B
CVLyJC4+BbtVr2kZmMSFI1/fIFik2lpfK8JxzIXrYVKI4LINbjPoAhs2eM0CGC7v
u7rohOrb8R8GOuxS/XJ8ULXtPu70FRtkL5FJqARuZIK2PIm2s22QZk1+7pfMZ2NT
tgz0LyoEuEKty7O2J4u3OBrIuc4XlBgGoPa76Mxv9YCMfiF+QN+afXJR5XEcv1kR
ZFDerKw2GpWP+/6QPVCsKP0G1FrQiaQQlEZ+kOcTHbISiZspqpLA3T6VNp9fBEmq
YB1J0Lis4dsjsmDTyRNaYGOlGutBIfoy49vGIZdOQEbKTx440LS3GWgLh/B18ivt
fiDhpYDxbOvbRZWZ7yraDFBUqSPxrggQm25p5gFDS88rTYlBV1PMw0iEW4XiKEvL
aFadUtDvPv12Cw4UnhhFqBcPC8rxlY4s/r30EInhrpQwn5EtFs2LgEbEpSfyTqBR
y6csdT+p8AB3QGdYp437wO2Bxlih3WEBH90ks79cvtmosRFMFJ/0p0esFZOsFPum
Ms/dnF+5rvrs36jHigdkn7/9T9w0htuGUH6Y1upr4+Ktw6e1wH1ytTMdlZsqkXHf
jU1gBB6gTeWP+e9h5yJE+2qKX1yDwv87KmrsU6tj4Pb712wywonneDqVtq2fuWVM
qNnrK+9zWtf4/I6N1/AU4AWVVokhi10qIQDVuw5+fw/d5ECNSQnezqRABpWmBI6C
euvgMhlCUifEgZ2YTsMqWpX9SNLi7/vqp0VTQUixO8V120PkDt7mLvaaVW4BAsHW
I14aoj9U58i3pcBoMMytQdQCyaeG5e1Z2Ly0ixWZFQZUup/xbwoaYSFWxe68a4qw
sQXLvsM7I/Jbo9QsWr7BH/ZpdHGYFZXjPQBkfrDKZB5vww8YSKk7lQ12X15Yq8EZ
KKv2i42Xemy3/eQnxk1M8Hj5DZ4v7ijaa6iu45rBDILnHhICB2Nx7sCUmir87/nO
xAupOxfUziLjNvT2PouQqxwRhF1PZzLu8cwf7bCGx7fi6wqGSnQD7gD9iPC8gVoM
WMgqufw8TCi52m+YSKut7s9JQ4pqsjXKHYp1Qh9wubJ3o6R+5t/fgCxOdo06gRNz
UOLFokGCroSM2zx8YIrRHNwqLBOEUq0nF1Ow1PelGptVLaK1Y2G+OYZQaN42jII5
LD8iKHbED13UjLcOhOUqKbmKeVN18g7+c0+ggagFUa6QsReAiuUVskEKb7zT49vT
0/lX9hDEFiEEkthIp7YuFPZtXTKCSRmeUxgvTs0r71uSFCz+X+BqP4hYjV4EOI6J
ljrqxNRrNj48yoMl9Cuct74psPifg+GaAzmrf0F6fa429Adb2sJLf7bQZVsdxbsu
qDCZLz0aRZyKq7N09+p2txEPy7d1vjKn+rHxlgRbECOk3MCMkykhT88fwn9QOKAJ
c5uTN60K/DZKjvAQjOhco+47NLZjHomtki/4XuM9SYp/ini6ZqvFlWIxavkdmwyq
NCcefp/cBJHS5+6h+oTaWQRfv7Oe+aFUhBZkB14svBBVEYQGPI7iQ6NfJndNwb/h
A/5byVZ9Uwo1uGaXUB3er/ujbqQjvt84KUBfgtrMy9H2dU2sgg73uKRpvWnIyW5b
gwyhChfj4R9NSPBZA6WnfYFVbLPWrd6QCYK2VXGws4mUnOZ7VkFDBv1/yQ4nw//s
wI5Ay0S7kLffcXuimah2oOEUuRhbdTq7mLB5kiTofX4K9Hm/tfpbh2X7g+vOAQrL
hgB/safoX5x4/YsWWSj1DMkZq9CBKPkLbl5nI1qeXrDM54m9PPLbedZ79A2tSDfn
g74GyJm7z/ikKRIxNhEWgXCk7FAne2n6XfuPy7zMyaaWKoE42awKjtyk8FG49NUP
jjS/5VK+se8sIwpql5BMsAgyyYXKLbnUOXsPcWOw1eohPGT3vCUWu2Xy7O7UoeJG
rdxrN+CYQixPfVY+qiUz8P+R7YiSwYhn/ko421ht6psC89dBTjGtkPC0qqcYAgSm
q2BeTQ9IEJqBc/0D2aIECCOfouDhjbk0ZBrs7fiXID1ggE1uiLnas+9fdMqAuZ3/
2le/sJB4WIqoDcfiQqbO6Xdzd50DlP9nJi7ngKi70jSNNNg/LcddIE6ln6i6yfDJ
5DNw/UzzV/g6hmBqnajFuggxr7X8+IJPHJWsUqljqrlmVZzLs4nXuUvIto/AfTFL
LBAlJgB3orhWc953B6h0CzAw82dT3G6hFUHya3CnhztLrLToc0N73WKCg+D3pO4s
93PNozDHUwvZyTrGa8DFYF8npcoo3Usmq90h3YCd9wU8IT016V9yzin+4xCeaXn4
efeoM8XKI0Raa4EChYe70/qLhojtaStLSRFsuntEy+RBwbx1WbsqB6F9WbsTGglH
CT7ls9y/i3B/dzvVNovOrkDYeEZ7fVwTgrb2Nfww9PWnbn/fNwb7JSnNuZPawPLk
zr9F4vLLRdE4kOOvwxAHf8JOQFwOYAa8XXoJJBIh+ibrUIVtC+f3A73G6CtZbuYd
jseVuOUH5booxUqgMoHAXWntdksvk7IU1JxyCiE2cUGyC57dU+ScoDU11qT7bay3
AOoORSsekP6NLMQYhk1awyrfl2NyjxmwjVxs4bTRfCVyPFcpZS0797Vd2zbvt/Xe
FhiyxnOf+GIilBviw4UlOePDqeg2V3FCFBUnJcZwJrRjk7mmc35whPAXa3veo9gg
Kuucdpr8bIDutUzeEVuABg4f7lZvpXMTeXhyhS18Px5fZVrFcxNbtK24pVVr2HAp
rfUuSFX7ryFvJRY+9t5NOEHFP8VW2AAANEyktC2mRTbW3T9zs84TxCdcRO560s49
dhhdwQYzpXSe8X6/Ea+BKJSaRmEThltrwEvSCSuSANcgtu3UZPo4Qm3w2xf9tvd9
xfmD6KzB+QbbWmBX0NQZgP5hmi6sK6R/XftORFBLZibnTD3rOc4hTJ78clVXkwr6
O4oa0V9H2M32482mlBjcNwibaT/rG+089MC87TZ9gvNc/XFwLhn5swCFD66jLMRh
ceZJ4BkRw6eiuSUuk9E/eOWWz3YQ/mgxZjIoxbGvYtgdE6EzEyKX+YwpB0JC7RSc
aQIwWcLRjK/RJh6MamICvsvGdfxeNxN82/JTb+FpIBY5aLWvjBq/HMXtyjLxWcos
vDA4EICaK2zig0u0BrPtCQLWtSRnHoy2RrUG04kDKlXqPa6PpTYVjMcbPq0/9pG3
K2duF9OR5PbpQqs+ohGBT/mu+tDcC5WxqqHn+bSY27oQwsKdMdcWZu5jgxrwm9Z7
JQJf6bA7QecOHjvKK6AufZKNPQfSg37G+uEYV6LHx4tKlxzqKmLSthBfVdTVIm5c
NTnI8XhmDnvY1aI9bKvAxTIRfY/0/0GYx5tQdQXYVZhHxrRuILKacrvm5DfDUHtO
ePHt/UIPOn2E3l6XTfkSGJa/mHwfFd59+6h/uJ8MnPj+nw8qLsyFD/TW2Q9uva9q
ha3v4iU1dgHFarBNb7J130ift1l/teV/usuJuXmI5rjRHwnnjLtZKhyq3WA1O5jq
OEOVUKk0qarAhZx4d2g5pfn55vOe5waRy5IeAoyuFsWoX2Ilatg1m+glDt3/93Ow
BFw0ABuMtslahmbu56JQHRtY3izlske+8r/IrVpAftxhGA4ZOid0q8jk0CyNcVBv
R3/Sh6fjB/xpXfTXnGsD+wx06oHg9d+eD5ti49m1Pi1edkX8JGJ2SkUSCBn5XTqi
dvdfPi8DOkJ7LZ3BEnkynrcSKUUdEg6VAM3ttfnpheTz1ji9oXSk4gL7Fh3vmYrx
9OZaj1mzOVubUY8G4fQ6EaJI3HETjQ9XFyz/zK8iq7eTEjZ9oh78lUuXLDbR7iNq
OMLC/HG3PqNQ3o8ZWjGJ2RIntXw+bphyxC0jN6z2T9iTLX+ZneQhFTp8BBg8Pojm
4QnXpGeqWtnWjjMLJ5U1EzpStsRfg9OcyeqkTYrFqBH1fUops/sVIp9gspaHBEPg
zG1NWYTRKTh7Cr86j43Z9Wf6xjP7hlKwxTfbuGrLyQEsDA8h7KCFLI9gGmmS8Q1H
nqBvw08DHShON8Wy7ZXPVxEU7weR0TUIISvwa9zahQHZ1risyVlF+d0f2RWMv25Z
Evod4mnUTrKAXIxlCx91rb+JjKLsRjAvqhJkdxGdkQdWYa7PBGci1pKl+ilgxzcc
/SwbU4Ur5JezX208ctMRFlDkDoRs1SPjm9iLeC8qQMSIY5ipPrY1t+WSIKbj+Qyd
wxme29b2JTTHhfvJJfLWmyzhJ3dZFoRVhTFietx3utHNVqG6aOKyBw008Qt1/CDP
dolDsdEN65dmd8s3HjfFLbaDGjkfRUc0Oby4Sjr5nSyu1S9PcvIimk+qTfWIQ29y
IPaz5RlOl77Bp1nIMX++O6ecNoGLwRr81hMPvwmoRXcuT/hNRblM43mZOPTp4ufo
xgrnlY336POGj+LUtREHiq0eKRkxCkVLhrt7lWwOXUH1qQlqCjjm+8rr6UEqaczs
swH9gjXQLmnmLgQF2HSdwVgiasTSLHVz9ti2/b/mmouBkGjUXDMyPiub5ATva9t8
lnZaiRuu2nqGTUwAAWoN3jsX1K7/CTMd3wOtGQqWUhy8Oi+d0fKcycrFDyzCWcDA
pcRn5nTWic6GBJfoZivp9X7jNOG3+BvUpde/XAA/dgQPwagIYDAZKPXC7s38Ufu/
jNJ+HAvTBt8YZJt+7+fldfE5sy3oX+P3JtZozR/sP2bcMQHEE52H+FDdY/1rokYu
iSiy45hupILdKU3o2q8aqPA0g3YqQ/lE1hNh3/rIt4HduJIz7nyUAXTHNI0JPram
0aWgylZ6qOVXfhK5UOQqKLy0X1xfgiNGaWCc8cfvnPxbmT4ou0bwvXifMAvsO5Bn
EnkJE9y+gtqe4VYc7Viejoj89+VxPN8dx2/2FLm/Jpms4YlfGun5f+2PbeDQwyQU
+aEpkasvmvMtcGRq2O0xnBQHy8Ama2UQl3vT1+iSRhOdbti+lkkQK2McRnlZ709l
hJ09PUzzcRUaTAVm4OsxlX+Ewn8Vu38Ozu5SoS+Ho4P8Q2ZexJNdAkpVR7L0GYj/
tmKg6TRUX97jTBeqLnBXMD8d39eTMQz/zldUaghm14HIbzzMzKV/pbQA9w3igGXK
BiD7cjCz1GmeTU9X0aZ9iiSpR4Bueel533TMFXY4j5+eJf74kBvgEbuQK8LOPRgC
usykPi+Xa6DWGphpZQ1RJZ4Bvygs/StPzce89F0SBsBdEjG4v7bKEa9rljacxZhV
I8EWKsSMcLBIrrSu06hK30Jmo83IDXUXRK6Vj7CD3yOwQ1HE4mQtacN4IfHHJhcs
05+tb9JrlGO77tIP4wwAnoSg1xbBNnk1ZGBlPSkxfYWnN7mvAitf2cnvtrdGLLt2
jlJUTSk/05NToOfB78DKPQzNchULjXkyyN8vN5IR1SfvZKvl4jpR3xEVtL8B9Fi+
kKAiDCsghu6h4fu6bQQDB6wYCP+ytfkpgMnXnt89GUMlL4I4TH47L3AVI8brzRs0
p9o/53/cHIQOLQ7aCW0wrYRmKe0292IfBmlgHFm/gojDGX5t2kY7/gAQh6DZCez3
pzHFrZGrXH4ko6WxSDcQZuvHN9hba/jnHez3D1oTZdHxfbz7OyxtoNE3ln0N3YR/
sRjeAVWQXMsHCL/QOPuC6k8PinXPJEoD9HkZi2+iOiqUoK1AXfYsXl2YdaSk6gjv
RKwiUqVe3JFnS6Dz7Pz5EcBFhtMRjtJHp5b+kKPc1gmGubDSJs2eOC3eHgt902Bp
sAOyVqgvMWpnjFpfot3KdzkKRyJQrVC7GiMsC2Gujiv2KtAjQVQKyNA2R2dHNJpJ
+kvJGikfnLGPqx5S/4Qkc15PIAoPcRHDGPL0dGHEkB3HAusQmuxWz/wEPmwbszlJ
Z+76Bye2uVAbWyX5/ATSdeXub5VvZbF6UXC2KSyUYerwbGAoRSbRmgGwVPJ+zcUw
3PuHmBLXW7BoZVXyocUt0UJ0ifqQVYgtZs+mdxmcRoJ7PntwPqjaDfW/xtTus5Te
MlvERddw+8OQ7u2xSLoPpcT/3bbtuJg584JtOyv54UltJ57PKY3F838DUs31hAkD
OY+018H/zmEeYEl0IOLazSQbnaG143Cfo2wA7q9YYoc1u9toI1pE3P7TiZKxs/kP
UzK24vczL9prqFvw7HQG0tTFhYoEC6y5pfT9iIjyn2ARSw/GTYcSgO7CljJnsSHj
zSM4uMWOBqGhL+u83fMTM6+EsqlcSOh1dehINU5UjnR453IIIjhO6P+9bT/DcCUT
BgdyISjQvHcAST44D0uqgZ8HlRXKFfmC/9Jgs8VDjBDFK4XPa3i6rCcj6mKuSCIv
Z+w7LLvNP+JueZkX8xMuOZ7YRt58hkhbVNZQtd8UvHlsI6ynvUMZ2K37vbhsj5yS
rBU0AjGSJE8acSudNLwtiAUCbzVfMalXiDGHFYIyYE8xM/Y0f++S15VCZt5lFbZG
8J2MBNQrA+JeueCjrHECbKTAEG1myCu1s4WnCTk5psbES3ejAjztNxxTEwtKupGm
OCkK/LRhG2uEZiRlx1EuoC+twnIa8MwF9LpsUonUX85rZwx3LfPeL2DBol2p8WNl
bRLyTyOzGPndMJox/gp4ZrKJDvf1QlNMQF675IuchDRaczSLX+2rrLpdpLcB/Wmx
9+Vd3a5lwFkMoDV56AMZl/cbjKQ5rybrTZAsOQpUMkyTe9OXwkuR6iPbBB2QH+Gv
Qj05/Gu6gliSeEri0FCEm73QAcYlFA7L6emcTQygCy0xKrhED0FbYVGa5jKKRKfV
bwJwS9aK1q4/CzXri00U0EwABBJZMS93BxA8CRrH4ZdPssf9xPbPKwMpew+mKQ14
zuPrIiu1Ys3E+agW3ngu4X7fobMnDQBxQ7txwJkDfhC0zl7VKnJIUyECGsxoKzOF
yw9C1J0hsK1b2l96PyMdf8hXaMFWbcZjo7YyJstlKl8yIIFqOjQYFikRV0dkI7lp
cRNV+9QfuzICOuFqhSoHaIm+4RJX4mOs8kzLqw6p6cBGmsxg4cY/FaAzeow2pqLf
0NfQRzKgfnX2j27xvaf09IQcsUjyOUKX5OzHPUn1MS/Xc3mQd0dTAqgc8NVES1OP
mc+o20Scp0Y/QM9b9f9kjym6Pt36gqgBJjT30HpNzguMtc5zkc6ewdN5pYCd6fEQ
8kPu++dK82mXuWcReR+CoaBD99AZ8jVTh8ChKT9v1VMOSLWiyG1NCpzTRSm62t+I
DIWWKvcu/Sn46iQ5cjKveoQRuF2sZxVhouKP++aD0u+D/m1uxK9+e+1F2P8uHNjd
51bLKfWF/lH7auQR8L7tpdmhOtQ4rtTNKiR3SRLlELimFtavnAqd5IHNyD++uclp
wfxH+OycHEQT4jf4R54QCQIv+AnQbOPm0f06xn4cY12kxAH5BlaFp2/c7n6AFIl/
OKJREj5VnGQo9ftOUyttCUxS/YpuiJmLUEGwcpv0m+93CTfAfFBLF5E4VYk2E2Y2
Y6wre9IC0sP7Eir+/DooFZ2ORrIv/SEC5Ddqh0deQcIQv0Z4LhbP0Hzm+kfPO75S
h6MzV7155118oCd18B9wYfhI4HXBXrD5RHzSl9hYP3Y/d4e9VFtY1v4X4IQ/cEML
7Bcg9Yr51sVYgbTKyoHv3WoDv9kR0NqEmJGz6IU1/Ot5rkHRxQ+jXqy2r3twFFa2
vSRNdaL/gAkqEkYsRebPHvmlClUvnczSWSeeL6Q30wR34snKn839z3PzQQKB3C1g
4w3BUM25PGZm5NIzNZkis2aHZS29Lix53nN3kegP4JS4uW0eIevnMXEm/m/HZbww
IjHF4kp8QM6gYk5MGkiH/AbW7p2r+mu7KS3BG7aV0ETeDFn04mesF/3FWvruCK/D
omyzwpQz8q00Aic1tNUYx5KaEbohw0WW0sWzz0kcxO91Dnw0cto25iidEFtx0lw3
mAe5qvSfuOJDPng41L2XNdps60qSC7pxWjq+2K9GexnOTVNvE6hF7E72ahMbFrKV
S614Um89Z65+LW30I5gOzBflbYiPS9oPVJwoP8PlS9ccGKZVlup426sKM80h85NX
BQ5ExHdNM0y8pqoahBURGC6u9uEIgrPpTs9FsrVdm1cNdCP6H1H1A8wtxG60CW+q
0HfI2TUi/9OURib5wQc3Y+FmBBBGZCtlxWop4XwIk0BnD8e5MVYQeoNiQvgu2F/C
6SFex+X3UGSR2I3UfJw5dWTDUp0Sk+Qs9JznfuyHP7V2gnaP6j+KrH7w+QjV2F4r
PqbcrXtJJ0dChwHNOa1WlsXcCTSWymmgYJG/pLvltVDVTgTp9nzokgatyGRxCSga
MpwkDHiMhwsjAgurt8WJ1fuR43pIagTlC4lMkg6mQ4Dlf7UADaD7UybnPtbFH091
JflA9VwMM6MAh/XCPHZQX9qgaGwR6m+RyeyMt+T5zX8/fje/E6sAshF+QXkH5QxL
PmALe2uo/eMg5EA1KNgf1mjq4BzJ1Kw8F4YIr7s6gQtgSexkOUuLZM0wCbHECwLf
FpzFW/6OfWr2Wv057N9cJ2K5tvYYCD5f02KzvyhXaIjmf4X9E3W+jxMkO32AH9sG
GRb5rrqGIn9wdP1/9qaOhFSJ0gCI3RG/tMJ9Qn3A/Z4TwM9QjAPnBKQYzkG+Pcz8
uFwKmtMiRDb73Qhr5RCoXh0E7krrWUVIpqhfy0p6KO/g/fwQ7fCIxd8ZWI/fb6i0
bGArtaWliWl1GZvsG9NfSJnXBab0r+/r+TmOcafZ1kb6lutLrktTs0QyjDwwwX88
K1nlr9Mpu6Lw17FUMv8/2RSTQOpXLqyLwxjBYnqLjlNYAov8xbyls6wHvOYUtMcT
xIVfoVnL+PCQGwcqmJcUlxoUWMQ9be9J0Vl7rlPs09yFZRi7YQnSgqNfRMpd7+fY
C8kUIAzGdyIsFSN8305h3pK7c28X/ao58gNeqPUjQXxWWQEhlT6lDTjS0Ninrouy
0htEL/XkAkb54YzaVbiYVFZcE21FaHIDBtWdZ5oCra1J4isB+uuC34Dq2zuY+Mf1
HzSrBZ4ymXfXHgPO0ueDhrrlegoFBWOBg/DS5FU29JPXASvqNQPB0BYgkkKggxdD
IGJ3YymuLEahWfJybgHix5A2xY0RjJgi1uwx6SkcbKk6bmf3PWBQHqBnKvCf5810
6u8UcqN4RGa00wIJQf5KRtO7/57kBfxlUPy37QE0JnEFQ6FzxCKzE0WPlMrpYia8
gR8csL68OsDAoIvFlFi9KWibhDOEN+rClBZRJzCLkA0qtYG0JmLinegUYJBLteEq
gFvlrz9sjPfxhDAliStqyDokRhq3U+53Lk62bBjgCjiygxHPknEluzzQ6jctj8H9
LYVY440lL3nvOsuUTH5mtYy4mttVyL6iNp/DA5seQvAh9D/ag6LXPSiOppRxSvkC
yWOqVujy7VBW7idvEgELQwUwAGSdPUvaIGm+vxLjK7rE2hCH2sQvRfEcD90pTXle
PI0NsPg5rq6h95qbhDUCbdYBKe2wwbrO5vhb7ojOZZ67TE89++OUdc1V+FkhQGIK
XngagS4ysoDNVDOM0Rfj/U9gB922PBD9ZBdOLZ6qoTnmtjYkpD12TRVN+Tn4yG++
+UJftt4j9EpOEGZuIxmoowZUGhBwU8ztPzubQrnDT6Jo5gofxz1LsdGzB5swaXCV
0Op84zXZaz7nbyv4Tq5FHG2ewt4ddPL+U84NeBUKziVkMf0nUwa+HmnZpxxEUZUe
HgdOPglvxzGT2aGyRtL3wbyJmq3wRbqmigqSTuHchb6PN6mQf3Qgd2MjPv+GxY82
eJYiVkkHiTeR9/vNj86zpKnlr6j4cDIw/Vubl5CAzetoqR7pHL7wNq1sWXThTQfS
cuSpYOwvhT5j4I/uKeWJMyo+xiKu/kBacjOlmYlSXM7SpkX6uhYYh9cX4pxb+XhU
xpfcWmRxjsyZR5czSt7+NaIKjkoekUSfyc5OgA1LdK/44DkV4EhqzGrXpKryyrf5
9BwzUu+jADZmfT0pc/zTFqnPpvgj/rr4ZaoIKJ8FXAoPK70vdwQ4ur4spmkWaF44
rhTKB+1UeHxVWMGYpXAW5QIIMHQit2jTlPxQb6oZT20lTCfqg6kA9CyKfxOrY9VI
CPki4izhAEugzSxNZDBJVLEsA03oCQrkTRdPhaOyl1PEn/MIE/zYyLm1wixxIwGV
RKMx/DAgf+dPA9R7zOkDbUMm86KENJUylsNQRcg0uZni+UZ48eNjGp9w8q/RTzk5
Hte/I0vKZGC48teca1UCf4+jkGtil8BgAvE1HVunzQL5ukrgHrhYr62duNWffzkU
FIkFAF/gpq11ho/XFzvx7hYJZpjB7YcXb/j5B3XHX+Z/KluyxKD0mI7n2PPm6hiQ
2T76q7Jbpb27kbs91KWu/6VTGLb0ofKz5NfEZPsOmwLZboDngrOxmvvGS9Uy0Nmy
vjbHY4bUDij5bdgFq51xWJbB/sGAIdtK/Hubuq56sjn/O1oRmIV7dnMi2+/blebl
3/GalxLf9QBIZ7XnfoelGN67cup449bmKgUtMX63DRkJz08OR3hXLTFda209cz40
hNAeGQdlGXRkiErRGiymnmydc7+PQT9deOAxgIJ7whgcwdIpePKkWsq+LUobw85R
1uYo0QijgEJChf2extCsLBnU54O38fTQmi4pzumr6PrXMAkRlbbXgejiI+KFTu+3
/hkc8sH9zGhAxNMmgzGY3MhQcDQsJGAh3eg7Vs7qUwE3Wio5tPZTb8vPlomL9NZ6
HQdQoUXI60eS0n/xbI8brIwtVPiMA8MdSwenFrjOoKc171GZFcD6qqxXh4h391sQ
Zfb6TjAWc3HF1s5UAZePrVIsEtiOH3RiyCKE95y6Aw5os88CXO7to8dBYwj4nD87
01Dfq3tGQvMedISQN9aKPZ0IAtGPrqrF8e7ggtPqcT1A2TDvK03YO01JDPOnHXhF
8fs5Jvmc6DePlpxwo58w++Kg7eLikuIQib024aQyIw/R/tKkuKxMjn9uKEDJ7zLc
e+HhYcVJxVhso0joSSvllNLtEAyn1ea4FkaPWugIg6W+BtP5sEZ3DIio1UzdRwWm
UJ2cb+2AAWk6Bc+Abv31gcjCYosXuXHQYNgOeKRKCkPVB+jbVd5CLYHMogOA4jbQ
w2lZr83mFa4GAz4Eoyhllhbccj+8CKdwhhKUNXux4bgyQ+QGmYDNDFESWl92rdzC
1POgiRnPATXfZsykcIs+qAd2ZhfPKMFUHDTTOe75RX75mjtM53evNoIxI0rIpIjg
aTlg9ZwD7PZhsxAwQKKQoWvgKedno1kxwF3Bxzvc7QZ1HbX4rElqEVfXzvoZwq0x
3hiY3IWJWlyc3iTjXTPoIB7VRLmwp+K/Lz+aYwph+bRIs1rCELMs6r3OcPJc+c5L
S8ZJY9BdyzYVXoTHEUlwXG1E9Dsawbsi3SyFH2jOHsNyN42OL6OT5QUuukupbbvZ
tgJ/f93ARGEtIeAcXsCdNVN2YPh7m/pYZMweq8sQ50wbDPUnLV6KRSHAESaU1y3A
MixeAXhEnnAL7ckoLdGeQVOK6vu58yGZtXSEHg6Xw+5z4Q5ghTrQUYxLG+vPo7nQ
ay2VyXZVoMGwI6N82Z7dBMAufjyOoWN507SVLmlcn1DhddsW1CMI/q55cTNxU/m1
RkxScRXFIt0BYrq3NC0r/I8sPWdGe36q9SgAubWngNiMiY2HM1cmJm6AWwBIJTcN
iEcQkrIitHomBIz8UwxArE/On0JY+WFjDr/PNRX2vLlN9wgJO2C/9VtRKRnC0ioq
bsrfyUZw9rNn0szaAGbSUo1e54eGPBA7qVrZqpPBMBt0siSc/m60bNYf3SBdfv09
JHJS0KsMCaX2MttRl/fhom/E50PqGBVro6FqoOFR6Nl6xkABYkJ2sOTtGeYS1fir
FhOvxyVGP5K0sKetNkos4Kp9hJBzw07w2bwJUMoECJrAq3BcRNLHC8lIZalzdDYe
V5mnpUieNvaEUSIIQvEg2CSTJJUTN62CcNgGi6L3MTLeJK2FiUN3xdD+P00UqBDD
8a17lFTNU4OuH2ZRBiGACeYQpIQMI+wwMXGAvBOgWBY4BU8vtELQ+5guEOngqhed
Oa7zSdpKyPsUqcI1/6y7cMRhEboBjaAqb0MfKXiesHHh5aja1hwcO+2VfyKtgod+
CoZ344NNPGPN+pcb2fBtryvXh9duz1idL6HTtbrqKigcL581EFelyoey/JXmdhcn
hfbnprcVXdCszBH3qOaufVyHJznjoQ+a5dH76I4VJ5oZgJJQrqbRAi2GjQn5mX/u
Ts6kFoT0WzJfQJlZ2SFlubRypPl/a0xIWUaceWIpNTPQtJwo7Nmo8snhl86Uj8fA
rmJp1rYcEfyKTk6zvXlj+CJsIkMZn7WU5p8ssPMRCQGq26O8yCnGtYG+U7q1ExjY
xZfo+yOw2gDveDQs2vfGXUX4zj0GQjU4/OR+zFMvg0E/3XDYhV69B3mmY3mtc6c4
GSH9MnSqwWPOnB6IM8MCm6fhxY8KoPdtocHjk128EFO5Wdc2HQCVhg1jfg2DJOpo
d4dxTBbS0ZpNzw8OU0r9UFbu7LbOmhczFLnb7Rz+H2HE5Koxnx2ZK7fy33pfhrvB
yqOXWB5Jf2W04REM1hursROyAXg/vV4jaR91DPTjgJzxbjEthTDw/hZs+vqRsIEp
WO4rxr6Jdk6XWo5ySqduCC9jn1pNQePUhUOZYOTfK/2b0wj8RuizIL3yUceCosnw
Zc4LkZFvx+FCevU8GDwCav77Pbcd5pdNscD4gzrCZrzXgF2k3hLUzo5mJaaSa8/i
1khGv/8Z6t94vi8wlxccdeNipGKvArCzMxQob2XqPaIrgOZ0PvqKTj1iWGg10zWT
9Qj7Dj3T5MRdaZxlZOsdPAEvdUeOZe84HJ+5LofkkADEOHaGqJEwWyolcWA9zmor
js7rM3AZccbFHQQkRTrChBTKCSh8QaatUF0DMotnsabYdWI/JCyWNyPnYpuD1lnF
46ldNoMYoLzPDoDUynq6fyTZyQzReJ2X3P+Q6u4ipxFpZtSQKJg3SVFcYwzDTRKs
EBcStW5D/XamBRqzldIQuTj45IT/NzlMSDO7xULjL/BTV8p6LOzKyGCBAFhoLOjn
7M9QNoqeSiFHkdkOekc5HWmHZjctVL8M7JpLIfs8qlYbPR43LrrNSG1hUCYEssiW
XU1TUOYCn9TMW+RKsrQ/XtAMe1b8wHpFr9nWT24iYJb8BmGYU6iIcFv/hUixMqRh
doOWKkQVwi2SK7B3rBQVoWzsB079P4hhM2iku3RYkklDVre03ef1u+chyJ4eGLKr
c2d/D1r7LoiFlgZiQ6ndrgYr0ZqtnsFK5Tgk8UHkijTnbpqvgeMKOskbxTx9SZmQ
2SEW8MsItBfLYssT31z2iG2R1eXY0Xfy+zx6TQrw1HhF6KvqbF0dCShsb0sDGLv0
7cs2ZuSmBEqE267JyinmEbMjflNzuMWA+o6qbQaQYT4UUINbJEqqjFMG3ybSXk8R
ENKllpzsLudLFZ2Dhh0pxp2gClSsl0XnnLPkLaKdA4SigsagRAwEEXCD8zplPuQ+
9oc/sF5/2Bq8G6gDkUT+S0HpjPANX0BPWitCzuDvmNZqZmVHXRsZXCMltY2hDHNg
IlXbtCNZv2ekJyfYMxvqFOcDqgROU57r/qq7QYlR2ubEudGf9Cugc3JVl6+QKPuc
rzpeKO6jIQaAG+CFQbs7iTqwuQR8xNFeiGCXDEYNF4naS7h10g1q85R1Citi0qXP
bZTF/bDi7Fz5k0rlnSvZDyCkXzTZGxc7yKeF90ql13bOnVe0FGNPdZNZ/fua8C0J
sfgdVzERyyuQA2+D7/Z7fHSPWi2C3AVQG4YCBByNqpK6+6+SwzErI9bXxzojTpXb
bGgeNANJeRQAYIqsAp7fq/HmqC1xmblHNxlHmK7teaiFeT60KYgXGnFX8h7QoDUl
yRuEvEXsVtg30Z7t/Rveh+k0q7kDb1w0B9iDS5m1Rn8ckaaDzZj4k27V3NYCmSPr
+g2vrYK5iWlAOVin5SmbWVnU08n5Yoo2/chtQ1Ofn2I8UYfPJgZinRIEOoTJOMfo
krWaj1u7i8wWv+ciunfSrMnrtK8Cy3LyF7dlmS3SNkW7q26ifj4+cPSpjFNRXLfS
ASxuDo1vtnE80SvNXGpJ5FUHhcLaGeMYmHQaIyxn4wW7iU8KlojZVh5pQEnDla5B
RP8DIs+1/6t1xw2ZC2w1wfunXUQF6dcP7+w2MMRfU6xw3pL6CvgN6snbZad1twB0
QyQi6YhiEBHP7KTPKlEqUWJx69lMDlneOAI0FvJeX41P323d3R8nS+3RIO2YU3GY
2LG2jR44MZcIsykZGjwcFDwjQbK7cMQt2qHs6vMST5VeRgRMwemNRsosAQWsDVJa
isk0Pa1rtwIqbLD196GvnJE6sGUO2Q7kNzFzaOvRdFQKjblGeXSa8LHd11k+ccJ7
vK6nIkYsLNVYKUobD09i3jmHYcvaWkZeyQmHuuOyQ48JhlqKaPyhBF53/Jdt4WBd
O86eS3Bkt4wu3znW/hcZHnpzxSVrDES/AEgM21V9Rsg/ITOjD5VOhBZvnIB6+Ru8
5q802RP0LNguxY06Ysg2YadG/lNN2+kF+Nwjr4/tMpKq+ctWS0jdmy9Qc8hMX+Oh
KXOcHbKGUgq3RcDOBS4sU2Foew1Za0lwCirsa2xuJmrV+QJgVAxafVOXii6kLmGL
z1kjSjP6kCARQ1KBUhjgmgEIPcUUmp5w8AY44VaZV9RYcCaRR9XNZuh1A3OL29zg
OnF6OyeGccYhZQwjMkYyH2o0Ymrz3kRUnNDJhsRQEkfOWeGhWWc8ZOhAFyJt99rh
+uUqHRkWIDsSzjYRMMT3XGV4jsORIW5/FXOUPFUDwQdu4SrrLd3jRWlRQLqZMSnA
sUZ6ElLxb0hp5UBQbMkChojBuNnrT7HHOH1PsjtY8GwZrZh1U3VbH0ZWtjlgHrUP
bziAySL96SQdlPPwnCgdf3KIj9PZyIgXhp5DKwGlMcX7e10tQ0a7NpS5xk/QInnZ
9brruUboak4FIWGyQ5gcpo5KR4MpONW28l7ve2r1h9NQWCQNvtIckCe3H0snpSH8
z0wo2qBwFZ9Iw6gWpd90h4DeSH/CqI7ENM46QK6T9LHpW1gAihhYlTpBEIS4Ri0L
Wz9MtipAsfEm6JwC9p+fs89XyHF0BfF3KP3NljUqkH56/BriBBLYouP3XiXCLfvf
QorGPyQne1YzaQyxd8xORC55ZZcidbSUppiZIABAG2+q6///PP3JHhVa8+7i2UiR
n5hep/FXzrDeEML2TsMEsKcX2LMExP5BB16/tB0VYuI1dL8tZQB4qh4VrVLnhlUP
75eu98+CJe9Ar6Ktc4+o4VQnN9F4SA+CDnjJ5UCdNt64cc9DL2XrNJAqlu6z4uOh
p9T1OUehq8IBmq+301V5oILUXS+5I+Gn+orPn9k9QuzfZunzbAJoa9b3h9Fyabvt
oLG21ELw1r6H+cOOrnLls8vKksRdIMXM81HLEpg2t+77dZ2gnOtL923OwmnmL3tA
GqmoWiTml7u3Z6rgE6mXlKXsQFjTFAViP3V+qcsjP0bKiLAVgR9hnTFegT1m4C7H
hdcBEvIq0+09zixKkwz6IxPaTqrh4vj9i5lD9AAmXm8qa3SQChlOMCCjRXMXzU8i
vlAqIx+v3iLG8G+PmrlZkWoPgQbs3afBPwt2i4JQA0QVFEjLuMgVMODA6yzIk31V
lBTNQmSZpzAMXicgy33E9eBum6AmVkn9HOmHe++OFjqQXh8SD1O3jZ5q9DbMOBML
WudCprvbK9+VEYX0mpT/IifurEAJhz+zhygoanx4FeGnf1aGpU+xeSw5zH9F8mvI
gtbNyG7h+oFs497YbgqvErq0FAGT+atPRE7UOOH4oaUMk/UYy6EuHbFsXM7Ce4Fw
VlFOtpJN/NncCQKd2ZGx/LOZDoTDwvNfjL++AsXHAGfZjm7bUG2KBwktSi4eG7rk
Ty8xR4aGDubx2qvfaPWrFm+H90QNvSJI05IV9mpvGKzAoEdi7ipfMGDR0uu/CrFh
RpGwPxO+uPzqzhi7YfeBVDtCSNaqSRb8uqRFvHvj2YDyCK5e4ZOERNAwKVByU3cF
zzk8q0UECzM8o9ihoOOveRhTI4C6ccBszkC88NPYZO8sEVNA1KEbo5WjWeCnh8YI
D0rpYatn0aMWTca0uDHb8/TuSNDCcxuM9IlBDikPQWEe4yU3Jhae2366p0jhiKwb
bNUYHE7Ya8EEV5cO5oecCgijezo5xAproBA/4hlOaM7u3d+yXWxo40iSKCWHeQ5q
/8qMMAPUgS6S6hAP4ndVYZiA+UJ8NwUu0plvG68K1HuYUz87L+gD+VVl9bmPPI/X
6R6jGiHJlobC3lYQ/8fG5kIySlV/qNHEAlndNY316m1/nFLhGWdMXSYcP7o+n9vC
dRyegtBznriHV2gATajNRDPUglxHeqESYuF70mke4zytO0NLDcMpOvpsBUjZD3Fa
lO1vbBSC5Euet8cFTNxlFlBwiNAg0tsYKDMbg6roVc11bOBDU47c12/FVaoWdSvq
M0XekAJzyM8mU1dS6csYYE0U1fOERIH0HTKbm8o0ed53FsfPhVDQ5apsfX1Gq1KF
0cDc+QTvWy7fVt0Phuh7HYfsQlIIJEDoIuraclr4kaIzw0xTbBVLYdjFMmxsFLP3
vtIcw6Lfa0pdwTj4yYB3TObX9rEDGLPQPe1sgxsdSseJ3nP/o8e8q/WcGjC+hQXU
akpHhafvqicq1YB+GPKfg6w1eWdyw3j8VcCDl1B7VICim8preDfmDu5f6BhwKREo
sEb4x7hFJPWG6kEWoBewhnNQtMyJHREqGAW3idG87sq9baLdcTGbBTW4pXdbZYSI
gAWIUBAQNPlmhg1+knVgaYGID2Cwok+pT6AuJPJER9xYBGDBibJ/UjUWPd1GX0J8
anBJuD22fzP0nuX4uFUm31qczRuxg5uCqhFH+ViQDGiGTHlWy+s+eUfuzaeljk3e
gkOFUNRxuhKfnPwvZ2rRMbotQvQ5qncsbI6M4Ik6lY+0AA6u2Tp5DkN83bmdlgeG
QseNNEGG8Xk27KUwqDorkNDCw95Eo26tzoQPAV84fx/Ti9QvQFNm7eCkompAILSg
OT1gEvjVQKchnCYR6GnI6Zmz1PUUu7zKZwQ5pLHfQ3ium10gFcBIAemnhrs9FPZI
oaDqs8eLxJZ8fg1uOzt5eexcRQeHJkoGVPE2T3ndHp/FPthKLIv+RUN+HV51YQUo
Ep7EbkFoJcryin9ULxON5Xs4BUs6xexmEt9Ek1i7GcFTgXmsiC+kAQHb20Qz5fjF
35KcznRDHc9Kvyblp6v8Wf4XALh05iMkob0ZCrh50krGKsZX5vod3ehksHlM1Sh7
5BRhr9gczZDoHQEaBNJ7xIFa3H0m6jOnlDu0Rra8+0ccynfH9rdJH/C3vEcQSkLb
bJlb5BKPFK9LwEPK/x/e5SANOR1zy9VWvAEKYTqjfGXX9jlI2N5wHAerysu/HJe8
D2mXjEf0d0W7QqYH1MD1yT/ct9bZXp8/P7eGdqyUDZAVvtnYCnq1vAGt0/apMfSW
MNNpwEJ5Hvb0XlB4I7ifipjdGEE5ZwWhHwd9ZpbyN+UVAq8IyWsBOg7JVjYUcGiu
he3bI/RibytLlpUDTgtCoElEHY4EkyfImpFgvsqhoPaAV2+5RUZxHHcPT/T95g7/
8Kji2e62N1S2jGue4bBpXiIC4NBrTi37R4Gh5X5SM5DzdDCCjHOSfU2Gjti1Mkrg
mVbdo8Riv4RQfMy0kJPIgh56DZI0GHN3j5XNEA0FBeFx3qaen6ohu1J7eDqlGpPQ
Zu0Gu48Fi75dpEv3Ej+uvfq8a6L/c5GvH1zTMtxV081GAh4+BggrMItG0H/QrdhJ
rEf99v+dFlYfgXWe3ihKOJ+AsFxzszwPAytOix0QzVrFc/UvrMDzRadFHQuJKFKm
TU6NJzx8y2XqADYorpS3oZI2IK4aik3fBK92LHX+Nck05JNxX8bCwRSqZyNg8IQY
vfQPLngcAtC3RWeuglOrDRXipsxa6uOPNePp/lVmeTppx21xawzF8woAxe0xOIxX
EpyOm04toFXIOBR0wyPpf/owJD6Y3oPnojASgFxSmH7yqDzkrk4U2f/p7yj0/Qsj
Nj2R2JGh3lMlHq//EAp+p1c9MQWT72/+t6lJV4HB5ipi9yMth0iu2+GKN9QGT2oc
Bufy2rxatqcJJBFffWRsZYZKwjc0R4S7KNABQ4gdZAikUIXd5be8cw2VstvAiY/b
PniRndJEYXO2aabgT3fpnfoksw0gL2SX8lmZiVQP6plkRh7Ue1arCsZH5MaPTdiM
MDmDL1FqmnZLFEZiZ7ka2yCsB+sj0j0jxNa4aOstTkiRUXqwSp6JUomdYEC9nKmo
JkEwcXw4lZBpBVMA2kTAwdVxslVCumC6lINwCvFdjbaDw0johlDGtC12OIHuF6F8
tr/bh0t68FvqwYjfiaHYfEag83reunaYgM0m2D10Hwy/9EcA23K7wRBlc1m8TYqU
184mkHQkSbaSysqUSBTN9TU6Z0XQNk2WZ6GttvcRYaVT9RC0wkNUNxtfKvOuAonx
lhE9MDJc4LC4QSWaqVCtLjl59BgBZPP2mZpZvnWflKcFMj2JWc7TVP/7dO8xepj+
S6pxDYIHlRzuvaJUnI9DwKQiY6jFllgG4uJrf5bRfp4HPr26rlnv3jR5sZF3v5BR
/llOyz5EF20T2dwT7fa8KrxcmdKYofBRnSiHvM44pkjv5Trx6VIURQNhMm0Dz706
4hElsWdl0pwNGv1IHUNpcGmijcziH4KphO42vD3WhbSeC0txJ6KP59EjB8SkvWZl
w71snoiI9hfjD8JMckIfCzQu5WGAyiM9pJOQv2hFFZDB0gJkbjNkybtgrPvvGVVj
BAmSyDMS0ZTBujj6prxKZ1VVJTpyWioKxLfx8E2gokQ9u5ss2U+WpIDBUGYrzCo4
Xo0btbWs5rBfojEqYUODtHdN6VvGSe977Cxmr7E9TVZtBEN6ScXNWRzMrVJe1kuy
CQd/2nzZVA5R8XEUmZxo5w1Cu70KZTuSmex/1mWGvX4tAwLRbgd6nuKVyPW3lPO6
6YkglTRIMD7vkCpdY55oHAkv2PijRKqy7lO7FzvDALU6DbXcuDg7uX1sWLosLJnd
SLq9sdJZdfrf3Q5tRS+IyRaBOIJQvWvtEMCH64dalk838xCm9+dw1RHVl4v7KwSk
HStjO97ljDTVEovEGUOl/lsXRXeXflb0EZXvWvTI3gG0QEosC8R11qu4Hbc9ikx1
PslfoKh36NiJ9yaEWgFEFWpWuX63NSb4anCrLltymSs/JZkKaNlICyqk+IQ/LkKo
K4Lzb09rpJ4k4i04HTcfTEeND4Z1bKf9wSG5rVTPhVsHEGHnNR4fOGMBa+gIUM1P
/m33bAN6T6sfDGr3JWPQ72ByWtQEoosTnCHPv32ckcy6abpfgIjvJvdn+YPq9DPr
yTvk9T4F7yAIH6SuqDptAG/KCBPNE5Et1cvOyn+DrEuen+9nRWQNGk+kC3fZ46Eq
S+Ir6wsNsxTk1F092xXSikvRiuuBI+pq+RFWOuUHcCwzHIfekxJg/9ys3Cte9WlY
fpBkrfkXhlai4epiaV6am4ScxrhMv0MwClKmjUaobidxEdx+Acxx/JZTQgFb8/ku
H65KlkusYbldob8qF1zBiCQtkqwOs2l4nzCkHCq0JyzgForMC5NwRgQbFUj6rrrd
1uiqTCcKVNHWP9X9mx/w0Yah+N3bwjs7RA3/+MXeQ6OOHWnuTPbTPhucJIB9KqoK
n0YdhRiPt7E6CH0aOe0Z6BZ4bcWJhX2U4lXBPjtAojxwk7/+q3nYr0mPl3t2rMTj
tbBydTnFK8in0SHaQEr2E2XSio7OoqtSVF+hqJYBP6UN0HUxg/MOYPrAeeZaHfbJ
IYITk5AB5S+P3DL5JmOOL5Ue/jAcH/ci/N2myITBx80w99QxAEG2vLvlQ7mIlcFM
P/Vh/QowezkqztWOey28gCea/MECGyWc+HCYdFzd+YUyfQmKV23qou2zZRO7c0GI
lsMpOW3go62tTsb1+OBmQlNrWPYGbZLAVC/9ggdhFPjdpbVx/6yUKZh8Fr/gWDkE
zpoB7+0dUTdpKWDJbj/p5B/x5EvIo+DkPqpLANdpS1jg0a/ZpBgbRnYReAB/LTWi
7jBLgPt0k6qkciWkzklh0qzBFW5/Ao276W3C4YE7WLXPMHEjLJO9UKinX6blqNis
22MVUQ784vZKUEer+aL7pORtMWIFLCw/jgjw+F5W7VY/8YAairLEcIhV9deXkoMD
yfTQY4yafTRf4JrcoJNZCglzXXL+XgorD+ochMqQTiEJ8uuStavu3S9K7/voDAz5
xn4tel6ktUnKx9tzuknKRcwfTPZxD0DeuPgWNsqA7BAXSkgfmFMY+heAw8Bk0gke
Tx4/1a5baiq1xIO760cIYEqKg/jObhAxhnrxe8erKvrcRO0PN/XH6T/kmykA2fhO
tY/pJhZbO3LotTKi7IMCNG7Zispfi8QEurL0fkRD9jiBR7m+rBynCS1dMpoH2iot
XlZmAjqP9LDSo6CwYNP0utMgHJBVb8eTIxu7I77MRbBxAuKF8hLM55lEzLGAJRw4
kNUqZ77SaKCE4g+DgUd1xRov1EM6Zt+Bm5w8IhVyQtcnR7ypmoxyVjc57x7D16X+
8bdK3+YOy8eNn46+gUWVBHydg7FjnDAMZ5cp6D8et747jOJTM2EU5iPj0ZJt6FLT
qnpD4yMdGu2zT6KA6eEQ3+5ikUgebTPWDPcLZEf9oKf9PFExuoDmYDXYjBkr+ww9
R21b1MvNppClF9ma4BVmrUxrpldr3+FOt+XV1fWrxdYm15FcN1yYLMhVxbpid+Am
hQ2/94CLG4ZR1sVEsquPoYs4m9neBQAMWzbZEmvOpOoakEl1TZIM/H9qwyfnWhaa
8S0BizMrKTlFWi5/ziww6P+5XLK6gnUFMlrB4ovWXiOus+jsJ95nIwlXstmmRoz0
CoeXMyFpNIBljgCfHHSg25JtZZYn7/ov/NFE9aWHXKzul8MnHk5UBgolSzZCjhZ7
bBe4oyk6uf8KH6q3kBFvhbK4G5ojXJnhDBIdF8pGVtkiAz5Ffy4K9r3umSqJ1e9C
vEsj31CuO+wdpyCQmG5ns9n3Ft9qpbNE9Mk15hzB+i3x1TNUDu5tyuR1Z3KoM0tz
XAXdLuxQp745QHxt0ey5SsxvGkkn+mzLQ0fJgbtRabB8+0rJpBGcBUKvbUXYQB4R
4agqAMdApzImSBdUfN7dDNWD84v0cYU36Tl/6BiI1pL2kCei6j3YPr1jwU9DdxMF
Pe5bbuXccY+o9uIxfaxANVEhGVrnbg0BwdhjeYrX9SnUTJ8HoFsposTUeQREDtCF
k5T4E/ElKJkH00MHTIm10zkW7WEz5HXpBAL5H4eNpPRXieDkdCeIAiRK1XTUQ3jh
cwaqFO2+y+Xd7czOwGpFGcVjU56Ecbnjw5w407OjYQLAMK+DA+ckgyXP8KJmj3k9
MbMzBqn/SytZ4vuAoBH3/PTtz7gZeE6Uy4WI3IQjylw8kguKTZF6r3Dx6NVGDLNN
qxCXBQqj/VSeNd/74ir1c+dSO03PyjnbzqvRcq6m5IqtqIZ9yAmML+paBqYUu458
mq1NparS6nj5f3F1VmV8gLC2tbdBv+8WQRqs4c1pPl/ie9Qir8F+8tnZZdKsm84w
g7sSUryyYYNyMRwzBjsKzkeSLI5xRMHQ1xezaKZvzrpWrH/XHAMujsuMLrxBo4yw
tjpM+yKJyMW2GWXQ0iR8qVCvqU+Y5L9rpPbNlgO/sadwwNSKuupykElNw+0BajyL
D4/GafdUWy/Q4FQLZHJiOajoZaD1IIa+PmarzxzReZo0coT3r2m63zRt2YCHsOQT
MgU7JfO8WvPZ4FlxKXB+MhKb+EBXFke5o+UvqaVPbpfUFvbauD2r5Jqly3YHxMFw
tOJ4DehAaQLlNavHiM86pw9jLCgeS1em+G29/DpvAMCIPhlhrapbRqjSBGrp2r5q
PDmwSRelXTRhbhoz9Qb2n7Jep4QD2Aclp9rGlZ1BPNZQtUWSp6cNY248TTL5kXSC
BFr8UM7mXh7yCO9TFez42RWFOdMGS3+eBIEy0Gwvt2ROufum8wIlP5PH/KP62i3V
DALAkJnHReUzfeHJe1kzeavio7iquHoe0qdRC2BKee4Y65ELDgNFd1D004dmEetj
NlQLXp2duutRVO3nQrO7dGC+u0SJqyac711tWplQKKxezWSffCAYyOANyQIugjSv
VgZW8zOckEIb4RfbJnrWUhpZDJqSF3J6DW8Y7C177UUqXuywxEInxv3LCNQZIaaT
lQhjNLDrQkItawzHCv82BDALWdSNfWPZhsPDuoQv6Y4d1ksb6vtG4dkKkqeOdWNv
s+ZqW/odIfCEZFJCnxvzTgpW6tTNBMAG6WKLhkmfjO5GwRrT+TL+ScMT7NmXgzAh
6zqeomkk+AWxEqrqWZJEgVt3Ne4LggwvNGOYuCv0Kv1ghU90i7Zsvt+BUa+ZkLA1
XFlqpO4f44OpF2Rozc7vsDuxE1g6BuGrPsHC25sTkGO6b/1w4srdffHQoV3xn2z0
HT/Ych5SOG9+E12D+NCncBY6Z+AVZXY8HRIHyOeFVcIDwZobRF1Ou2qEkNyU2O6+
w64KqBo5Srlq0Exiwvr0nZEv5ggaU9t4TlkMuPUaVXBjX/Wa7CB7ZYHJfwuibN+X
7p8Vog99+MkJcmcQSiijP4PGNLarN08I9Ye0e/xeR1otrSZh6946BwDfNdceGaIx
dDR8XXUw6ICB4QQF0u2W1GmPaNOtWXuGmt9A+J6/o7mLY9hNNNUdXntbEKheYrm/
+cJvNiF3s2k2hBGZeoJatsO8+NX0etQyh2vch3GtJdFvTF0A+XtABMXG34VZQYU+
/IwsgJvE+wjkhQ3i0MKALP+q1hwTDMANglDFqbWa8dr3er1AtZJcqTSDuBKi3pLM
F7SwB0fMNgZVA4kL+12h/D+BpUfV/xl+/rUA6ZVFYqgyI2ZxrV+bJmLQHK41oaM1
rtpothE//jrgU7q0OIyl1neMSbTQjlRsqDJ3AiXREdQcl9vgd5tTgeYQn20GCc2b
MP4rNP573ZT14lCPzBHwuCiUR9zTG2pnqAal5ZUZKAbT5KFQxsDumfXJU/AzQsDD
MP3XcEi8TlM+EOdRrPIBtmDGRUCgygGCvscmvJVRoue3Lq+a+Hhf9k2iToJO7hqQ
CiT1f7Smjqes2P69b96a0FMgGdeXLhSEJdnHu4UddOkqBb3cVjC7CThdq9l32yqx
ylx7CApyB1hGMMDML4xoV0iGW5P2T/fCVtROEDXxGfBh/WuEtSkFgZDHbS+hMHux
AU9sKb6hB6FnISumv9i4omakUv8P7OsUR6sByLoQNdEzzOeH1KTKcbWTJaO8YX6R
/q5oDKReBWDKTHRBF0vrd/bnKcSi9IbNQCFK4uxz/YONfRa6DNWt9BckFKFg/nN1
9h8GmkKal3rCjgdTpBW5deyyfxir0eymRnH6yDOuGZpsxaEQIaE1vzpaGeE5816h
QRiNdsGzVCa49JgaIDv//87TEdUYY7pSAO48AFLpckFDeTXt16LEz8oo3UAoXWEu
GNYfDoG7C1LFKaRGNfktkfVno6ZB9Zej7jfmIRzVgpNX60GxBH119ItFxOd0j43j
6YtCjPpyBirbp62WRIt84jKabPe84wQj4q+e7DOpXLWjFBTDtUKJ/a8MW3gcdGaT
Wol+4qm5Rbul+AI0tHDcYzZaZ9gPbVzXTP2LDghOqHTIlnaRb4PwYKk1vHDpZjv1
NTWHuBQmjt1iQbDeU+nwDiWcBLZ788wnTylU+n3x3AdTQmzSt87awf9jXqsgA4aR
4knI7tlafVT4caxMKG5/cPbrl0o2+Vl4smRoseceCBD1gux9X8gFLJgcxYhnJEpY
cVios70A6Uv/jGlz0H9hApeH318EFzssRs5ZyOmOht3ACjXxWECmH6d4QjoUPpIt
hbonXfSF1aty6C59ZFPb1vIfTmh9SH46nOzESkWHBxuV0rg1cYaLs1VjNGm7FCtj
xaN5wnql5jEl+AIYZWbaAhPgTVi7PhoYeGfrSxBvdbPeXrFM1U72Xs8gP85VcvAn
J7kwSguYOwnXdMC8kkTp2FMSlvo5T9OEu0eIefGN2lNa1+3YY5TTuHcGuqJN2tby
QPu3f24NQvD7svlLTu1Tcc5sP4k4WxoQEHuHAESjI9N68jccWtHjmuun3zJlmpwX
vPXp1bqjfEkPTRPvce/m3qyXww9QkTJ0UrKPPGQInqorSW9B6bmVRHT3/EPfTVJ8
btTIfwJHjHBEvnQ9u03OTgey4Slox+KBaTw51+jTrDugXI2dVYVRKR21OfAtlhY3
J/ASYaNllXLyuUBb+6zvFbcGWEQHKNeTQBBAujE/rl2BMgHcCshXCqFvD3fM4wtY
eqApZcGSZbczbTaChGsYvK3+HT5Xl5Zv/UyQbhMnwlY5eq4ZkCJvtTP6leXnEKiM
fo9NlRF/+byOwonOk0sMd5VKNUnDfvRt6ZXI3/93qivaocgeJ4gYziJqkX3disyz
Ug4WHLmW11nWtuWki0ycBr/o9Lw0arQh/BUVs+5u13hja0lWoOH78YKF7rzLGufw
VfVJmfqwaGC8fagEXo/aS9f4UT71Dpmj6fmoZkojAIpNG1flhj6gL3y4MbLrzwhF
bzsbHElxxgf33ICirJb2GTOxKIOwEU9QFqt7SlNqerP1AsM6qtug1qXsI+7OxQKs
B8NmWgyMwScq++PoloRi6LWeQKOkdbWeLqDt7RSsQIGtUdaYf8uOWAAhT7i/rMSG
Wo7d5Hp3WpjpRtDZswlxP4YyLpTlX4Q1Jb6tOjicSrnIPFfqGxy9tpU07g8cy39k
DIIIE2KRn9PqS0cpz84xoU8oW8AJIt603xJeTQRdC2TM5rzAGR06KJMLkCSJ5BuM
XMc+tGQ5OqdDy7KYShOxpOTjyjsAgqRnt3kTi5pvuF7FJkiZp0HWtMhmU04yUA40
AglNe0D+tGetTyuZwJZXIbFUy7yaB8b8tKYy8QqhU9dfGx4TUtdsZdmCMiylhRQe
jZFUQvQwmG4X00a/sUFuOa1saSFf6Ox8hFufcbDkmaAzQ7E5ZAczUyLc9K0Z+doE
3IaZPv87R9V861Jm2nKCjDT/LSO+KCyiUmWy32KcCd7Hvedes+6HacxQ2+H86lrJ
8Ib1hz38b5sZMmp4VUtVNln/+VtfP33Z104vHb+bIcr+5r366AQHuFDAhD5l/x0/
OiyxK8tQXU1/FD/hHidYDpCnjaHraE1X8xEdNoWa8PY/yCl0QvTXoCfg6DEV9AOs
tQMywCcEcsw/LxwjM6ET5NxncDpnI6q9RoEDMmF5S3lT8zpno8Ag73dEg4aUubqU
dxiMVCeLD4lZPvl01vO+Oy6kFrGuXN1PCKxYaDBxrJtB7CPUs5EQyP4I1ijjypbU
giLnAoFSm6oYYKUZ/PImcFGcS4xiGz6uAHyRz4w4lg6xOdVgt8LaX65YSLIzOe3C
gOpd903Lvw78bbD1STrOK7uR3mTD/CRUb2ASaN/5cmUw3TgDo9CbsdXoZhylDlcM
xYsK5y0ziu/GQczJ0j1tg04HU0J2QBxWOXyDDx23jd5WYtZXhBKM7NgaqV1ls1jg
/KQKSlS80Gmm2GBz1LFua0oY8+CwTG4nJBa5Ag6nJNiNDr/FIpZtgyUZGu9jn2jB
vzMS2D6Jin+Obiij2huKGw++cVSeyuoc/Oi+guw4GRetu1JLwOmfFwbH7nXlhTig
CNUU16758u7MkHc/mNAkTvtT1UmhV7g9fjNey8Sb36rCc3HZlUcGHatzh03Kxtur
b3n1Sfxo+EN3UQ6lb412OQQ0gSEihrBhhBiujSj0nPhkxjZCZQhico5gjGhmu47h
kaDZevUaJVVqkSlGnfNIWRMk2DqZOSvaflneHoI2Uklh9maI7SIdr3uWNn+pGWYV
rHKypMqXxx4xDBnDkXNhiSYY0mT4iVQ4QfIFD2B/34a4ly3LKiyrirsH4V7Wj/a5
XZcBHvmtANTFSnQWhDoYSg7FRiWPau2MHwltZn6+n48PRjY/G+rHqowk7qUS0oMK
PmCPCd//GI0HwovMLx3/Y+I27YaOS5oQ9JaWxWhTBvNzYn7U+He04NjUXnIEwcfS
xD+C87GGIpnqUiKu5ba3zDZP7BZIzuU0neLMh8PXduNoJfucJX8+KF6wyKIuoJdq
/5G/dwOPMKKk59p/FXYHA/2ivYl53LXXS9RsS8axFQGVV8DGjYDsqGHfGUxAkHP8
Ktg8OVh0WTwGr7w5Th/ZoqjxiEEmpg74bDshI5uN870nDtNURbaoTotBgVy+tRVu
+HXjUoL4Z+9TvBqDHBXsx217/dJ8gT4Y+2+6o+4Uut+8AoU+TZxquSBx7T3oLTq6
uX4h8mXLIRc9k+q41GEc0vRE4E2DgkyBeRZtt4lnHyOUnUS4Wivbw7Rl3npK3b28
oLJIU/tc70CZou9fmvO4apmGBR+TWiQMiczt1ZL1UmGvm1YBp0YNAGmE3Z9rd3qw
XKi12tj2TlU5rTr/zkpsxtElpGYUMgKE0qUZ9kJ0134B3Ud3WVos9Qrg3k78lWzN
F8iXEfzx+Kr8S24j0JDuXRJ3am1NXPW5mGbrvLtAcpALFpJdbnha3UAocl2TUfG5
NA6sLzBJxLrM0/FX2XjioO66IDzt3wlT5Cnt7hmrJ2XDKuFSIEmaBMu0a32/Y3cU
wtO8C5dWo3k3phWAixUKsdmVmGXaJ+g8P0lhclt/y1rHN9rB7Pj9iwLbaLz7prkG
PqtLUKaniLMvldNp1ltGs/B6Dv5yAAck2IQBVcGTLpr4xd4IMFltTygibT6cqL5N
41BZQJmABSZxILDdzN+7jptPdinx7uE9BzmgtspIlw4eDM/PyLqik+ycHOmaDFKc
WbHGd7+ZdBmDCUkGvRVlanLZ9XgNXuEqnzrQiRB9ky5zkhIJ097q17tBzcZ+8q99
NmUotcRvcjn0L/9NCDpXQ1EcGIqBd7sFSyz6A/4dNlQ47vGT1hu9+9paLRj/Osqr
lREUCW7ECRPq4Yniz0yQfalJQVDDybK9fScPdLQreL6JyNp7EJd5dMyh3CVp9PTe
WeKOvwGnMEpFLYxZLfOstQHbMzUNwfKJITVacJwxldIduolTBZmGnhDtwl1tbMlM
sWOGkHQZS7NWAUjx+Aakqe+zpq5/8M6IEaan151z1ptuAfFfC0o+xOyzpphv1535
v2f2BqBQ8OM+TxCHTp5YqgEpHFwopvEqOAAykfBODE/JtyqNlUj6u+fOyLqE3L0H
eTfX420h+xP1nJ7U4mjk/SLjq3F1lIJWqSuha2fV7oavYGmAf3z/HnB/yzcjJQQb
QlzOln/0gpQKFPXiONvHOSK5aLCDy5tHRfNWtV+v/VrHXcG458MjWVugFabTQxo8
wUou8Wv2GnqZdPguyPM8dPHpTlH7YszvZng7XzF1UDhH83jxoPZd3DuQqSsxsaLP
dBDAhQ4zjWT/dociMUnyfj2XJETnXUPIRwWb+gk41UfwMmpZyBgTNivm6wFln8+b
31Y/NrqnBvHhNLVknnyGbDJ7yDTsWEvKC4ly61j8bEy4ChkJ6/7rQ2v0fNcJOCkq
A5z5Me9SHEbms1aFt0HNvOgvXq3xL8wYQAKGcORmalMLbvMmL9zua5dROpPAtE+t
c+GcEnPW9JUeJNLJwXbBlvljJu8zzHzRedycekM/HeDzGa1cEMePCUg+2+ICfvvv
T5EbRNpQCM5o3NR2CPh3+dh4pkfoZpvmb6WSsquilkj106s5W602gOUIcql3o6nZ
PXyuG/nlpnOoK/rvKg2pp/C0cXJgEmCsseuEkz/VNBTHimMOhGMItZcOT/jfnHQb
DCsGGNvHivg4ycK3Ud9ACjDtKbvf4dbUhcZh67GB1ko5dlAUbwIeO8cjt3Iy6IVp
88t+fk2xraf/TWGAZILvAVuA4TOl1KsJ6W4eFGpBIKc5jon42m0+f1CwzT8hvUMf
jxP0ISdcNJvfp0Vf8erYC48bcOysNv3VnhLm2CvgPz/+/Fb1OZbMJMiNT/6i+mbJ
Ysa59cewZUgNny4VT8TgzrrfR+QMKwPPKa9aR6TdCO3nMcw5W3+7l4fm6Z7bDWPv
ZsuxJpSH7rWwD8a6kD/nv+jy80xYv5Yrj45jGlph7rnIdwrcM0enVffhG/bfbvtJ
e0iBgcxOchuH00LinsatsYOcY07geJrtjKIRDLirXVzJJQbTXbh0LZP36d5mQ+qC
boiVvdmHS4WJ6TA+mfCWoL2cI1Lps5iOkluUGhNYkOqNcIfSSwj1bgx832sybE/n
neNP4RcbZJbgISbibg3jMuZwqd6aSbYRl/EFYHV293cgGO9y7TwtOW8SFpewcj1E
+6DyaSwWdlR9w28GBBwOWNsxQmBhQmAGQXj5T7uDLguvPxJ3CS11Oo20hNm0Dsim
RUrPHvDzgKSz4o9GiuqIpRnOzr7LnpIMM6Yp6keCFUDhkNHHX2/5xoawgUYeYUka
9+C5nADREyr8R7LJkDwpveUua/10jvEDnbal0cFydu2aKQ4v7BOLSOzNr4W4gmBw
0C0goXc1PO4uP9Pveg7qOZwzIgRsWC1yj+VoFNdxILO0XxcYWgzNXFNIDqXrOAtf
9QraHHmQdyuc0eHBtWcSbrSHDKRY4cXPn9cGJ0U6G+g0bGjk5FL0i/hx3vd2S/mp
c6GJ4zRkjivESPIpTCOUQ+KQAItC0i2TQN6HMXojwc5PvfqnDsn8nfxxMje7XKGT
zmdVxoiB+V66QsIyCznNrW4PtwGwRXrcEPuQeSOv+2VTEd2w7fCweETrPhAfhzq9
zinMOCMNY8s4Cvu2T+J8pM1Y4RWcRzA83TlFKYi+lPgd9yDaWf5CSIHMq9167GJX
jonYq/X6z+mSY4VUQ2yFddm0c5cmP8h0N3pWNcv3rFdztmukKBjE/kuoRSVyLucS
uYXnmRFn+ylvVVjiacwHW26cnMIc4YbOlmmafaByZKU1IGbcqqb5zi/pzVMRamu2
ChfHtOac+mPJV4UbixKHGOfBhfUuEnSD1dVmZ8+s2aD1aISWMwt6gId9SuGNLk1i
xAE360fPE0yJpykFRiZ3FqKEuwSW1N2rJQRetFrk1Sy3AxkVb4p/sFIZvlfgdiXE
RV2ml95J9PERXwOHVe6FUMXng2/hDKerMOliCzeKn74Vr+RaSWJmywHZp3fP25VK
fEmLcxyjqoTk7ULnGGsJlLsuYAKyantyEa626YoT58sz3y0vFhiJZG7rJ8bbUZbA
DGSy1UT6lvxsOB3/LHddKADqqtuI7cAr7vhVPkWTaKnSpNr4I5sX6ugG8dOHV2GM
gM8UKQtVAIqOCOnk24zUavhGue4zzMrPtEY25bK/Ysb1n6HgHddisFlSd4oCYMoX
ZEs86JJfYp5e18hv9mo3HTNyXZZ7/Z3pkzrHK6uaLphTqhfOuI+PN4jbTrOalL9w
1irnCnZ1oxhreaF8xJVqzMSiqKMmhUSWZsmDax1dl4mgzsUk0GNbMK3Mlls9ojew
tgaxmbFcASlvA69FyxiXOH9A+4PgQwMY9DjGDZKJUgT056ILf0oZrhoTaEdFeSxo
RRRbPiaBwbIkN23YJ8c9X6P4wOYzhPuFgDM4F7oSXx/M+45St44WIS8IEFe9JOPG
ii60QnPf1+TD0JR4numZKc+BnlW4mG0himhyvX1UxisE0tQkweuTeLxGzLpmBkhM
4buR6CrPexs8KSBhnwgs+IS+gDj0zAYWkuZcP9XyW0VfPlcZAvMgAK6RmnAxnUPY
2Am+L+MJ4uwrwbeYhc8e622/U8gYY21hVZSIMYDsLsIlY7/fpelu7aHmeGQNCfcR
I8qhhcwo7lbt71dkojWvmhXLng3O245IJnrN6xIg2UFIhT4RiW0Kmj6lyiRo9Fi6
4u4xbOT/qS7FFo+ep2bBWIqbeGuY/gj5BaEUwUxAQ5SoOWi0/Nm4Cg+XYAd1EADw
1w6Fypw3kmossRiose+ZqtHQAqBHmhlXGQld8QBmEkp8cfjqd3kzLQjy9qAqNNuX
KW6QOxwrSkaQNv1kwAoY5RkwLU26bBXJ8ICbvcMkQPjEw14K8zZalMjFGEBnObxm
JMNxV9+S8bJnTUhFd6C+YrVmCc1PbxGYsAucRS9U3lcd7//2Qc34NZvDzb22c+7t
dp7avCetvfYJvCaJl4mRvBXl4VrGhl/WjezVGFhemOFdyYroeNzHghDrA/EzzU4b
g/Mx5dRn0Z2o4/X4+ZeBm7d2nbCjd7BZRAWBvN4YvAbRrQaQrURpW1GI3rXI88Z5
kgSxEbvI37QA45dXDZ8xPhGRKdigvB/+GFabeC3ToZiK8FazgEDa1U7YoIQxMDBA
RFWShExHpnUnbvobth0ztUBM2XrndWEdDy1w9Oh8DmsJehuYTQsuPYOn8Lve4wg2
KoEa4guB+6MtJnuFowGNW7l/zi5iXJV0z6hZnqTq4Zpmj9hMZggapQNLmDbWvVhr
NQ2/4On4Ic9rFda7AiZu2vtAcfV9M1eNB+orl4BRi4dDBHGZiAwLj8Hc7Ii+kiyT
AGdRrPDOXv59kbQYKOSA5DQJc6TNAGJ33hH9qm+9Dz2i4b89hLfXmCpYCogUnYEr
aY4RllrbOVLDeRrblE0RcbHUvHMSTtc91y0ljoJXS1ffloR/X7fkJayW4F/2nh2q
g69im+VNVj1VusKChHH4UTyxU794tS0/sphklER2DHAeJPBqRFRq4TLcIFN9xdZC
F/8oBy3j7FhsVzOGHa+FCaqlj8Y8cp81fjlAZvUnAC7SmJ9hsA/EMvlj6aH3vpMI
0lrY2gm++vt63GERuhxYjXxM6KuxyNWuc/BFhsYN9IuytMDC5p2YWWS5WNmyCJl8
5b0j6fQ7ugSjdgeWHA9RYKUtgEIH7XnBLZH8oERZzjoYn2t6jW1lXUJErlqyEv+C
kb+AKGUZlL7Bk+MxNKDd7kqfvoW9KyCHQ2JaYonprSdCL6Vq498TGlWhdKMU3304
aNUCqW8drTH875/Hod8j/4D2B/sMPj2dmu2JhoDuxavqW1hkENyYvmPeb6cfSOS+
XfbNYcBZzi8JgWXDJAaRYuAET9ltbxKEoiaE7hqxMJjLhIuA7wp+qTmg6UpA3R9d
rZLepmxWBokk0jhTnn/4OJjkxJ827fUGZmM7/bJvJUiWwl4S6z152SDDPdbtJsUd
ZLziAQ2SsKcWwMqvYnZam8mce9T2wJQ+wY1K2crO6w3EJ0bQmgXnwAlGiZ5c7i3j
jo5QcDx7UzuFiZrEx9LZ5l5fm8KYw7tqiZhTG1SaObbN6VvAf8bPcTxNGXraX2sb
QRaLXrffAK8MVTbGy1zgH0KUe62ZD8ex77S7QrtlrHMdA3r/47JWFLmHW5pt21KL
wAO451GHGFIhuUXhE2o3upBAG42OsyxKy3yKcVH0FAKQl5pqeq0e+7jcItv631sy
uJ6ucLzZYLPeSTIVvsrAF5Kd2MVc5bXDfQ100mv5c+scfNlRmsIJym/rVIjNjzti
gz+/KHWuFN1Kqpw+0yzGEtfRUUQp1iazMvrFPxV4VOKOJW/FhWHObenoEwc9CHP5
FhosudVRELADodjnW1R5jNSyufxNA0kyyqbt9EblmujF/QmUM3DOorkXznsclXBb
PW4N3ajV5Hparg+W6UEi8E4kUQg1+d64dD2CaPIcxMumuWjmKNhINgUyPA5y3qtO
3fOXtBXmMTfqx6nQ3h2b90d/dWU7FGlC/CwjwG1U0Lbeh2YYuqRqXvD+Z7y4O92c
jNqGbqRgnfwI81nEv2X5nhiBe5fX5kDLMzS8pxHnJMdeYKL9m4LHME1OIyKtrxwk
C5g9SFumQmENX1w4a7quGAFmZy+PQKWmEioyw7ugo9KYxFhncZsP5PlauwWtWSaZ
faB5BB0Lo/v9ylcH0VO81beYKlt/pgxvqYyfNzub9GuxGbJLb3MWv/iin4h/Mts6
Kj5VCIxhF0v7w0tWMmsUSXsoHxVvoogZ218VboHUhjAwapYBsUKrR12vh29U7sLs
Zn01KMW3maLzelitO7Bhk5bSMYh6YR7ddC7HX5PTM0YQeFOzT4FcPagV8sfpGtPy
VEIo53CsvwHtTWQuM4Lt0a0+xPM99JvmYMwf7R0kQmCe+4zLv/HCTVQ+nII2KClP
eE4WBDX5+A5y9N0O7egOD+uAwBVf6r/mSFZP09HEEyPnFzZ/SaEfmDYSLdITYaSR
fcBlcJE6JUP+jMX1Eu+hLNoTH4CSB6fHmPdpSIvTBAy+z3WQrh6cXR+r2vujF6Ew
DfEpXeVJF1FBDFhbeUrD5e2+R1pcMoGCNh2KLiyU1y5jgjBYfPYlfIrf9NfUw3+x
L1dCJCeanjZDabf1pTSNfyTtu9Y8rSMJfPqCUY4XToCsoIznvbwlLjF43Y1Nyr6T
X7mhcmaTVSxfGrcbZsZoLHnPU80vowFSjcuJuCm2Cw1NSg89uogezkdMJ85+RFOP
/xSb4TZQlQzRThuI/awgQY7TZI9CQViesx82+cSWMqENeHa5UVXVWEsQV+3iiWCp
2jJZMruE7ZuLt/ychJRbGD5CWOouPe6sH7gh2y6RBERO1ivkeAlVfnoMRi+91GGE
iyhNJHHe5jCtp2PykqjK2AS8+ME8dkz0xsOU0SU1ZrqrdXJ4bwz7KVlKGqVqT8qH
nNG4lsyk9QadbDcp16Z1mIq4S0l0O4cf3viQsp0mCZxYxw4tkwoM1+f2an2DC2rs
xBjGCSWocD70VKNFa+Vd2fykUe174jZhzkM7+Q8r5bVZ1FrAI610ZVaA9Gpx7q2t
vNGGFiMP4EzA86vlL9MLhAgztJT3P2czCm0uHx1Q58dcWY7ECHr4V31THQKsUZnJ
hSv+LYIMkJ7F5H88K7vR03B2uiZ6DuGnpK/XdpNqwoz4eV+zFRRc45QTT6dezLMt
FdSCtVpiSdQQuQd6dlavnMVLcmZ2IKuuyXWMWlolv177e5vI0cHRokasuQKjbX5X
NtpecTZIqGURRce6NCI7rxvYdVp1ob5+fp9v5Iecfo0J3YDExnnE47IRWNs+2cGC
kLsEg6uxVGbvzZ2RCh4qG6Y8reRVwzys0oTmwP5Z1WDQH3NZjibO3sjCgC/sdBld
Vu4/pg5Ksu/NTl36E7dlCUNrexvhdj0Tl2ztwQsy50P4tSMQo3wr6qfIX04hA0Aa
dk7DWBy+tptEbr867cqiuvAJhU/tPVFQuWlCGk8k7xLGgBOhhSe52i92zQplk/1z
QI6PhVEX6xwdoKtqcSNvoumk9BD9+i1t5yJFbFtPH9qXE8ZM3CdgTuZdEKYu12en
GCdifGVkJ5vor+EUfMW6adfXbnaJ2BfbKcA7/abHHeoo8KzaIxMIyhkHROTPvMTa
Wj8aKF0PAU7rTGvNzT0uU5uVKrhC4C5hoE5t4+b9Vhgdemy8oY6ZBnQJjxr7PFJh
purEgqYGZxprDNLsWyVr7erpM3bKD4uegXF/Xp0JPYqTdeJKenAQGQHAHCujysrB
1zUDzAmOdGYp/f/axe7gRuxKt8M1iXNo7PLVD4QIsDeid+RSYaifCMsLFLdYpBpt
B6nHjMHhl8AXyTxUNEA7A3MnaR2Vk6Ll6oQ/CCzjr5c5Z3EX3mozXbgL9j28WqsM
hdrlhRRYXusNNrbzO7a6+UxXhoddpVj29ZIfL0HuInbHaquQdXVcIT4LQcal0SVL
FgA6phQRRTP2y3RTmjAsp80S5Qamjys5AAq26W1AjH3txJVO5+LE+09c7UcEEXKN
RSfEdL7BIGu53r20C3PH5p0bF20ofY0EaAln11A71t9yoOpXa8CanMWbGzNIxSHL
4kPiOG5k7+LWZHQudDGHKiW6UPTGPxxsCG1BdReUkFSpS7OHclNxq+SKIfvqWo2Z
HazTJvDUkhzEir709aMETuDr7tFrdBttqZX3ZXWn7Ecn5bwNWMFU05iZEbVpWh5z
T5TBqax4fhVujCj6MOy4fbLAmvabCLRjT1Dv0K2I1mFqqa8/kYGBDqazxMmVCI+J
qWRsl5Ybj+JCWgB894aP8fpc7JFeL/EbE/DziyUfMO6nKXRazUt/FQyEJFEezmNh
LgLzMjF/0NIqY75ZiB+N5E0+0JT44k8Bmq2wlTPvapBeaTjxOcSbMC+WshC3YPTx
uLDbO2yjuUmwOU4IS2KYz3t9WbNCy7qwaME4R5vv1j+yXpkTFo4SwLRCuYsBPd2x
qDbwRByqQfl2fdfA8NzFSyNTIE+hwO3yBoI+2qd81dWgIZKGqREY/i2HD2wmD5P1
vzgOD8hABw5A0KU1rqphAgqPsNzYJz2DTSXpCCrW8FCze0yAkX61tL3N84w9SV1+
ZuCbbsK1x6SfpfDGgbNAzuKVzZKFo98CKRwxklz6o5UhfKrcjz+xY0DULG+tKhjX
J7k2fKYLccFCHglemoVmamFU/fukc+eurpAxgx09+oNTj4SV6BQ5B/frJmDfrLpx
S0sNu8jKk+nyPmbU62Sobki1X6ZD6y7iGABLGMZewIvUYbzCVIh3JXgnbZDZagvD
JFnIE346T19IBN1+KwwodiwNxsnkCenhJa24Z0HPuHoJpnBCBdm7QBLd2MPKzXqr
CpIk3WcbTypo9ZoIzenxSPJkilY4P+pJFZOWrqVYeGvriGdgUeygT0sNV1KNHnfK
nIYGhTiATX5HOAkTJkdVtfKD/STo+SugiyN5jYHXDjFk5UYMFN1nebkNyORHospX
yKGXxOYsBSUQjidHDL8BBssn1gtfeQAa63ErPMKqDCEoKgNexlrVZtMjhZWqyeG/
Pr9iZCwgXbxKstARYNB6LjLmZ5FUVo7svzZ8HOREeSPlzz4fKVmOAkgsFmlgXObI
L5CvyiqRj0krKrfadoEmMRHbrZo8Ii11T5b0PNj4oCLvNxQBGY2w3RRhZvaCMF+9
Cj6pc7gDBPCTcKKxlnPd+j6ftkkLFS7Wpy00+e/QrE1nXX6JIJpRpZFl82ObFbwS
MW3d/5dxFznXn/9ke/yHA1S+zQgmsixaE/iaiKLh5xmXuKL91BMBdXRi9LY/kQl/
sKr1fZ7CFAyRcMxz5bsW8GYMdKam5RIP/yGMalF+RBMYxb6p7Q+L/pYP+rIQpQ5o
Z4Re7tiWX1ZBZMSSl5wS/NoxjJjmfXEvWuFmpxrxsjZR27JhAg0BZkJeHOS4rAm4
ruC4oWI5HWj24+37gseKyL6DYW8euPfWTYuwbieyFzfg4U6HXdo647sHdgnQQ39u
rh+rPwVRvfCVk/BFlJzIVLmlNO04XCSCoQOTaKhPxM8Ka0k9OpY3nA/eEaGHDNt5
PgH6MvsYLOdeQDDBAUcMcSXtXFe2nhNOQLrAZGMf0A/3KQWTo+KlYJFghK0RlJaW
junBtOh2owFszqvnr43HqHiZZNT70TQYJpMfavyjf94AWMqJLvNfIFZVKm9iVWkT
f1048277XMgjR9BPypP+rSs5E2CJxTjvNlsk/wIHtnClsPAMYfFoxk2R/UjD71kW
KzGjahCfHyuqzXZ7Y3c1gHJOjz3HxcMA1pC9o/cGTyFCw3DFnCAnoNGQUaA5nZX6
1MnuN4nVeQ9bOfNRC1hKrO7BqUowwyDe5v78dZQjWDv29sVu9vfcRP8xShlUYLJX
dd8eciBebtGzgbk13zxcCE/3eCdnAoShx3W9CFvVbm+KEA7SkBvt9F13+0HP3Bv2
J9K3xReY3/3dOS6Rnz6uAs3ENkTjkobnwf1dV07mNFSV91MowF6ZYrJibtlFWsLT
8cKywXEGImaZjA8iB0ITNq9F7VPaHRE+PD/S0gyx1VcfMaKVUMfPz9cmUI2lRUGZ
tqwcKoXhgjzGid9rTaA7x9XTecfNi6zgNh4BAJZMduwcfTJBPo3+FbUcssHUZx8N
TrlRhg57BUyKsnVkIIKy8ANa7jo7GZzAYI3KtlUf5FIMRYxUj4+qM7MOdRsnl/Rn
KPJhT+r582XjSeh0Tje/sjttGUvNao042tMTAACDz/V7T1UQsyHDRFiR9mab5YMl
Kyy58fdSSQUHG5dS6oAYKU088TL9P94G9PP7rSr2mJ7vQFY+fHkSSCNNH65ouoEP
KQCIZxh8oD1AuCx6z91vTQYCLuQksH0dOJsP5zDPuiQIml8869ccb2HPDnQZdNn0
6iqjTMO21omuCOlvUa737MDeMQkuZ1V7FGsiu2Imc8geOFTRCgd0NYs3g0TbE/co
Y9Aw6wENW+sfaEseLAxoNMNiHuwHHElFMZu2WCrbc+KwoCSqgx+WWZjRoaNwSZA1
Md3B8rjc2PCOJATWqgiGwkOQuoyPoBkkDU48dXTVsJ2nxZ92jWX2Rmqiu7e+RtEB
QP5NE9K1mtQeiY4Lg36++n701GDain8CGbTKylqejBQn3JfYGrmq/lk4VLdbxdtA
u0Mv0yZp9gARJmVpjsWWGVHPvDfsJo5OwPidyIVhmLnglgv9gvPBzDfcuK7IpakB
N3OMvW2nVuqaQLg+Oqqo9pTk5DHpAaUbpyzdc7O/R8OOscdIqBpcUOOO7IFlSZ1t
iQAYESYNotPHNzARWYmYu/stjgSE6fEEYeNdqL08QHWo2IppT4IqtsZ8TOYZ7M+c
kG3220F5KnCKEvmcexz2k+nzeg1SHPLtl5YC5lgJPnGae680CeYAY8gtQ9lAWMpn
WpFm9ZOZ+akzhpem6fvQJt62a3YXLnBzzYCxvbSG+VsR0VbPdRXArJtup7MSug9I
ONvOMg4YojwxTK+0eUsmsyvm3UnQ3b+tYN3ypw0XRpDifQ2ntSDxZ7orDZItuqn5
qIAhLhgWGjheTB9WphfinKSjwYIgStWfXm4QSrl38z+Xa//qYapmVtw96OPXogQP
I88QyCO0WtQj/3ercgGFdxamyX3Bx/weyYxRnqh5Gh52/b2wibxarbXUgxsejJG8
Ic6LTRDWyrylqYldo/HPVtckzfh9lujibVqSfWXzI0dv4Er+lRRz1CKw/RYn9Mn/
RG3C9gYMhKgGD7e0WPyM1fUsuAOqV4IXLgexVEdjONotkh6g1/tCfxQMs2YOMkZ6
YEZOdwYidrUFtiuMF4pA90npQ/A/soMxz1lOxae0l1Q1w1k4VzOp5b0hAsP6nTso
OX7bgKs4Mh+EF6XLgbz2B0/4WduuZOZCijeNSszixauhVfZouVfGca57PYJuOYd+
QaadL9XW6UFTBFjtsUwciLFT6OgPQvaDXg6HU5ugSUQZBlUHoZqTYLU9yyzOPHN9
ncZmAJxPsAAQWHnaZWNsP49l8abyXxT45KoQb1NIfB2RMO8/+ekiF737KLidptCI
Fy2C05ZgHah5hZbkMfDCx+u6Ljl/Quji0suJNhOtn09zRLKXzloYJKuB6fOHTLLF
xC4TiRdsmc3O45kdAkXy/Rqbj8h/rE3hNKY6EaAp1NCcB01S/qGVboyd5WG47cMn
SC4OJl5iXHeIzTcGoAIi0vRaWUVfVLoxd5BEHPPUuOZz+V4oezETvRLg8vW3ieCl
UwOZ+kfKrTdZSbxR1yMT+qjQfPJH77Q60540MHrPpt/o2nKJkZRWX6cj74pggqw9
Gcgm62ZhNrEVyHRHn31FX4QziGhF4TLp7saaEfQ821Hgs/apwiwcA5jLhrLMuFnp
44ho2r1L8DihTVQuVkUfJwYWcmnmIa9YrFYyP95yplMf9PyzjRQtAAnbJNhbZKMg
np79uPxujPbl2E6a4lRLZq6WBKvSR2vupF4tABCMQ1qgm9jE0Y8lYP5lEuJlzWhP
huH6LSl3QxN3gncysC9dYQ2yBOjX49v/ALLRVKbpTplIbZDFJV3/3ON1U4aOX55l
58uTosYdxRIsYfoa0PMx28rfCORcI1fnYSodSfm2OVNL9iq0QtOjO95khnqAxOJr
fzLUBvN7VDMa26L0fnD2Dj0CiYnkcizdGJAYAKtOhj8Rdzd7kFIS9I4cK5lf3MHX
EpysoHXCfmLQ3btk2h5eVNBzFCYNlFpN6mp7y2qeTdoKYWDTs7zXUIW0uljkU2S4
WsidPGVGHknMY7HOvI5oftb+6SN0CZLJ/NUmpby39OaOAuvDlDpqV+cRCYHwmXzD
MusgJ3CxZvbrJXVjP7eUDaauKfkY0TUjHURVnS3V2nADYW85qicBt4NmDdJe/+AO
rPd8f6/o3Hcm9z2h5KOgSPHDSLIn/WuBjLWHypnjn3AlhPrRNgI844H+ah3+2TXw
88Yz+ZpWCknvWxESHJhBBU8FPnIttQw1+SX2aNNYvquR4sp9I5Ca1Skoj9fIToOS
U8YKYzPb8Cer23f9WEfxSMIGUnLAAe/YWZVVoExZ+XXHxZsStAKyWsycez/6zltX
e9KEkIybkFImgmeb5TJK7jx6xH4B86DUt2yKLKuZqipwdOjD/XFrEZuUvmFtmwcY
sdlmGEiUeglVSOGj35m36RsXf3UcmHkJkneXYo0Rr2yWauKqALABMY9Ih9OcbY/T
E1/1sWwSTQe697IWrKzqv4RFm+zyWcg9ZopnGPZCVSBkYs8DKJh28n5tGAYnw7Nh
T8mO7nepAYC0kSM7Jq07S1OHTDjZz45m8EcFIx4XgTcw2QQcOHpo2odCzBOYIWGd
yLXrd2isiOWTIP5RMRe/SL4Ssiuuj8O9zBdzlFpE4EoU4p+c8id6uVXPnr0fIdbB
kqbZrldAuQzG6q60UEBzrRmwwujwA8Vzh55N/wkmAM58NZiIwq6OTajqsuWarBBi
C1NXmbmlER+xj0MGyrQQzzkdEJmFw/hbN74nERqA9fIWNYE7RcFgfojIGTPGBYlH
14vx4L5B55YyGAk1kCNuJaLOT+NExziCvwlrBjyN+PRYfS0hQPJ0/05GIjxq+GJG
MjyGitmim2LVBizivUpnmHnfvV8r3HHlya7RYmoHo9do/1vKw9EIsThUPz+2ikhM
YP09LlikTvPmbjWM0f4etpaLIFzR9sPvXihodiIQGX19ydMNeqmZeG9fh2e7V9WI
CYButZy7WKiE4rMpQ8B/TFBUgWJ5Yq7JLZXmRoEc1zQJ2OYZBapIQ/+GkAHEpYzU
3VNcqrhmbH9mwF6REWAFlqIo66W3670KH+a6qZScqIaqHzLor29ChamjfeoLKJMn
f7fglN+P78UTEsR8plPbP30F7XAwQ/hLRq8qDRcGk7c+i71niTlOrOH6eWGrBKdO
+ehqi3HlnTDhsOZ/Hj0jaxpZKDZC5hka4xIIRKEJifm+ihAQFUAxSKRpnrCJwHJ2
d4amAnodzo097Lu7k+3gDFdgIFXMhAHSM/75tFRw3xeBgxEwuPgVxTKV6A+ha54w
pVRh71Yjtg3Dt94dEopeLcInbAEJPxXHA9fY2o9QwdhJ42odRU8S6nMt5b3LuKUS
76RlvAu68ESoKbUFVM5rn385CpZdowJU6ochAeuYrFVq6K3+19tEIjEqPPyw0vuy
JTvXRwU8franqk/7WDXEEx1u0FqbbpOFAk6vnx/7HlbPTHZeH/x+uSWZfveD/ktV
uQ2nk1g7IIz8ZZMIPN3vrSrFsX8+8ATgUcBUm5wmDiOKhhC/vQZYi93gABjabY2s
up+DsvHx1Zxfuot6NWklm7+2nRjZJFjD7by79SvlnVg9ldI4orOqGpbN4iXE4vuG
tR4x8UZiEBHwY/aHsdIC3hXY78VCCi7BRvS+6FQdbJNdA5P0b60jrTNSqYEnudfv
gSqEaBFcy15AiPcstNiOkhfVTSJl+qQvSDOsPLTXlqxez91EPh1Au8oAN/x8FDoP
+bAuOZ835KfGG+vwr7MjmAwBNVFSL+lUHAMMWAG+K0miFXOaQcLp+jBS21lgtner
qkKnP4SJjTwsKshGuwXEN9cY0eoQF0mi0F/g3EjxFBLXWx6wf3lFuxmTAfqwFbNO
OGq2YXSu2evyGtjtTA56HPtV9Hm+w0ypLE+SN2OeUx558pXpnEZQ5f01dYvWj8ly
io7MmqHo7m1qex+g9m4T2JjEdN6N0IT35aRRa2h/9g6qe7804OusTouToc+brNSF
7oEGFA/s6B1D+5+NpKJlqqGiS6HF9tEjxPvu07grnfK6GQtSy+efw/q+8hozz2IN
isEBqnncezGpPwqUkZ0Y/qD0qm3wBD/ky+1ixf+S5YOx2wZEBOWpfc1oaKeK4vXu
K5NSveQQd7tAJVXWvCR42LnSACiyQGKvQI9cLWLXfcWiimAtleaGzMjl8gREJc3Q
x71Hq7HbXGMSa++3r6it62VrpHwAnZNx9dtg4HkVFitNmYLYSj8EISdHT8tAPRwv
TjI9Ec9raUHR6ONLobtUw/qc2eqbNTANt12kRd3rJhVhVw8Kho761pW0ufgjdszq
3Ao3P6Dm+fNoKdsnAaXUie56uxo9SSySnB1GzEFhVQumLjLAviW4obgJQQOC1UW2
rCJmF4NL9d1NWCJKNgUozAeLGqa4f/2KtLD8TlLNliAuxeIIJyPtRvgaA95RX1p2
aK+8l2fStdH9N8PKVvk2vBkecHIR68jpQmHxolBqfq763lRjZ9qqELnQw2UIePwL
6M7FKGEgY7jACHKsdoFW3OyvSaIn65GaRnjy+if4aFGMZPJJViQ458lmVyz0quEP
Qi04wWi5sxX92dNi2AK3vNV2RJ9EH63d6jJ/P9HtZn0cNfiQhkOTjEGwQI22GRbU
jOXvhbQFGpuIM1NPdsMAX4Ea26fOpSuhwYObL6+mszTaRM3n18MwdeQ7MOqnpUH3
9qC611h4kEpTrBrSCxa487lwB22ODk4d9CtoJKZLZsK9DekiaTjmFUWAogV++gg1
5N3mVor7h/8e4FQ9w8sV9ym3TQ5wMpjTV8D/hasz8XzQxKTYWoGzhnHexaWsl96G
C75zOukjsYN2RZHTSPjQyLiehI4g1aP8hP3h6jED9VYq3iozpE2qtchAL5W7soSY
zMQZk26I1HLj6UYwuwB8yilp7VF407uQS43OeyJHKMuoIbEFoOTbThv4Xv9OPG/L
6IW4wqSFTgs69UimSb44t6BULyTHly7gFFYp3qusu/SwyUGjQPcE11YjsPi8ZSqL
SxT2mAMoCL2WrSgB7znWjHMhD5kgeenfLsMDT0WNbe+XmSqa1uzbIii0aiBxPtqI
ghW+RA6Zj9gMlbspOHZZG+OmG7BGO7dlJF0tXWLpddHK1vlnWTtzPgSnsnjJPo1H
o5mrLly04LJtV4JJyWa/DInykmR8nqnVsQsIUAfkxHBnsoa2sTJ666TaTfbWom/H
TE0AV7jYvapYR0mxGzhd+B/IocVHrl4DJVmtfBjny2Ss3uXm8SzwA6E35AMu4dAf
vTKTN2tX19p6BLWtAMMhga6lQ6+LsoaHxKYTR1y1sMxRPOrCM0FC2clCcxV44aTe
MyzHDIx9VbwdEKhX2tHIkDFcK9K4M2fN+z+Ppk1niew5RR173kmzIMj9RX5vX+ae
9LzTEX/1FDSpAmxFvip8cdsSEaagTCzz/NQfq2/zac8DuX1WOk1fE9HWw0Gu+Oz2
OtXwimfT1Im7RD1ASCcmaS4GFuvXyE6DzTRUbkoax+o2Vo9SlxWgjJzBFCYuDob6
wxGzk0kz2idCBtjhjl8gF5T0byqw4KGwJIKDo7sAmMhfh9fmBqlW/PZiQ4vfNwpP
3gIbHiMAIE2H767ohge26+YaW7iCH/DrxWBQXK+VfC7+pOr8gWCT2Uyq169gb0n5
574zjn0zezWWvNcSZeisbkuTEGSF0ueVQozJplUrkFoMRHm3h5ct+D3iPvn85YCP
xLfsNjILdehMe1BVyF/XID2i53vlX9tr8g1UXjYuWUV5LlvLkmHwmSQSsS4eOnyt
vhzFAWFbRqnmuoimR0bVx27mOnKqkh9AyeO7rQPoiylD9xilzkUD7ohYvxTdVMfd
w8G32ZciG6TqIoCm8su43ilcO0Wa18zSlks+NdviFsHImpHVLyihsPxdf9sAYa/0
3hUKLCmp4IO33Bcs3CnYOParzWCzA2DMnF2AUYCHAE3cBOrisGZiiyyh/UWQr2Q0
BKYIsKXV8I1pKj5HylpG/QeQOuNfMWUdkBj94iBSAJhyKvcMpb1/4hycW/Imbqi/
Y5LF6K8mrIWiy1mzMRqfUiltk9gL6ZdcYmWzfTXjiHTnsPCvRyyOFTeopNogdU0o
HJCF+eCEBvfOXQosjIRICZx8TulTvM28nI/xiBdfhnAVWsHbaXzQM7x3tpKm+Bq3
RjtsTMDshZOJW6JvjLquGicnajkZ4Yyr9/FaxyvfFP7Y4z15fdQYEXaEooPGFHOO
FySbDIdHuIq4kGDNm+QcJjUME6CpXNlqyueLpfJfj2BhcVqYIELAxmcgy6LDUgR0
UmfFT7TjmV9jXMx/MYJpt2rBadB0WkyRcAJH7DLVvXUKq09NUmvPp6+JCoEvQB5h
bt8ApFfa2koztgu56k8JmxEycT5fYmuuxSMDJ5ewJTW7r4uTvI5MWDw5aucAamIA
rPo6P7xCBUivHSFNbohByzWM2VW/P9aWPKE1bAj1TQZDV94S5lIlz42p4Zs0e9+V
lkc/rWFI1lBQuRzzbCuV5CgtXJvLcQ8gvAxM/1lQTpe+H1UpYVh4HMz6BfgWeLPn
AUzmkOmLB9IZYcYOOgbt8E6dpacxaaCmjnSBAQiu4OWyO7ozd59+D8KTj+gopvKd
PJX1kA3CL1hJOPHE6x0cQ69aDGmtXe0twdv62dwJeC2WxLwj0mY7EuxTs5vTbnpr
q8dvOvWhrOL6SonhtsZX+o1Udi3ZvYUo2Eq6GEmHghzNnEI/zxQjUJZk3vG3Nu1B
YRiZCpTHeLpT1mFD8haeLS4LG7SpICKHbXPCyKxa+8HgA2Qigu0yW85NEq/L2CCL
ShUi5uRDiUjQUHgHz2B6zQKCD1af5lyS15n4K6PMZ53gUkxa7vQtPCfnoFhyuBzm
h+FsTtFDwmJXZKwQEvBU9t7etObhWOLKY5RxTP6/Zhe/7ioEva8YjVNlwOWFvsys
Rr2upeK2tfF63DWvTiK6cKkoWDpUdxVEu2/OdGSNLFsUevmZzvqyjr53Wt9Yy2UA
jD9tAIULATJGsJiYUHsX/HCGtLE9DRUJfI+NeaD5B7JFqo5nHfUE6WkLXLJRZNGo
+e/SyuGtbeo2B9xmEBmA88r9zUkbO+L16Rc69rpGsWXMekSTrUqAxi9L4N723E7r
Z6nwClT+iIDRmbjwyVdKbKRGOaekA+eTXgwoMO26uZC/5lv0W/nu1qMWQGXrm5B6
zXibHNZpWAIMCnUaH0qre9NnnES9Si+nv6Fb8NoUsWrBcYR+sXn6X/HtdCTCi17j
dQUdK60LVb/D0cxB7T1vhlR1/qmKlCN7kaf1nnaBS6TracLvhfXVt8C1GBnJNx1I
SxxeS9vIlVGRLtw8EPq6TF2V0/mbzoPdzWIFCg/6aShgGRs91NgeAb7EuPbwamtV
FqwaA0kgYJmlsxTUvf4PhcR3jpOcTmmYyPMDkoStvzJMaM+OmNjFlJhMCQiNdLaM
8HCnQu+sWQ/vKvOgAxynQV0s6CjvobdyMQ/WOdjp5/lIKrJRTgPoCHkqTTsf6MEt
zf/t351MrIxRsuHhOGli3V9btZNGZQj7kF9DTPXBjuxwPmkAR6zWkFxUeLQ3xhdt
fC4Xp1PTgBoVCIenY7+KOhPXllSXyjnL7dI4/2rCsfvoQ518a0NDJ6UIroG69ptX
IiEmX/Nj1azmAo7QYUbwxO8XK0SdhsxB5qTalmeVdBa9L+D17Ac5KprTZiUHA6cU
bGCP39kzpUuD3AqBQMO83npdhIxkaSHMJcwAHMoJyqTlLVd3RWORwovxeuyix0+y
vhv0oiKbIwuBMXjH7gOqIUUOw8LehGOF61dOFrE6/kBsz/XYIOxll6C0MuHAdUQM
Vi2MQCSFtpUxwgzH3BVmvCB1m4Xt1BmWqDgTNXKFEQwDq7k6QZPiIIhxDXGj7HbA
m6Isxs3gYIOPFapFL2+cmksD9agXCj25azqyim5WTgD6cUdRqqaFVrAH1iPba2Bw
WLl+FGVlfcKGqFMPJpHk/3xC6K/6T79o+XgUVshUcsrg9gcKxAbyO1DBW19HngJO
rOuyFiaruv/z6AYnQsIkdkPwiTmdd5guetOUOxeeFVc5710CxWj4ytXeeOkDSXXK
yMHGxj9pJNbDCaPBoMZi4Q2SB2W3DHsYiEQZgeZwsysIEQS+eyOoPrsMfqJW7HF3
lsM7MQcRj+5KowLwpTRnaDWTylwjAU0lXoGYeodqLQ5UWcUOA09hGUhMdWtDaNaz
tPCRjDoRNrPHOmAW+WzFzwIgpVvgfPbcO0+WW2visDgoPf/q2t9otdgJkRAmdV/y
NA8IDdLfcKHdA+OEVz0LmgWDJgqCk8X23hPoG+qjXiCqg+rcF6+kYG7CcmWLgPSH
lBgTJoNoJ3NTCZ8rfrHdfho3HOqCpziRol0ygU6zWrJm0wsYrU+1fhKCNgvtMMtG
JZzfLs0UjnIrDCVPETGnVylAK1sZWJqjkDo7g5+e50GNg0IPa/FuJRXiS9qO7G9p
FHOuZ08UaUbGDGd354119okIKZ1hwwjyIqT4g7xFemiwiK5YLVd9Q44fApQ/Y/zl
QLZpFut1pojLam8RBqT+RMGeRBb4slNhwuiOnt/LGDXl3KysiO88GmPYm8qGLkU8
nDi01aWrraeBa9VFqUrG4r7r8BW5NYKYMhBLuyDJ6nnf4ax8+UnLFOc/MFEn69Ed
Z3VNQxHrlrwckLufh4L6mpw7rw2a6Hnfr9Nf7nefaqiXveksm3Bxqh2o5Gdj+lp8
stpPRdI4G+4PSsW2NxOMJvwebMoTWPqDKp25bn3bHEgpBXY7x4UqokupVv/26v22
5vGViNBuHJTZi82fpX7l0EeQQQkeCRryXbuK6WVdqFHhE5KCk+OZDye2Scte0nv6
8vh6jZGw4QMpWDGCyp/spuXVjxE86WK5QG+XOD89glmSvBp/FOovCqX8pEWkwuqb
X+E270v6Nv/YsgcHLS5LHZ3wUqDlKNt8G1/ZbQcYJP5Q5myLLw+AXEkCOFFeqLBc
Mnk1mGq+RgYDDcTfaGpJ7qc18kHY/wXNnQLCNYxS8Q/DB6jp0pQjX4HCq/9MP6/s
IqA49jri7X3WGzz70NrZDkMKoEIq6/zcjM2Xe+TNMbTPhN3bmD0Pd5K7Amh7XUru
FzC7cukRCNEFiC20eKi+bfmaFnsXCdlybLuglBLU67jz/6qiHDWV3EdjYX5YaBay
Z7t2KmaabPTly+z58DnCgNlQYfCoLU99Ki291a+Mzyi+0VdAGPTuKzYlrdnQug6k
1I4WN9M6ltBUKMdhN82OJ5qGfeMzfcv9SHZVXOa9a6ORdwxtSNksqxi3onJ3QsY/
qUjVup9tC08fq4BCB88xRAecGFxAKbhPUD+3vJ7/LLLo4lsW9h4upxaKapHnyCtE
0rr7G3umhZaKeJqXiWTYUxQHY///q6x3whuaAucmNTMIN2Fj9M/L1SekBcgSqqkg
L0NAjhFb5FbYIYYqKhKzPKYt1F7xjFIxN8i7koKNCCAowqItneoAxSxpvGLzre0Q
O9JULFWIX0JxIZfDXPz1s8GSwg8Y+ANjKZrhZ9Kvr7bVqHB+MPdumWehnWmVdkTP
H+wzEUru3oBGje6TAHqKGUCbnUuNGbtcpDcjVd4+Y9GUOD+DcEQSgPG/bRdoy7e8
VHvSAC9Ao9llc6ISTyZsbdS59XDEobZZw3AxV6WRcUzUdqhEHxYAJBXGgKzT9ON+
fOy/uldQ6XgYg1h6pdBwqmZF0dIifjyAQYkosNTIYfIre/sy+Jry5QYYzvoE7qBy
acH5Hazddd9SUpo1yQ3AKvU9Esj0YjPN5JiRkfp2FY9QuWinswCZuJU2Lr7hof1P
u5jbkXXw7VDfw+HeCqCMvRpeBRmrVJsmE3k061q4p1zOO5UEUdUN9E3D1I6/aLse
obBPt76tJl1u7yXhkFxlicvFyEaB2/GRJCIGHyD492Zou1ROMvPOfnheeF0gL13C
8cxx1qzQDasNvAm56RSA5ziYyCfDXgifE5I/oXl8vroDB807jicxNVGwQryRk498
Aio11y8ZD1wENkvLVBKLui/csI3R/AE5sIBviTlNizSrj7oQ8vCflyzk7WkHGW65
ou39puTHOq6wcUBsg6ZUWGQg0Lpl9y/8cPUGSyU9l+nqy9h9SnY2n1BId6Ipd/ZU
RfjTWdiolrSTEciHt91h3zp2I/eL4zvRqybBMIxEf2r+FYpW984iHAZZtW7qX+j2
bOxIn4cDIcaoQf5BQVwJBMccIR2q45qRUhtpeq+bkjG+hOnOEUdvh+JV9Oe6IMcC
ZYmDUnlpY3B+1SNHwz5hkn1UUyKIQIrg6E7qC+zo6NFTr+iZkcUieEm/Sr7Eb/y7
tq+/eeSt+0cKdd/HO6Rn2dfqq57KzsEJvbvylZexsaVOiXve8wlT1f55mjvIy/2g
gHsAZKN5oXm0TAnG/I+xlwe21qcMm8UQv0sM6w/XF6lVyRZE0JT2nbouha3pUfPP
IDPmF4s+jZWNaXWWCN0+V9a1XW3Hn6ZLUMGkn7Mibyuzxuy+uzAbmiaaoSPqGx+r
VcSfpFAEtxBDt5elUtfkTefWk0uokLtyCceXdUS1C/dMeR7y6XfQG1sO52zBswwT
bPFv6vnHXkUQz03sQ/e02Oi0xwZAQUFPbVfRs9DPCw7PneBmK6Ro3lgB6otNjBOZ
qqutvnsvI5wKm0ebfsxoj3vlz5AGregr6VyohTOP14gkWs2HdVINGVGOK6ig5lIG
3PatpJI/m7bCoan5fOzdlC9KMGRaPeu7W2h+cJe+iQu7fxxyonKqqyRhihmsy+0x
mCHi8geoZU9H61tiYY61GJVzO5P1y/DQt4USOrLCV5wIkapsdUuebzEU5WLuvhYd
PchTFftq+RZ40eXlcQqgOkaTOZEarl6sxRheD4AfqlCf0I6SrYO/rJ9n/JN3ZZzU
hQN1kImSWfkmDsTNKnZ7YOOrOf/fx2MP+SldrxqT+HMAOZO5SudoN95gSBsqFkLm
wlk3q43OLT0j4qAjhi6+dDjkai+EWgfd0/B8Y0U2pQk/3apchz/IoJ4vjYtIMa5r
jxPbjT87lM/Z7Ea1bD3/6gaKvnn3DVRZpk5z95vZPxZPNmzNIFgMvkXp/i0f7RJu
5SLDYQlFdWCJDNYT1haPteAvHvaRQ8tHYkyCL+LHHKME37EXKaY8Apl8Muo0Kmys
EJsYqQBVuD4+1DTe2iFukGSuK62vnb46hr9dhRqFNmgqpandw4JvZAGEqDiWSAYx
xoYe7J17Sdz+cfD+zlfMMzj+aMohiPz1xtDdP1BEeakxAlq/XwZ8aZteLAdBP4ky
pCH0XBiffi7+/kmuRp6WAyRxq6+3TrTa+8/zyvZM0zHiqIEs3ZQf/7glWSel++GN
cY31MT4Za6OdhRJ+s72uJNjjqko4L5tBqx18ykpCaq/hjkrZ4OhUXfR8ErKvlwPD
LdotcYraVqFJgqWMsN/Rqqk3WJ1UU+sfgoiH/dax6KElyUMQJCKIZCXHybtEgxhq
SP55XQKsN6xFFKypgMHWfft/zFAZiTBegBSj+Sn+zipR8dYGLE/Ch9W63J2Fj+He
mYs+X34LaYz40FlB6pXU6dZibQk97vt0t7rG3yjqZwawJFfXOdr0V6AfkskmZazd
9ygVB7FVlf6iCnqPrbYWBj6gE4zL3TXnWBdgzKMBTmIRic3plzWjnrzMWW8pl4ce
c64UY2csJb9iPInU4Qd/lrpUoBZlXfb4Q/jNo+ysdv7FY4L33Hlh+yyooTnr3U+I
IWVIWk4AwmALwJb9f16VWS47DY2b5AOu1rFFjzlqQ5F7hup0O4X6YY+3Cn05iZ2o
+4iSJhq1TFPAxqu3xs+T1oBmCwmKZBDj/1GR+BwA69NBP3KptcfW3gXLpSgwCQGi
/dU77gz1W6Zve/YonZxWkFQOo+ZBp7bStmU3jRwiW6sf/kbEgh3XOKtCBP3KfKA5
7LlPGlFKKQ3uQMjn+iC5msCD8MJ5IAJfWX8MAv4ceZLZLuSgNBygOAWDT8rKf011
2aJbNvHBUmskH8fwILADyI9emrt8eadJwNZsJcNzEm8drc0s44LcxyaBg2iPHt+1
kKfhI/3FF4lBVerl+gRkW5Oaiqq3bR3ULleC3RMWPWuy4mjxKqZUX0uogytS9Spd
gVbAoq5kz2FoLmopMJcP9dV9eSbKXfwBMp64Vsp5Jc+wMeSsb+eayGK8zED+KiFl
Uux8bPL9a+ICbr+U8T8EsfKXmBDOY09lO2QGjbrMkRS+F40CB+V3SvRKtbuH4ydg
XlOU+RhiwFkzrqsKbc0aMTEfoiKP/rqIHel3okdphN04csksxMsHvokeMupCtFhJ
cBqYVm5cG6HEZvHvzUXS+TULqoAYmz4XjbVzky6lTYKY/hZS25SB9dHmEHCvo0yC
UzW+ZaE/wP8BtOBo/wk+/aYtF/9bps9NSXPAjfiPHrDQw64cMRsvlkPxyFIQ/xMw
BXdk38rx6AVgqkZ/rbUdphjouZrS8hMEpfpABVWO8BR1isJNZriRAuhvClXBgJMv
4+GOi7QEJu6A9FFe1t5vEVx57Z94x07AbZmbOR7OoZvnMrmpUS48pY8Bv+nBK5Jd
vZGnQPKPTtsMXcl0/TbQE6/a0Iy97AdNGhAP+Zsgm3+Nwpq5BK/fJfV9xRomry0v
HUX9jE23IL/Xh/D9vzSbgYBdRXkOD03Bc0248ZNYanmu4MDdScV549JjLibxtRem
xJdpze52EoahF9nX3UsGJG5xCr0UBU9M1UXmr3KmPQBLotq4lSMjQkTjEsMZb21B
RA1s2du0yU2YqhwYtfklOmjJspbusRutVFPoJVOrBS8En9g8zUhc1jzMaeDKX0k6
cOnhA8VAueCi13CJzuRTl+hqz4yNiqMO8A08EXsQ8XwUFJBB3gy5nFkWVbsIK+sS
jLbRrp3OYjdZQ5bDENPatif0bhukQA+2/L/L9VGU1JPBcl6c2aN56WEXkDrdB44c
und5LkaaD4y8oLJGAAaUtD0/ZV8pvxLnqlwXV5wlIBKHPFRxnOQ+8o1NFMJefGKe
8EGt90dAKoK4Zw3xdnNDG1waWuChgEwOpdGIrJF1/pF7DVx8H/6C9aDPV43yRuIE
TSakf+ui7LwD0lTyaWjBgHthjTJ4Ddd8SxVS1jDx19EuvK6VNNxjWMa4L4QqAX6u
BwVccrroAWYhEwxHJ5y2VEqtL5ROKlkkDHIeI5YnyRWc1a1nupOsx54QhMydDHhr
BcySsLOfIVIt5KgQJYjqZTpwIXVh95kiGoaZxH5GfzjSWfBHlPdmNVbvEUpdHgcg
opdQGDTikOTRpQm9ihjQANt1UKfZBV25072JmQnwAaZK5RAzH3Z2mr9OsCFkymLJ
7sI5OreLBRLf1rg/XKHg38dyEtQ7/tqxOK4CGsScq6dDlGrVPOAybxqjdKGq1fzz
SKCJ3ozVJjo42G0bWr2AYuNQgn/surgX/IDEEgaGKxW9ABZgE2uIrVnoQn+Wf56F
BXQ4p413Fj1z+2Sh2XHV0iQjJiyxDytWPdH8qfdPzINI+4r4EzQgTd3h26hYLhwV
fzPKNv151b00dgb15UCo4aBMB5JfdNbrn+gFaGOBqcYtRfS5FCDBztrZm1c1YLDm
hYQH0Qt/rth/daPvXzBHlA/hLoUBMLHJZE7UeCvYoSCBhyFELepg7lLf4safFgv1
xqt9ixW4xoyAuM/23N8mYUc1G1UjPQmbHKvu/XloXUZV1caFr7D9B86+Ux/cgOvN
25U04Md6qblKOlgmSnM2stpqWOGHyd5OQ0Xs7dZwIqecL6rMk1qSq0FUmsBv/FUe
U7beezvY1CtjLw/KGv+nlSDRfkRquUAaUR9ClVjgP+zh2AX9b40eRjsK+U7KItnH
F73c+SxzvsoH0VfFzAAelKprTBG+vnGnGyjyy3ckzlJmAwbGOaqUfadIFgR8JUJ4
hrO9z7TdNLR85WcshANpn5Vi9EohX6jKS5YG4K5JgyGIJiTRaPGC/bPZ7cW4qzRJ
Hwc/8NjZE4rOsXTiclZDTp0zunHYJIX6ciWZgDe7DEehTl8TTYGabyafL/xVEu18
eZ8P6KcwhJsc2ZkC1n+TJxJ/jbadXTbxiWGDbMqHNo9B4BXpZsvwfDwJBOfG4JQ3
p74RYAJr24UELZfHIKgxIrPUmINWETjBrcVU1mBFkgF2zuVrw6EyNpyp9k3XYQQT
0M7Mlg3F+8GMV7aRlrhdtVTc7cWROjNyglZueaiwHEmijUdQ7TZJ9p3ojOxY9nx0
TsB+a0/fOwhgt0kxUuIVZm/szVp1kNDwEeXo7PUxi4HotXnPaqgqKVCOMjGP6MCH
vsnUK8SEVwDfQZwIDGZZc666+fFMYf+CNC8ixKm/kxnZnchgTr1N6u6TlqWOAv4J
Zy842H10NnyOO3qxDdKyThQcFchcerYq/S4qcP31LrBj2NI+xn3AxmAXzFcTmRFm
i/jY5o0Our8/QPa+gKkkwe5KVRAAZ89PLR7aWOdcaIzzV4LxEUaFZ2I2IZWqCPHC
emuq+iuXytJJb+KImLtv1nAtFVn/tsnT84MAlSeJpmjae2YJIpVkuPDSbvSu9NXr
Ku71o0ISDJzKNw24XXKnsABPHwIZ06cSHLWtkkGA9M6oxFkwhbcHd+kVFY7FTpNu
W54f6YAm1o2+KQpeiGHw93GiUTenQm8/jNK9BhgiE4OU6chToKBjzp79w6AgD3oF
xur9nMqnHjzJJDzggdNuW18/IblOMK1kuj0xELJBuUP58BqQMWs6P4U6/xcvM8e2
OK1Fo+Q54sfawbWuibcKx6+876Yz4pAV/yrarcj/NdVTKRChWcAQG31PHh69Xv54
qTBzJzSqpshnV+eGKA8siSInc84FVCYLVSO+uni4wroyoLs0jDmbwPAJT4nnAiTR
M1Nuwji6URt1EaEPrkWjffAHtjneS8J7eCn+00vjC9tMH02mMqXTPE2DL6Q8Amhf
pkJb7J5KiBMoNCrjIhh9JvKc8/Rgg9bQrjqGNJ4DeUjE1CGEfHTICQ3tLbF5sAvn
A8Dbih41/FGZNWmROhjn+nM664kog3WY3z1zvv3bCC1V7EL99EaETkQGw2AAmd91
5BsHKlmGDS5afu5z1sdrQNv/zIsWbsCXZ6PxLvfFh2xbWfgZuSXI75O+/8yH+QWF
4WCJKizPeCtqhovYTrem9mYQ2EMANTLGrQkiOkGGFdbG/0IXpvy3nsXVUab964VD
eML9w2mW9vKQCHcKHKN2rkio1loKAeB6L/c6+F8M3EaB7jy/5bpVHzfGxdzdYBhB
1hLYLjCyUr4w+UEt9tQpTF9maLr1BkNvw1Wb3tXpVxiVH+N1v3jX65DnHEX8XTbP
1ehaXtwpTJrM7AgyEcUxy7c8PONQqd0DwJyls46mlAzujywrFtOUUUkHfwycMETW
bn+7Me+ApwMrv/I9j7WSeEwqBfyGaIlzbecUUyU10T5o8bcNAwQyec7VpJKK46xu
QjcipfHH3sWfBPcG8RG8wwOdOaJMhlgHMxsW0A8JlxbYigufkLuhilRec5C2qpXa
vsewfGuV6k+t7QESxE79IruzaApICmI9+RiIt0tA9wOyult1iCOA/hMP7h7C2yX1
4pad6Tcc7EeLgJvcdByarsKFnpZNT2gsaOliV11y/X4bwarE8vejFMckxoSqczBW
3Qk9Hu3yZe5SX27l+6DoTbEPDR4iEMf5ipRU7YDdOQeuI1KtAjNSfrf54Mg9w6lY
kuIGoJTn29fRr5i0Y79rqp9oLvf6hIc09uoqAcji6uionqkzh+UbsdtRnZL9Uf9H
2P/iA0oxO+iidqV69wqm63dRdVpTLnXETarwvYDub+1ib/+1AJ5j3CwQyjp3Dnn4
BtkjghyNJCze53raNHeYEQ8rI41bWXHeGt7W4dtsRUYnYZxaspbU1wDqbMzWc/7w
ENAuSv5jOBekiTFZeZLUNYeZaRbcBDXfT14/TUvPeYfpyAJjtz2XKY48c35msu6/
UylwLItG6XnmtvJniTJQMnxcF22qRvNWrybIBhCh5TPf0tWnihP6B97rumswAL49
UVyplDuupSbOZ5upmxI/KJaPCNNFvF3JRP0MRAydX30OT66sAJ83D9/7Pj8f0Bb4
hwh4mDDAXBZJfHcFEXxpaauIJTWKuzkVNtbN6Q7lCySS5HrIS/yieOTNwILtNSjs
/cqilzdJxDpXgjzvo4UNZGrMB5SONRkGZlAHD0udyAdnGqyGBnbHwE5GbVhVOSDI
XK4CZii7vMfgadMatjVGXYaMJM2LaD/JKRG9P1sHge1kfOlO+1kxGCqSscKivusg
TYh01udnEnKuUH90pHmKXfWv6nsvJOVz4Ivzq+PPBP4/RXE4b/mvqlB9BX+cEC+Z
wKAotmhYqvoE6sER/Op6ZsAfD+NqHi+xZSsmrdO8L8VXB55HF4hJc/X7iUVXQdYV
S5Wr9fRZEx9f5R26qG3gi2I3uHJ3BtcjhoqZf8pZ3DXeTxfVFJLjsfDSsl0e/Jyb
S0cFM3l4gesJAgqOzm9Bh1RLPZqnF3sRKpYyLcMEdQjwlKLDPn9SvRoZK9ywacqW
u4+0fytzPvyXw5fBh7QQrIiUrxZpu1IYTazubalg31xkGEeTi16lrFF2Td7Gw7+P
4WG9OCUe8Uvvx24qk9xJ6doQd4WaowuOD4PScgFZJqorcXUmqZ4rekOFMxGl/gQk
Y/AtztOGdehrEt5Z1Zw2IRd3rQMVVsJ/sTxz0OMP/9jd04RqIu/1zrGR0z3jZuWU
RBdVDCDQ3hLrtw+juicmI2ABYcZNN7teG0yKw8nkS5o7jg109p2pQrE59pFZquX8
xeKCFueJpwmhq5Z6etRwjnWasNd3vw9Q+wncF6vsQvgExCYIAv0HHN6LmWPqoJ50
D0Cjrgq/GcLEWdVeHiPu4gpi58Aa6u1eYgCMbDEzrR9CpRPwHtLHu64m9SZN9Bup
rtDKxyONkE3E04hCYCsYXc/l+1RxP0sSS+/PYxwKL84RBquJBT+woslHBlg6GIBL
LLNMkzjrNj8EbEtyj6J3Q1jAerdJil86L56mfuio6WpYsexsiXke2WKFMpX4bDrh
7T6fi026aDZh541+2fMZzYck244ynBflBaf+F/Xm7bb6esCNmKoIZn6fG2Qzw88R
9Mnzr166DYguAFFVv8DuJJJfO2qRZSKqTZsNPx1ia4P7bwTCeG0p/fAuZrR7D9Zo
HtlfpkGpN4jERoA6UlVzfWGPAVWpAvYxQ+7Hg7OfNLrOvqfwcnaQ/dxLkkI3y68Y
wNLQAN+f0d/jUHdpWGOIRSs9L5gcuRoHlylRcEJNNhda0syjVNyajh5Ci14KJeDJ
cabhlNIL+QBvb0MjD+a5iedqILQ+2WYPUIsFKtB31p7WB0WNd3u4Pud4vmaH3P/f
HdHj7Zqf0KdIz7YaJcY0rKFoW7yJv3W8C+t7ceaFRoeU03K4uGfeGxzq1UxFwUz8
wWR2ojdpYBvVR9jH7cb6mnOklLvCQHrKcYcExe4uJdKECk0JHrDu+TZ93YA0+b0k
+F8VadcaX1AJ6nNPgaMxhYpIwKC2Hpmq+GrWuvCKrgsPp+9uBuAA4VPm4ZytGDrX
cnbImzO2rfqRJG8fSpBJ2qi3BZMDOKXD8fDspS5ZexA1w2xCmms2Hfd34nw1Qa5i
xlg6CIIIEwh/ZHnB/Dm8nEhP7v2oWqTxW2QNtyhbyDwb4QYjGlZUYsWN20NTypDm
5/4jICAMHsSevyRcCN0NoouDpmH/6cFu9itAX8mJwIThCR7LAl+UuzFeXNyvMXlF
Gl8L0eRtdjHHCJ2prnHIajfNK3IEZcB+aVagqOlo63iGeJvqNpaagAhyz0+6zr8r
4D2nN+clQbp5lJ5ZydcdBJ4ySPBv+bUmeImNsZ8z5GO7bDJiH/KfiIvbdcBkYOIT
g+odNlRy8Cpo3icxwfMTE6tzDJaPgiMT7zXzVSzXNXvNNX4bdZaqbmnXi1YeNZdY
D8Hwkmmr8dwj5OR27wsaURRr+P8Slt/UB9nFJokGyL3ITXBs7J0Gr3wVI1TOXsCM
u888bY/ZqKP7V0zmz5SCHTxNR3ayaWw5KjaKE5+DUbwruR8elQH+ZYRBINAxvozs
LaEA3ModcdwRS6xEDnbXCB1oboK4Fla+yloKJNpXDg99rs15e/Ybf5dScRvVAVD4
k2PPaauBivUU+DciUoH8vYD6q4K5TU+xnbReeoGzRj7+gn6eCdHy/k66YjiI/7iQ
+YEdY+s4iscPgq7zi4WWJX6CA3zaEA1XcliBcQuPkhKqYjX2VqYZ8WkHgjUMuVBG
unYhm0cqkHUmbrUL8ilII5qb3xdBskBHExL4adKtGp1/+tAFy9/o57fQgm3bMfHL
XoX5b56R6Y/zc3/pQlvTmW5BhSZGn5djjryP0LG//Z+6bVoMiarICfBL9yXd2KPf
DLTsnDeF3ZBOCpjsFCpet+FOLBMMLkYnPbjIeVZrvtQnR2HmorHqnmnyNUycQkC4
ZTDqJsoAZgdX0ioLdFt4FZdNIDZwBGCN9vm7Jh6hSr+GMNpLF5fDhYVLMKKHX2WJ
oB3Gt+MP3Fen4x9sMdpk19ynPJD1Fz6lD4n8hNdB3khGeYS81x+ONM0u1vCGtca3
4DxdGg1jh4/KuvnWfY+7qffBR7FXbJQrQaLEuwFbP4s2VNazIZ+tbUcU690jnrQy
sM3iPFH5xJFuEN9BCf/Gf1KQTD73H9rpor2RdCpXcwS2cj+nJoz0yisEtS4boOnC
UjcdlC+QHTH+bMW7D5iav3OgNS/8+A9mRsTbrATxmGLiAXwdN54TUqTMA0sUBdEp
42j/qE+X9pUPFRXPfKd0NPIb6qoZzwpTM243Fk6xiK7BPYZHeG1VZf6pC4azPkXB
M13m/JE0068cE3OIeXTgYHFkMaxICLiX6gBhEw2ORiOMbtXW9GgbeiNOwYX9AnP4
gt0JzDgtOrmBFIqOdbASoc5uRydsvajfoA6Km9bX/ztMvLaINHwAOhLbCvdNzReZ
jtH3ltgwd21r1JpfXCiz4Y8dN+lxw7LVoWDV7hrWkbNqkg603mASjl5o2MAWG2ve
tk4lTUKZbzjRwXxYK4fd2eAGrESdAmBlZziJCaOffK7Rp+ABNYXwwU31TRrrd0aM
BnU6GW2X8svbKsZj88CE0B4ldfr2JMxd+EAK74pITdTNSNM3HghgjiJVwVbCsIl3
ZevN83t66HlBqK6fLrfVJy9xITfPe+aArj7ybdwFJMqZSdiDKQ4YAWUlKRfzDbWj
Xj/upvgIjiPORNmcxLSbmYsDZrgUGASGxVCn9xqhvyrB/OGISUYwRjCIsV2esGwA
MtGASZJ7QoNF4q1cMkcgOtBxjiaQrvI3+qQQtV0ZFSD102aaRXs5Fc6ewts2zQBT
ZqsD9/nO0pP1ILR1eTd+SCticR++aThcrYOpPw2PAXUzDVtnOdzVIX8qlyCrgjXC
0a1ZK8sQM1EsZu4xduFQxGnWq6vfQ+7QJuARx8mL7z4qpLQwy1J5vzgySUiXqmsR
m/ai83JdQTyQgdeAPdMM0t0Dn5GkTBfGIC29e3aUsG5XEhVX51ihM5lmkleJZv7/
FFNcHwLYllNadUmsI5TMPzpO4MukxRJ+YeTlZb1PevkCBvYkrSRl47/lS3wjKQ38
NFfrtXxCtpirWi25pZsSVx6ykCSszjY0BOT5uWT3CeIVEnRLpMnc+kzbNcyOPYsl
50vW5IgUnrGURJMUzPiGLqNM2hESjeFI+tbsSu0MIV5Tm1HCRakIoS20TKG2gNzH
INSdOVKyUAV3zu9ldrMcWAHS7pU34ZoPDzx/25qtrIrXEi4ecqd3165AzyJMGB+C
p7SiwXQQdoD5onYYPhyiFruj3Sj6iOhcZ4xl1tuTHKnrn4tFBMbZ5ct3z7mDjvk1
gB16aSyibjj3uvl+zONAXUV/gRMvMOqydaJtCmsrviGtLKHxqG5rfICspoVrXZYZ
7u+5sspumSratDqqTVQfHxvtxEqWT6Q0GO32Jud4QNhwWVpggkT/XgAkVWqd/PgG
uZcErM2bqrdDVuVaRCCkEHHWi3EtO4eeg6Nx/KixAORKra+dVfBchqd1pFfjqemp
zHW5tfUQN3edmSCwR8bQRjjkbyuJTD3O+aru5xtD3C5wEDXRMcyEMYuREnrUQ1zm
INzTYm9OykKNOx1yskQydPEn5DZwob+OFk7ktVLogwSvtxwRaCeu0LnK9u7mj4ms
u/Leoe3BQJedJfUp+In51ypLrgDQ05E75DiMXZGJg54fefc1Wk1G5jSL8GCg6awl
FZHH6I7xPd0JjzcrRODNg/Ma3f2GaY8YF5nmv7wAawfLNui12GvP2KzbyxpAxeby
4GUHwHgd5VaF6wF+ojng7SfNXZsHtW+pDXbdYrZhWrb7gORypkhLugtQMNc/AQTo
SjmOJ5eKvT9xKBKaEWmpa8hqy/sZFctezCkX9axsxw4zaeCgiJhCLSk4A4Le470b
ZqfbxfxdIhjqDGL6wZku7Api7RggWHnBjz76vBZQ7ucM8/2NxntTUfiQTMGfK8To
AuqDN1+FvwWcQ4UeEvVgup0rb9yMBjzzYUyG0Ah2GnAnUA4h0AVvrOxH2M92SqcA
pvslhjKLOaFJu/buZuAMOFudEzj9HK/ekbIPCkSIdtBLA+1JV7gsXv90jn1qgmLa
Igq1ijkTbF37MbHESZAqtO609OUTVRT/i/5AOLDpChcnhJ+nVAuRSqkAp0AGsQ6j
NY9qq1a1mtGtIAVw0CCCU9r1hR0eJ8SFjCiocJB8POBJQIDv9G4B/L3KzauHHQzS
ffKtFNkYOKdubgfGndIaleEujGRf2xLy+HVPluyZ1e4vdjvzFI4YIsrySSRRksPY
ZBDPukLrtkipMz4uav6QBE2/tgc9/w/kSz+OenrVIJPNkq8qdB/pGJfof0kSz3mn
3tldEvojp+Lrb4W2gzrALfnnlmxXvgkSMCxU6/6czg4Hrl712OIPIe4xt0hpo7VX
2NNXNVwXJOnVyRKx7bCk+Sjui429VEZVm2wR2axSlKE0vKJW9srC2LFezp/m1kLZ
seuHN86oWB/gjApCckobBV1EQ139rQHSHiB3sHdvZa47zkielfE2a1OiLZAhFCqC
S539STEK8L1nKsKLqssI1ZnNys2+SZ7H2Km4cPX1m9yEm+X6RoYTfpthIIzsxCS6
DeLXCEQHWlXMgoi+wypPBrvxR0LnWiF20mVbNxXdjkEm7X0a5U1aiMzHaArsbZe9
efSCmSyS6zuB7salKodL7QChp3jtjnUb7/GshHOxHPEcWIjyoZ27hih99PGWLYpZ
TePzqP3mUyIyZMwJ0lpL0krJqpEq+PLBgmTsnoA9UTmjJvrIREe7Z8h1GB7wVQDl
YUANUcIwy9OofzKtlzduPtDZZS12j/pDr5TFUMtBUPc7p5l4Ju/wzR3oQiFT9+gS
nq8ogHYxgIu/IOo8nABqgQVjdC4JmX48mqhlnTr6E7RRJHMg0KNEC6wj99XfvzFS
W1SrD+u5uoCwN0/oW6qiuuW3NjQZVGAQkxSqT8GOJ6puPyLv564bWDquqFzG52+M
SmVXqGq5TRErjN8+uFY/wr0Y81qysGYKMyvjho+OtH/S3zBT+FfuBtSS7zz+NJHX
e15FxvWgu5eHN7hVNKo4Yx6p/XO7HUa7vhNn+lly+sAnAXq2AGWu7LaSeuNr/yz1
paPucwziYGOqvla3Zf2Hs00YfA5ojESWxW97GppupnhJzx7838KZP1uJWV7HAh58
kJnLHbEMmIHmJEVi/jQhBtWfq1+PrUhQ2R/k+mrgZDTuGaSLMwzPtG3cL+erxxx/
9BmgExDa/IQnfgOLS9eTj/nw6lVX+y7cmln7I5jGPXchBa/J//YdexopadU8/wBj
jTK7frgTzkZrbe62V1O5s1ZUA9kNd9sU85cdfE6N7sm/fZycO0d97wpiQ1pH5Dgq
ikBdTUMRcDV/joiLeTdGmhw+baXvFBnAbm1l6wy4vZHlKs8IB7RMQuZ60naxsQVQ
Lool8fPCcBw4xe89I/MWtQf7CHFjbYzpFja+/miovjeJaCvz0NrQP0LcKCml4hE7
V5hcMGOz03vUC+FXFs83auiP9eX0+z59VL3EFPy32zge36lp6z927cUbeWcAPyPo
9pirb+rDZheuMTXKI5cY+gRQeqCNILPR78mpayyBx7U9tDqhh6HjsZ1U4eDxeott
F5mQkB0jb4aqMzzYMdyfiSukoGB6DbS4/F7OusviKJgAcI20wDKpnB0NJFIT1fZ8
a/FBWuO+spWrws0k/yAMTvde2zVdFMl4zR1auQOzkgzYmPKkcaNH1NoLDt+0Kg6t
oQZ3HSYq7S1bVV0kE2XLeUwi/4W8l3Jx3NJancu14C8Fq79guo2L6A77cZtXXW9V
QWCfIcgD07km5SFFn1z14d2lRXf3PMswG8JE6wgCG35T4RKrlVzRDzi5TjR3O8ge
YCeMhZx0jh3Xv95kvcCYdi/tiqrDQKHmVEvehwH2PL0iGMVKKdQz1O4WGoQ1wky0
TgPA16O88CIDaO2EsfK4kdDJQU1lC2ViOx0cEE/56vEMyd+pTqwIhYgrf8u8zWvr
KXLhvMUB1TqOaj0FLJsf8HcaBNjadnt7myrhUDZMXG176hM0lA1Np8zzs0Jyjuz/
y8zHMUCeH1Pqogo+6cy45SXllRGLgt7j0de19YlX820wjB2x5cVwLC9fYvaU4Ul4
ByEHwugcZNXEpuGcn1qKg4npBNnI6xYuj5R8gj538gvgkcC0lm7zxMCwGd8usRRu
Bu305cH9h+BwfYszrUJBto2v3MFsNTDQSyy/vxlINnb4UHM3y42pn9e7ftsdHHwl
64OI7FPu4jmTcGsx8uFt8HDmDltitgu5RkO8q3RSa1uSEjWGJSxr5JsXPvsZO8WV
F38u1u6vn9f+tsB0+VAW0DNMpR/5Rl+Ww43+GApel4g2VewdGpdvt2pIV0Dli3IS
TzcQLmiYXKD54GR7xMNBo5QHYk/tXfGiHXY7g+fBGWmoQ2ZDHcySdIbhbU5CYJJ2
1x/HxKGap8B5jix3aR8NiAAXZiZ2X9cntrV7Rm8mPM7tfcREag9a6pzZ84lTxwI7
4J8c9xSrUrCxUK6SAra/P5la2A22YDRKjIrv5z0hsGA7HOCh7WcIkLO7wBvCtFp9
M/95azrW8+GNaTZphbfaSGk7duquwPGjwILkQEONuLOX9TvIu8ED/MvdILF+/7yv
jpBIxwX38ecI+MdFVe/lrErK/+ZpgWtn6XidLhS2ElVXg6EqCxbtGwwxwSUkAGTx
+ZqBgOqDYlRrv4pWjOMmu+LOguc8zIELNidrUSUy4HzHl/bx3WimeRpS0yNMmqfr
vBFBL5o/TzCSTG5iVUIjPzA2E0uf131yU5qUqmlaW0nH6vVvcJGd7s9ck8laMm8m
ZxB126zgwvAoSNXGO6K5waQkwb2kt7HHK8PDhqaXz0Nkv5cHTbj3hkkGPK9b5Y+g
DgqLtc27d/ARSpm6qGPzczcBBOTm0d2crcz9edSO3XUMFIKu601vV9OeOijA1EPR
6ESZxsBniRlrgjzt3v7tjlY8Rkn7hSVd7DVCxdtbIbGoM24Sqys0tvNWItxwlhMT
/tXubwEuHD461OLCVQI9CE8+hGYJOEm2BQxB+15APVvUwfOPl7vljzY0vSB8aF00
4QPZfLdI/BQ5udu0fiGrTFnGXxXuJbVJ2kzplqXCYrknMIbgSGMaxJL1/CmCGkod
DtDlpNVr6+fasVuHY20bSPnRbKQs9GQxSfnkaUBZQhL50fSkZ5Ax5aCJD8saQw8C
feuMHd+/rhKDyAnRAtKbzcG6EyQ77gHB2l5/yo3dJJEMgyF4Xmy7VBg72Oe8nPyy
b4ZI55bsUT0hR7EhpzlkfAoAXxuHvB/IVqm6JieIg5ShG/UA5nwQnZ/nzr19XU7j
hGVcbKYvzbgX50TL8jnTbM548/03e603rM1sien0tDPOX0LZZo7WCHhiHCXSv8+X
S54TnUJDxeE4nL5sjtXteJ4dbSwWgCsiVpjsb7NTobbk0tQA5kTkgpEhuctHKwhq
IfXTOmdeXl1G9xJ1cHyjBOs9VJDFv/auMkhS1F/MkE0nVgoJLJomCtow+G13nKYS
Kn/f5bA+kHJvCiHh65BNoifW3RNqfWKNXqKP6nwY+XGL8JXQ5GmPp5Ss1rOnu8Mi
KTn6PCtdTNhnRcUUICVmq8wxdkAVgC0bnRuHw9DwdPlF1UPcykQA0hpKtadxhpx2
ZloR9nN2//w1an4fRwMXDjGP0Sr5J57ZQHYQiMC6cGJfhdhRY0HRAq2Y1Kl4jfAN
zhw4+HbExzmyao9JuTBBa3S1tymocQ4FnClr3PpU00F/SIO4zZx0GzutbxPn9B69
8N3NV6/loFIyV6M59U6TzNjoltXUjJ1OBFU4dhkiH+FNbr26OINKz9qZ3O1tadWg
gMCb8Nu1aWRuhInPCF06ycve4FFdy0yebC2A6ODdvKElD0fHzhBZ+z9aAnysBN3R
vl5tRPuKhMbozYfe4rukMJtgYFJD1ftxF0WpCLIzaYYDfZlRE/gjL+H6Q9S/7OPK
gk/ACbccUPdhS7tlJkK9cFbLh3SyGAHgFXgOJDZlAKaOw0OT7i2ao2TTCfVpHWhJ
HFoUSsnAFGuxw6Ex6F+5UeBIzCQO+jFPPisxmc68T7XRpt6X3drXCtGEUpzj0osM
l/+Ul8UzLuNy/OxvpQD/ksxPJP1jhiLz8Z4lIkaPTHOmsiWOuosiFvhuhl3En8Hw
ceRd4ydWoRwS1V9v/MLmvAUTmWg6S3JwpA0skzVAkIBOxClTriBED+omKOyoYUbw
h9u8V55K7jWWfaE7UHLkk//tcHyRog0W92ugPzvCL0dw8wJP0jOji9whvVaidVFS
UaDRNI2sCKDnhnuqcnWdElIVgVpWZQ5oPJJZ+IXV4inuaNrSgM2owarmO7wMBxQh
R0M+rQSxod1Go2Fbc6YjOva1a0CA25s7lZP04YhUeoWBIBAyryV8bEM17RM8Np6U
Y/Q7eQLei2o8+WxiuV1kRfZyACtpzom5ldBjW0rdv0qvTiUpSFfhgEAnnp6JjTsn
fISlfCRMOZwPeOmukSFv33HHM9LdQwpBxZlVORAcQ0E8QCFBblCrCmXBLMYLo7te
fZ2cUfsS4VHaabXTwXFXSkOp3oh5ZIqp1LM638VGFBDia1sGZ7ECBSUi/K9DJZv9
w5+d0gIlgii2j5Lyad/U4e7fG0crDK7KSWSxjjJDdtK/rV/EOGMSI1ypYLQNDpOx
COmDDjixeKnXQ3ti1W1psBISNXlx6Kt+SlQq+OnpQULieurR6JnuvEmTd/vSFu9f
ZwORekv24Qq3FVmivA/eaYgJoox3QwAt3CFy0qSdsC6gTN8QSeemn8EcDppNx+M/
o/0kkVJ2H2wUXeVog10jbji10OcxvzUI1AaA72Rya8Z57SM9J2qORbX48p0NCYdq
2Z1Pjt5WHFmKZlhca+oFszYF6OnewiC+SdPtlvkxTVXOlTOENu4IMmXAvOWDIPtb
fWx7qOVDwhD5l+1ZopJwFlXlRMLr/5St0lhcqCdijwavJrptM0HhmA7LSzCY0diz
qz/r6v5gdz4UWJgkCzHXwd1PTT6OJvFSLxDaY09pxlVsCk1x1/juy2oH427lW28s
fIKU3XtjMT6fDMJJ1Ca2eyuib6sWr9cwDN4UFtBpPh1QsgGvSCbgPLY3vOAGFSKU
JlAfZwVmq4NfI6pqrncQXwQW935b6zU1d760QaXJzhttI9s/hsXrMDN9hZaT+BnA
cO2AksUJGUGMoEcN03mrkQvG7ZZ6pu/CSCs0do96+oDbAzrV0IgFr6gYrWSLWovZ
WpL4bSMx4hTPn61IRCk/L9OF4yCFNFQXuxUns9l48odpXYnYKroeerKu9tyWBMoo
IOa2lP7fV7HVxxXgx69k9vJpLZUhljQw3QnhFfeQu9Flwyx/C0dDOYbdxEVPJeY8
HEYWQviuFuL8zXZ03bI7FVteHYWI2hoNE2cva0zK22x1BybgOmAzCd64QUrjYgNO
H3dD2toulazjEqyVhTfLj56sdCKu4eiOU6JbUEno/3zy5AUI+QtzMC+sbdxL9IGn
cB1A3zLO/0hCN5RW5q3R5uzLI1SXrSG4qVjLsJBZjwsWfhDQC2SUs05Gw/LR+o/F
Jwca6rOnHN0adwHUzqFhSK1Jy+IBS6hlYW8kGekLltKxxz2f4WF7lzsQwKiSUYxQ
JHU5kBa8tvLGyflu1pmTnXsp3p1i5wJJN5KMkJzmqJcTWD87IV7w6cYtf++Zf7oY
mFVbwAwDHOlX/oJFy5fXxptwN1kSJKswuugcYPE98LO2IyBWpdIq0txleGAb4ruv
JoQ+/giLC8hamZpl7ZZeEyUR/AUSKQDpmvrokMV79ej1SC98RjLNNMu4vjawKf3x
8skwU7kjrruKZQGOmwNMuCLRBjmd1OnyN+Xm6HeGZLfD5ZTgm07aIHXZ9xF6MYgR
xtAyX0RVnPYbxSqDluQnkrTYF+GU6sjL/2K6AWFZ5pyO7igvTg6ryUJAnxeYwlqE
CgP/zWTimZ/5WkktEqOdWP9YT/6ZqhxirpB+36Cj4JkSPSkBTJ4pcmSxo+ACqJE0
R1u0wXPuoxKy0V4HHW6jnCsWGIytaDdC7oGNsrcCkjCMYpVw4gwmVDASeI7k0/Dh
OohKEtxN5rTboT8weqR1Szx9tR1VUy/tl2cAwwpMl3RZ5sPXBx/EGzeH9EOkXVQW
dMLzj+kN0PMt1wTpbWJY4Kdt78h4kK1Uh5lNNH8jyAkLuRp2T6FQ8cEgrIT/VbfQ
76fcLH2ew2EtJGSyJMLgm2O7uiI822VxmqaL9pWm0XOG8O13OzBxb47hCu2944Ql
dq2qi2XDM9puMYkL2YzJseSYhi/0a1sLbjO+ao5x2iVc+1VMLL9uKYYFGyhN5ObO
574vBw3nCwsSm/1RNuUitPFpfY2ba2qE2txHuRvqSgdQGAQKAaVrrF0v5EaLam7F
zd90PAXI8on+PUOuqAWc79KR18uRq23SzLM3NPJZtHozmcSY87AuGaKl2pMJtlvh
0zBbBF79n20Kj0zGUR+mR1YvRRN+sphI/hSoV1FSUrvaVB3KK0ZkX1INlGcniNK0
9crfJXY2vrqHhvq+JuplEVOAYFgyRmXOO4diduqjzNIpz7w7kx9km+u+tvFYFqGy
dLvhC65I6UlA+qT8fXOx+r/8K9E8KdihlZF6OQqHRbL0pg584jxxFAs+0XXHUpnV
TcbOWqX/q12TrAVjigqFkp8WRxbwc8uE6Y9ftjArlfOKxFiO6/fpF8MpEe8ghAHI
v1u24TWqfYKh7F7/YMFhGdfhc2K2EhX1WcQp4luarJaysuIaBhkcqYMtelzfZUPT
rzv8crwpOkNtMfB1VEmBLPw61DuqWYapQQpFh/CxxVPrIwheraYq1OHRKQaMu7Bs
hqwhal22uG8kMUAyAjuX/iLy/3uipWKqF6Dv088CJvy+g3sfAWV6GfmNl3rvjkbb
AbxGnjZuJrBcvMvpMCibHgfubTJCedVvet+ps2JglVM8QfcjvfztI2kGzHa5O2W5
jviyjP0J60fRSjJoWWaer7GcKumuVvu7XGT5A4YkrrtmEM+6GvCGaESEc6dmXs6B
M/QIeQKC9y3m7NQxip+HNTWQGHB335r8QeKbcCMCMkbGIJKzpna7IzTQf1EJ/0HV
NUyif1pmMKESUsY53gM/caBxo7tcdXtxYN73Qpkp7xQcl3e9ZNWsVSy3VY8/XmD5
/LNSBNuhYSEdrF0+e5wToXw+5aycay84rmsJUro5LyIAme1x8vic2cdxPxENOw4R
pQQjZc69D/zNfxQ6pf8TlEA5hkQxdmyqOmllYHd438ztqfst39U1pj7GEpZqctks
SWI6AopeyYXuy5sZPhe3X3y980dnZNw1pAYFPMJII2j0gZUai9Dpc6oax6ExXC8I
yOydbB0t8PuVV32P32ihYAxWD/oMAg/kO8xzLVMIbZivmuElNrHMAwm4lGpG42p+
ZFPP2oiKgLi0rNs6IPzNO0u7EkNBZsfYWUdoQ8d/AJdodxu6u9AkN7YDqfnurprD
gxM6WePfuITXCPWNMOrDwHFmU5FsrRSNRQZY2zSof+Vw5RsFCBJK26cp7oe1/tjT
t3671NOl7EdVDsSElpMSoWvHxqJzATgzx7zy1RfLRu2LYZ8O6RLJb/9lU1PjgTh2
DSyZf0Wa8+Kn+UslE6SvX24Sng+I2K18Q+I8RclAAm/X7yHkZaxME0RqBSJvcswf
A2KplolHJQJePvQw8cxP9sYmhQdh+65tBKIEFOjWSFmMTR8p4jGDpNsNAcIVwGjI
MxPdOygfvQlJ61bpsP7aCYpeoUiZq/xcM6dNolzdoBSNjer+TLEwYL6MCqvUhUFh
BzEXxHkVeGHSHsitZCDvg6cFxywOGrFSWwQsAqMi98f/bYJAYblvtH/moD69KQPL
INrsQZ7SAyJu4g8HApseNFByu2miZIHLjIme8k2JCDDQHbkxXeb2q/Ycrv8Fn2YE
SiGC6z8OdZ4aTsTDdN9ZpXDc2dfbsWohATNfonkb/r2u5wIGyFlsNMy5n/Ugjn7L
W/A8YUvRcrCebKzcTlCsoamv2gSzHFjAEqtDcP8h1nLQtdANSWZpq4qr/bmRXmKa
9Df5eT5aRxqS5MW32Q4KDA00tlP4dS1RlnCGVv8PLszeb0GXlvANX32iiGh7DX6+
+EcTW+SW/hGYWgHaxEafrlJp1o1IssJ19NOF/aHA4bzNCPT9dzDK7BMG7O+1FUZd
NnZ/THTSUhWnYJ66GJKAXg5B2Rb6fkn/hPujqahwfseR35pr3MVy8Uh+nHdYwMPi
6FzshiciTJSU+i5dF0ANaLN+ovX0K8NPOpRZ42/2Xe45vDUc3kSy+RaTbMfgJJOA
h3SrdBvxA12TViM9HpLafPNgwHcxZo1WCXKHxDMbX1cia0jXd1gOUlvwvHMwcskW
jZ1OiNgEQ7rNyl5LcQcePP5S8efh7UaAgy5rtlqHgqWkCACokQ64A6QZRr9r4T9H
nSAZItFBxzupaZnZrDl6DJWyScQt2iH1I69h/z0Aq9JkiVj2HQfuVwYlaoYcCswH
7PVHCJBO0ae6eGE+LwCexYJHW4sI3in3NuxLqPtMoNIPWNAKDe1HYkaQFqE53VRQ
/py5+s/VVc2IKeFvRIoQDQ2kDAS2BvTWsKsWGLFRI1R0SD9Btv05D/meS2YIGgeF
hdsRGWlWSnwNXBTO94WHQ+7O2AQESLyQM+pysyDXoM4Vt+wbmHIZnOzmbFa1QvzR
PfZ3oT0e8LQNQ/N7vp5CpNGSnxD4P4XhrrLEfSKcYeQdKTEhxLLTwA4nVwfGOmoV
qP9vGFzdtzIeoNnpWFJB5gLcP1MMgQVsBihZxtdPaFWogc3OEbGqld4+6j0WrkZQ
JsqtG2S2Yi3lkwavpp+CmBHlCOSY09thGh5nXRaYPeoJ/6beM0BMPqg3NQ408lNI
hp0UNybF3xMlpuh4k5GOsn18fFMAUFWQpcHeosdkuU0qZuagBaac70Ok7IiaboSc
vMxW1d+wAk9Se+NqqpagJl9lHVszbpq4j1lfiJzw6yfbcURU2iautoD0X7ctxbu0
RdMMXVbMvngEbQEhaqSoGjm2WE0XrJLUJ7IlV4HB1jyE7hXR/brnyhcHPdXJVhgL
Lgf8qF6A1Up/KdyEjImRrgTUmeItWiY8aLjhB1qTsK9Ubcv6Q7Km1g7hlDz8GLyO
cgufB4eRQB9dxaECMPNqcURokB9u9YpGUN9Ffg94rIrx+BFCdQAIMbqEJpRk5ZyY
e0auK+k0yW/uNOLP8Wmd/2ZQpMwhC5qIXiZIhlCmM5tgE8n3KbQxUmnVze/d4ztu
aE3+64utO8xinN459OBmyKdz/z9bUWBD8T+tR3A7bZkNO0h3i9kYAuBIDSu7MzTB
mFQOeAiExPyt01hAuUeqntr5wcoh1Ea8/Dtwi9XjWA/UtB48QXWvBvOXosGvPTWi
4C8hMmooBvPtmTb35/7IthT0hK7Jlw8DYlEjBI1aLEhx0NLJ081L3+x+jSqH+hhu
IBQHFFqSZ4hUhqwNjUv8kJmdYexQ6TLlB1Bo+x90KiCl7CXDu7GVkxvW76WCUDht
psdN+8/XTaulR1ZOI0IkiU8o6uR11lAA6TveYDp2ur+ztrrpLz8tu6Nr9wN56Vcy
ehmjFrHIKZMcBgZPRYZp2Y7NPhR1li2stmMboG/ZzlVtU85lN5y9Re3UhtdAC1+h
3TDnVCIGtg3ww1wX9waQCsm/7d50J5CZQ34GUdNQ3k+oZdvA67f6AaXS2hU8G6wP
3MpqMdx4OYptdKnJL5FTEtZFVFveyRbjE2LZ8KzwkAFbm3gwiOmyEUX01PvD/59n
w6Ot2W1UpN59LGkIoCv7082898y1KjbDXDoCWNjzP9zBBXXtp9lRkyRNJccpcW+Y
lOoL1A3LM1xu/t27ZSk/wWE4z4LM5rdCTLOjYUhr3jyDv9md/Iyyki0BWccATT2r
VcGcY1UdKFbgo1UGzCbn63npDTkz9HHexG8xRh0k4GuVwtgtlxSqzRH0RWVV0Tgc
WJdX6I61uWA5SOPDO/s+QhykkbfOaXwTst09MvaEX8lg7xHKWaYAZYgkKfBsGVoS
bkVdl0Xwb1Euez1FrHrPk+CjzlyyLcJzxQlnp4IOssNYp4VmnJQL/CiDltlzeQxS
vSbTBc690OqkhIAp2Q94ly6FNAv8AjFdovESEA2ABx6tyJZ6kqva/Cyx3W0n70xX
8CxCtakCNO45xiHCAmBiTLF0ouUx9sutXp+GbocD6PtixG3B+kwNL+QbeIQTLpOO
FUrc4V9soJeN/qLXzzU5TJXiclH5Q6djQDcR+lr75YAAWQVg7oqIMWd3sAp7XxPG
SWlm5De3/yYEGUfbES10TxpmlSeHvHJ4rLoltjenuRSjyxm7In7Zl48/SyVYgPKK
t5WWo7hnwpt5YwGk5ivH/4ynY+PBc6j4xzrtoaNkK1d8W3xqVLbmQRzAUuAxQm7A
nIpMGZV0nQObyj6/1WfpZ+y2td3ocJkudWewDW6MSZqmNzUnw5OxX3Xe0DI3kT8u
I2sVn/d83BLqw/I7bdEnfaSDG+EtSAZ3l5MPGbxxFGWIm9imncoolCAe+tzKtEYz
ND0y24e1OUB9dZnzhRS/079h3PucbdeBxLbAb45FEdv5w7JE4FeB9cJC6AWmJpZY
vJJNC5VUFJQWKHv+vuQk5u4NCwVcFom5AjkzI1tD+zCBavZSlhrmPr6oOFfGE2MU
rFD5z2CIc+qtRBgBEqEkDQsH2JTapOY95hdUOEExT/JrQkOKH+ZBJs/5KM46u7qV
ZNHiqS2ZNBcs7hzXxEgqYmJ6F1mx8+yDzRPi8+sxbo0AEj+LX5SURBLjrF8tFcgT
bsupulPaJy3IjLvRu9s8mrhM5AUUrutUfzOR5Jy1dKx9RTJuDD9KSraT+ZznXG1z
VDO9+hyWVSRMfHrObjbWtJSiGo2aYfcPXQPk0a9SOwGLqEr8N+0tMIRj33qoMUoo
v+nMNBYXFomQ/uopiutLf8JdDTiDFiYZItO4qVh/GYkOejDDq4O9t9WmT60ofKjQ
+7TMau8sRVPh7/4ycvmWmfMwvw5Eydc0yTnzrvDlSLzj4XqW1b2GYw2cvAGcED+T
tUjOwhU6OheKggPD/jEra8XXPDElTu9CElZG+Wx0lTX7Slq8o78Pq32bVGSXOyp8
n2U/iWLGVkTOYpkxLppFuNBPKq5c/QDyV3nC5DUY4TDm7Uft2+7BuhPOSFaff2lA
2awgaFjtrKww4wTAU4MCeaTFjEc3Pu3nbD79Bo/DGTREEXn50FRfpMmu8OaKgdLN
ax2Ybe7WWqia5nu/IHpKiAIhSGBikDxqbfAWW0NsQtyuQrG5Eh1n4axFr3WrTqJl
oSTxbYSuLXxp3l0dCJ6n/vwHSUVvu7FGBjIr+4pAJfvklU9t6CQ7/elOvfqMLy+L
YE02DWe9AswpCDQtbW74J1GNh5VHwlgvu5GwvE0jzK/xesiJSg4/uvTjzxKDAWws
AY/WGdSUGv+PaH8TqeTisggv8QddMNa8QeZPjMVsOUjMHHKeM0F7QDtXUVKdipnZ
aYa5PN+IVaAUCliJQDFXu+GaXxX2kdFnN+BdXQfsUDfL28WMFheluRjNjMGeCKU0
W5szgW35WQdmsOYBRjjiB/JEmECWj9Bpz6BfoSJ9j+I5Fl9shweHVVFxelJ5u87A
C0SoXXlWw80ieToj9z8/vGkGFRTbzaDX3GbOWhPBHm0HteUk+ByEDGRwreV02TBX
7bpvm5rQQYVqRLKSnHheuHGtDoiwkM4IZ1mzMTYu3DMSrO1lSsBdxqNt5T/YbTXI
RBfiPbgwhjaltixKBZQz94XEMmFWVpakQvqbLF52EN1bSGBJK3CVcd+OckveKr6w
vPU5mU2MKDRP8hloNNcrKH4S7be0TqWJlxQ2fr+mpeNn984HJZn4iMGecVQAxDFU
ZMM+McDGZNk7brjW9SdyzXvRSqn79sUWWcSdVyAvp3EFkUj10K3lB+nlm1FQrQZ4
hmfkdWGhlYe0Qrb1CnA1zPJPJ8fH4UdxNbUPJHC+HBzZv8Ljxi6i1HKo2qVMZ7g3
n9QLucwqhzUiQQD4RI+jPXgN21Y3SM2PttgCCYTLTz2FVJ/1CnF0373zrAxWE7Fz
5dKeG2tsNi9c2zWd6XQGL6WKeTN/K+J4+xOv7xNoRTCiibBz77DKhlCe7e6XSnRB
CefNg+gEpHbQcy9S1PfRlF1TQYLfJ3/SJ82UoCyEXSD9mNBfeUuL1N0Lwv0gKwhl
KhEvON6K+0a/MrHQXmfngsnC2BZCN11aDerC+rJjyiEzMXi9+nN3gkY/tyz586WL
NghNwBgWbc7TgfVKKIsfsoPihM6eUo09Yc9nps34UCU07AWjLssBNumJ4ZH467Pf
u0V0j3/tT9udxURnyIP/IHuVdb0nMR7lnsUnhJwDi2oAt8+ogGE+dNACz714TkyF
1gPRV7HgSgzveUnZIINYfqzp8QpLFNBhIA2ubyu4xjie7GF1zbXIS6/3JDzA9D1o
r5HHFiT+Of+RDSzEb/GKNwhVBQwLjwhg1yKgL1csOx2AofmhEjfONdlLLFG6PQBy
ya5G0tat5U8guENRZp4Rcee3ZcJc+TuMVeTbCDro+1NfDwWq3KZiO5O47kxXAyvQ
GPXkZxSS2JxrHOEfoT/GGaosVJOKGPgo7pdVWGBdAD4nFMs8/F/pr/Fb4/YIQHGn
nqaxCbcWgDz7rZxGKkkGtVELxmqqymOsLgH7VygcANnjcXCFR0GNCfN1x+FiaSND
HmGK2/n/yuxmTel/vMgBKXXgu1BVFhhvQSb0ESrncaCMoUZTltFDOofPS4+fuoQ/
F3p3Nl2SOmsvh7AM6rRFGdLhiPLhdyjJsqc+B7BD5gGAAjwb2qXgGIldsDQmtTFv
KHgQx6hOpL5csEOFx9k1DqgnB+SbIZwiXRwtMYYIGfip+xe/vnPP+fYjPxgv9zWw
Z8P2kW57opQbbZTBY42ajXOetHdsUP6KlGBtOlg6ro5geT5AL7LvaCT1TNtkcObG
o5psePj7k976rteE1omu+UuLQ/amPkrV11Uq3EVhLkvWrc4YpP4DhKDOJVLKVw3Y
6vbk48aYqX1hMaFOql/SE8wHsSH2YCf2J2kxS93d3mpHZG/6gAIW0uJQ/SFXy1G6
6yrPrwOeNxFS2T59de04CWcugJbBeQbhDGKn1RxUAeWXqHuPOVgQLqjDr3YPK1fR
jGgbF09cYQV9ndY+D4zTeErMBDm4GBV8FIcowb/KFrf65UQE++cpPr76uO9SK4Dc
Mjs9mgy18sz7m10xdVDAhhVsCJoGqY2LcHKDlkhbKYISNs4nG17GypX4TTyWXaHV
OkZ+S6OZi50Pz+8Tbe43gG7mqqlwb3HKjMVt7owY4Pt1xQRdHqWkc/8K0KD3p97n
0TxkCV/VYV9j9QVwMY3NLjhg5dFEknQUUkRYHy2WuwNd/eZsj+/l52f3DbjaWQ0B
HzPbkyl7i0UGa6UruAH8CjwfS4BW2t5sUYDohXHnmHe7FPU0youy58XDB/9JI5h7
EKN3z0EnQAzmYkMdwA1CIjlBslExHRY3o4pEBQneGw2upWYoe4tr+xjKDO8I70RV
w05Hqhhec9vKRh8qiGpXkI7fe6+bcbEe0pGOcJ8YAjj8f1WZI5uMdF1Gu61Zap3Z
Ld+73QIWKXSYNhc0nS6WCEQvw0wDf/NbzJNjewMHE+6Gt+YvDz3zdgzSb8V5hrAc
a+54LFef+w8J2xSQYMt/xV80JkqgJ0enBzqukts516Linzv4E2RAP54yxLHMkVr4
md6+nz83F5Wpl6lP18hrV7Mq4LYLVF3okMqOm85bGZh7yO7L8IbWwVzxM9k0VQtS
bakBZtOtUpiH5mBFkCx00aghXmvid0k4qD3QnIoWAarzE2Txho7woLh/B1xgGZ2L
uSJAJ1t5XMam3jFCqZnsEKI/M2CXT7+VR76jPQZNqvcSnIiU3H8K8akdtUTLSDRt
MjTChxq5P6H8SJtcTP7UPmzF82+qznKDgbOWBMXkBMxoiZuA23X6PVMwRb+lfxJF
ITEXiuMrc7wvDUSB9sMHy86e4pXthAcpQNmni6r4hMxdtXkv9nezMz183T77qpW/
4+pjcPyU7v8D0ygIN1z/uRKosbrua7cANIEanJO28kDoBlPbJ3jSgnPQAEAhmdpb
X6BlsBsyDN3vGjabUym/fChq06TPoSxow2YUqd7BmCWkDwX68uGQcMtj3bLF+kq3
JUS81YpertuTmnWBYDdFqStpkc7c8K6WfzenTzm7giaHNzTxJQMMDVDXkVTAbsVE
I1jxspbod9HwTqOG+RA2jqCgj+p2mu00RCzVd7jse0MytkIJYDjQY7GeUx9nzVO6
sanVQzRBj3l8Uex5hUSbMklgsmwJH42SCIMDbZt00SX5j9nD4FtxBuBATekESD6J
vZ8VYpkmbchPcklh/RcxTwOQcCvAQ3Dl2yDyzv6g6L457byRf74IIoXM+ZqYSVfJ
mcNFr/WGeglyB+bobIHkSrckI8dQUv0H9+kgI0TG/3BdZ2L34MC1owBtjivXi/IZ
x4UVzXf1+h+UuNxBNUF0GnGhj4YTj/mGf6q1ykDDixVUbv7IWg+3i1ttuNhll8rn
c6CxpJ/fvzvorg8kGO8AXBMsnRqEEAs5EnE6itCgM0tlpEIHn/emZWze1B59qek7
xysvIQyeNsuIhdypr1CRh4zaCrjwDgCK/In5231ErxJqpsOsZ2OrqVFeHKbodZmK
OpfwW3Toh+yqeIyFYRCJyw0QdUswAhz2BoIE2ET3A9ZcDMsXTI5qsbet9mXFUCb+
+u9t/io+iK99mT5JVWnQowwmIrPmj5hRu8eHIz/T6tNi8r5baN4cQa1LbvgrjVWx
iEqy1QDCjnGxexASyXxpbRSTmNdwg+O1/2kWenXX/lKnnCJgyDGh4smB8hRETzsn
QKzqOB+LB9saRqVPNiGe3f5N795paQ+1lvk7uSJ+/PDVfTKtsequ+Y/T3oltUSUS
bOWd1OuZu5JqadR/1hL63bsZJsrokTWo4IuVvmi/KVhGkTDqyYE620/4VtM/9v06
S2Bd+LnPZUjV/BewjaRVn939i3llCAotB0flBr0VhpB5sZvlB80TWICWXtECG6FC
ErAfFGOl7Mq9cZQNZRpgh4wmrhXome0Ni5j5+zuespkEBTITX1T0GlkLbYvB4gb9
m4G6jKNcXopcpta7zlS4fuxoFAwOOgx5kdpCJRlvaAnpo02tY3ZXjyEgOt5J5wo7
6WPebF3D9ZYfsvrxbNoV1ZNSji0R6fZq0vm9cVlQHoSWSQkKaknmOcPnwTlOUML7
enxBhFiBN3HrNR8lrh7vr/afHskN4i1kYMsKnoGbuzo6AkZOdsDdHsouu/3ITvhf
kndpIPTVYuQceYklsOBWZuOk98Is1IJKGC/BNzzfybr5DrMW19QdvotFt2BqyYMW
q5Dhr2GLtFGozhcu8opvK65hW9jLAQAg0/43OPHH1H4hdsMhKnJuWI5LKnQa+g5N
i5Yg2xGwZWZ3YmNeRI9mDtqKdA7/2Y+MdZrKnGq/tNWJS3W+Wt90cylZp/EbcoyP
PuYJYme1/rEQfHKOWVCiz1yQMonikqynQV2/Z5vA6PO8xp9XZwGeTj2SY/Oak9of
mA56P08Ujwf5/m6Q27hxZzV1/1PkK3IJ7bk4XyS0ejQQhrPZWg+UV6P4U7oTuIOB
2/aNuhyZY/mm2dI3CJO0uvO7UNoCTHSdcPYHb03J/U1yKV4AhX1sNvv14wO+mj3X
42/gzmVNAWOm4XSnCZSpD8rPWHsB9mHZiyqGYKeUC4qeYBhUYsLlsNIBsfs+aBc9
grKnLa21rCguY23wQEGPseNjv1cQrYl4c8dY/a8+ubAJl6b+It0R2XQViaQUS6oS
/g+rSNaO25ipweAdecWQQ5A/rnmmlpFNjZl1FMj1lLLIiZ/Uht6jiUipG64ukXTh
GUniuTuDkwG2jcU/kkjqu5W2BuWLEStWU8WlDHEzuhE66Am29Y/jQt5y9VlSAMnw
Cz1uae+v//btNnXnRKYS7n9QRZGii8oovGuhtf8Mrdk7OGHlrh+uxVWAjG8QIbfi
Ffjdb7brMwhsBdvbYKkTkwrjgl4LHyOk76mh7M4Uqa6piMjiuBQ16796WQowoe5/
9+M1INiJgwvQTRuq8F7AFnrZrD0E36/xkDFsE1zCNLbVtnkhblrf6R8GE+LrnSrQ
DPigkDEkvojrSc6E9c42qSxtz+LHuyyg00pic301OFD6WFvJb8bZTnFWXpzth9tG
7YWzDPut28396ORSqM+FtbG7AsAOLt32a2ofIbM4Qpetng+OKqCRrWVJDRTXz4B4
Sv/jL1+b2uUxotwk7MzvwsCzrFI5MT2JksTDS6NVBO1SinJMsRYMnXsa4suvtP8F
307JbeUjg/1B3spVgp1+bUv0wAH/sR1x6B9pZR/np6Adkh/SW1cXoTghtt2e9enT
B+OA9gXldgaOlfW5PiEVm0LCL9MoUtiWzT9N3aixpdcqPyuteKVehA+blDquiCG0
bkuhdYwuEScVRV647hixkfFiailqT5pgG2eRaOPPFvodHePkzEsJXbaONvWLag1J
priOTTMCbPuqzDdaCQIryS86CkjFCuqmDJ6PpwrrcMx53Dw/sVdUCzUxyli9F2xK
TNbvXkinwCbnW1RiU5hg8iuvpJSHFiuy21fY59oIFMkHvU3FoYjW4sGD7x1V8y+o
vtSsHDGEoIEFXUqYCmE/tPsegnrMJOOLY5GMh9kaStJGLSfhUnNN8jxKHg8ykpAT
JYivr2HKISSG/8xAXC2uR94bQDLzrcm/XwlQ9Je5Ad56jK4FWPUnbz0ygZ3UxWq6
XGQFm9ChTvEAHJA3sCiXW1F4f4n7gEfWw9dULFfo53MnBx3d1ySO81ebV/2uFgiD
JmgFEzPMFMVzx4UG4sZ3C05HYeansJc1HgwlDb0vEVvXwmsC6ZMImzYGtcc0Yc6/
lm8kSDPLpfDnnUo1vVfMnOxHJ6qcMUlP0s5keH9lZlLRrQ18KN/lTqQ58mcanIF7
8nKj4BZx8wbBV838zLiNcYK45mk03fdNeC28oVLwj+HIrcs+As5kI0expeyquZpG
nceMKTLNYMfXSJyHjds+ooH6zn3aGzOeLNLDGra5Lu0c0YIWaSZy5gBZN1UzMSI/
hSubSoDvBg3fugs7cw73sxG9HQ2OhYrVdtn3iMCjq6DmC6qhOreGcYAIMHivmZNO
ly4+95zWJ5k7gd5p66EqhH5yCHfYFD0FpkxUr6tohrqIanenlC/zPwwCg2qynsPv
1uXJXOPXV/Mi6ycmKZpPttNtUP+O+0OUrubeSHKxSBdG7Q5ctlV1AP1DvH8EiI4Q
gSqNfZV92vqHeDJP2+b2T38TGT16SBKYtIvzMAlNdMUMB6eKh7BYi6V2nOc429cU
kfhzPtoHEvT2qFEM5FNoWql+pXX/4r/ugUbo7313Ki43zewTvbjnI1c5QLNZWYEJ
pnPy7+P4Fq8VDTtSDOTTEXGJXSj3xZy63dJydbvIXdRrbItOwU9uiOJRFwwpI5yu
xI4ANRsfxtL6iKTZPOhjTlMEOB0TwyumwBsg1AjwKxtbCiZ+Zpc2T1F8pvjdKUZV
RkAQfPOp51MaCy+9ZZ07H8cn2WpD4Ks+V/zD2TKqIqPapkUaHxnhgLzzJEetM3Mw
/KEAtVCJhv6geJmIBAds8GO4capnMsWY3mHB2zrOLKxWbLpjtc0lqVDolZtJLjIb
z7vAxRbVQKrCSlMdI0sq581Rewecdeg23Ce1DxTwTuuiIwr2DjiU82Dy8DNoJJwT
nATrVRdBw6opWAIWV+TH+DTUrLrnowMVanEI+aWIw4E2gTiPIvtx9g1yQHgBvoIh
jhNKrFNNM14KG529xjkEtIUtUqJpWAKgWL3FGIBdjToSU4SJidq72WgUf2CBlAR5
GF9xXpENHb/UCIX7f40d9tRTjamWXjj2jb93wWmKoXmx+icybTHja6swCZaBEVsz
g8iNmFWY6+Q6hTCwsOdcfdJDIzML/ecdIw8DQrmGq0EQmzgQ6HcGbmfSUojO+WRk
Z2FRZOyBlvMoYz6b72vIMbA+Oi3egmW8S39RN3BslvSBVN2IBkC7ONjkdixbWLiX
AjFb9SaLl3PdgOZjdKWtKAAsbj2iEfHOYcG2nto7otqUXJcAMHkgwGoX2gVpynRC
+5HehpFRCkx0UteoML0Nv0oPEubfiDR/8qE6ns16CXrHAqNCqJHOHFPEVDgFsvxT
/WsW+kdWf2zZuYkCql/jG+8uy9BLA2hgocd0Z9kwczkc3WjeXcB6wmOtz/yT/9tA
T08sb0U6v5QHo7tTQvl8LwMIHDkWp3Qw2SShlVtCv1yhIN7EbkHaO5aBjPIUUtaA
xKgfwMXeNguKwCN41yWoTCBWJCRvpuS0KnJoeGlMusPqaZXbSCTB1TjRTjjuc39U
BsklWDRwSvSe+xfvzOaXHUztGwlu4n/48fGnWMd/nprNdXPQ5fd97lL7Yolj92Lj
5qS0rnP5v2aT0RZ+jm6EMcrnhs13hA/aCMyokiDR9SgIJGghRTxDJhYI5+ER8+6s
jzH0rF0wmPj3Gm2HfMlHBfipshjPSZ12cQhet3FmwJcLh8kRcudzGDiEamgFmtVO
+LSysHDeZje4smMTOsAoD4h6cP8MzsJhoXneS7ttVbYyp/vILcVCcV/RtTqtVXVx
0IpoZEwYZDDMMpmHOOzuLWjd1b+6YWrIhdCdX++enwcRmivSBxVMqtIaIUe+1KJO
1apapVNRASD9YFvcGlotlE7ihffrWD0xUizkO+AEGYc4MutHJpgEnaoThB5GuuF8
Ai2xr2bY7vfMQRnf/9Q9BWxZpEgNhYPkudGcyhekxj85BWC6HBwYF2Wj/XBCPuJk
b3KAcE5qRr7GDIpsp5HKCtwBHGxt1/YJFxrwTI5Qcn1koJ98FywChVb7nagOaboU
o07nTUU406qO4JE8aP9Gvclw0nbiGbwX0C3aEsKUD6eM9BA6sAQCBcHWBoZ97HBD
qFHVQvmh/qej9/FMRpbHi665y6XRtjIMu1xXglkSiA2EZehlw68oufKJ2DRqKWGq
8v+rizdTWGu6T2E4YUTD3kXSnednaoxiWJyQk+TAWsOC5S0MPbpuA6U/lc+HYi7b
bwPvc3HDDZ+LGyC+6aRolpLehhp5I/Mj2lTs0Oj5kQFSwfZEpERL07IVyvHfi+iA
/2uzO7l+7xvg7GKCm1+nl0C2tiQd0lgllRm2UQIhb26WsWFcn7LCp1laLGgp6y6+
Us7aoj+SMFRC/EmxtxW/IsxgnuiPdwPXF8wM79b6WfL5WJ/FihiCbA97mKyp6PVE
Jo/OSuIg5VrLrWgRULTT0mnvI7IOv0CSaPVD/jXJ7va9B6iTrEIcbZV019MKVmSI
8R30YIqSNR+IfL4UU2bbbPGtbe60v1ssMv3SIjP7rMPa03SGyF0d64ldptDRtVL3
WE4GHaKa0vHo9+ju+rgU63ovGL7vEtOEu5xHiTAPITFq9Txx/m14qGGNVqIAvOU2
hfc3YaEi5b20xhWdWpmtB5SnXHR8QQ1a0CuACBg7Fz6blwcO85tllg0dVXj3hj1C
r8EA3mibuX7AlRzvVWFhRIM/tlA1HAS90sZfGMy/qO9tlm4Kg0LJ7fuiqCEwHX6q
gk0XaedFHKofddThYunBaelqzIfnK8UlOc4rUSV2a+1LWhbkMQG04QUIYsTUI7fk
7Iv7bR3roCHGvSJokAIAkkajV10gEP8Qgc6GxBytNQeWAT9rVUwvT0JoNkWDonB3
YdATi8II6vWy7fEIUR9LWfF5TCARtQqAEAvw2Ji6K4NxHPJEN0KgT0bEnqxLpVnO
nV55Y1ET3Dw5ODlW7diLhUwn/HdDhyAfegmoFhqOzAacrQtxLN8aUqj9Vt4718QT
knpOM3ehCGmv3B0MZDIkzMWyZgHE74LcPMhVmirt86gYqCejIzy4UIIMKeq8xtRi
1bEjK63To5UDOAOqoqROb2yChwqWWGbQpDikBoYtHvhKBBZBZ63fWtR2TTVERcTG
fiUb38g6VmjAvyjw6UFOFzcSDLqDKvwm9qnTWOvkmyZOCryCl5aAQ/XVSQhSSyFN
j2D32PE99OmtXKS1AcwCregBnL43gReELWvTOmuBXIKCxle5DgFqKub0LhFLc+qT
uPfJ37MHjonaI3tIj3Q/5gBbUXxaQkOW4wJ+hVbyTcihL/eLTVlKhz1FqKfIF7Br
FsKr4guOhbtoKPsnumqEFjqNFGi53wWRpcu8CQNehJeQ5V4sNQN7QWiBD2yK3+ZL
trWpon5emoVhtpZvMvkf/FvwNbf+PvwFanxvKl03Rztnj1wNomWdkja8NnbGfrxD
dWy69Qt2iE2OLFtIkF8J8kKhxHdJCfCLG5S3Cjt5n5Kk4EUVre05a+dcV9KhpgFi
Mr6x9/tnXYZS+wysGBTHWxmvj/cnHW+l2G6Czkwjao/2dK3iwGHZlI7zTiQLbrHM
EfOXcxGDFHbQfcxOVuoPs3QdsO9FrPq+kzI/sjNxUAr2lU2SihXB2oThY1+Fak4H
zIphJ0xGx7iROWoyPPdQ5z6fpmtPT+uCk9oTmzPTHxFWmKZ/Ye0eaWUZ0EUxCZ/i
ZoES03yGU7WD5sJ+E14nIknFf16oahxgnRH2Gm9LTGZug1S2xHm9w3OszMf8OK3a
dEY1boSCu+QX1YnTdnPfhKEkB+N6PIMJy4fEmPlSykx4xFRn4T74zlGcUb1JZyhy
fnDsMKDMsaH9PoK2j818M06jQmvXU8wmNNYN1kWuihqBwFBXXkAqNV0QbF9YZhcR
8wPaxE8voKEW29jhBnWN/b2CVc4+5D1P34v5oDt1ULe7r6Rxb3psurPVbYDYxHtE
g/73b7+hiC6xVIwylwEoEbjepo5S6VM/+0fdw+1AgQCMp0MlkbrIffGgJUgI2QIs
q5I9cWFP+JJ0mzwTgkLt2rgldsHZhMu+3Uzj6gC6W6+hZBFq4PiHMhBT4CcykQA0
2I5VMjoa6nDdJ1o5LvImpJyF10TCYkG7f807wg32kKDYmCzUtCvLw8li6CmF3XL6
gJ7Q80ctiFOzNNrv3QklVf2N18kxxb0Avktv5mSN+LBL6n6cu1dWg1sfufEUfShL
sSUprnxYtnOwicnocQZR+Xc4GAsWuY3u2TVp+Z4S0PvuAxpdaZwPZXc7h/p6i2l6
IyiDjF9kh7kZSwUVEAN013NoeW15ozNd3g44BfySqHwxD05oxQKpKpelRENWdMB8
4iksf0NjHWMEqcJo+iaYO/QFSSJURlAGB8pPkfg66QVTHXjj0Ok9/t/GDYVYrib4
627c2vl/PSpSllsVo37hOD/GXa6rdBKMdDaN72W1WSCKx8DojjM9ViljQTKex7fm
9127sU+ic5BQ6YKTvX5dm6pA18doKdmb+Dn5fDgQFzcVoSqyCs2ulAycd8iSNEnO
+8Mv1BEWxOnXTEVsh1Yz7ctYv/pXTtWr4tuCr/GffuMCBDsK5QzufqYx4grneKwA
gMFgnrPJk5A3kYBAt1lMQb+1iTUQP1tKB3Zfb9STtOTaQzHWqe+q9BEQNVyZ7E1b
rsfpzc7vQsgPZlNA70UKXrNW3RptGbkOyH3upS8RmnmdA9mQ8RWZI+VkrlUvQoul
kfsDFBSNhnZ6ZvnKZK+U0GbglW/oSk1jjHef/s0zcuWJZp88Q5vM9x3k/Ul/3U2g
KK2PZq/KlNFY7yoywvnKHxY8VB70x6TLUGJKio9uXkj5lGzmDaHT6OxCHahp6WLX
Ij/rFS3V/fjA3sbIK0d+cfIGYFEWn4wsJRIMIybZrBl8nBAtbtZXhiW6hJuiWdKh
U8ivPo7q08WCyVO0mIuprhnbLr6kjj60XEaUqL/PWEkKmzsm+fokKmFa6KxTHWHN
1B3f3IMkfXALxuQKo2+A7nbSJS58cxEH4VTmg9tYuJsCujjWLhuVMeKHPTBXCThZ
C2yhCiFHiLjecj/xaZLBJBDv8/UHJ9fThbVpG0QDy6UPpQ/zQ/eDH1v4b7MB8mli
ZRmfacjpJJfQLd9y3cZ1Tl+XK3plPk2s+OJTtRXAyJ3tv/93TB0dOFjF0xsVO/ty
dFrygCQTBJqrDVFRga3AQbhYOzCqL7jZuJW42DG79FBthTjv0UGojteAOT/ZlIS1
ikOfUCEbGaHBYdx39yDU6FtOJBintHUY7g9CDWNf9KORaVsWhf+ScLpKBCAd3KIS
MAosfBwB80/ZxbB2kw+U15hawhoh29FpjgewvpHqiKa3qwIFnHCzXrBv5ynsol5G
nnwhsS+00R7W3dMOn52pRCscUTb5Si7vx/ARv3sl0Vag5LVxPFuhFxqgrO1M2sQn
/abS4QnPZzY7xdYjXbOmsa55Xv1XT628YeTPLOZZbZcDzJxyDGfJjs/Ce+eXzPrg
5W8V4o++3YrW2+aS0tZVoGvbqtD10TIrGPqoq3gUXx11+o7jEwDmqOXlKZsvVmxw
2l2684iRXpAwe3rCJ3CEs9hVZRr4kDzZUyrGJmNdrlgjiea49OUOYnd9LgSLCpV4
npGDoEEASn8U1RVmm2TosrWkYLL4Hq2Vnq+HpHnzT4vpm6SpHXh2JGB4DYvo5vX7
qhbep4sEcdRjiX4mvGmqbJ6vaAwMn8Uh0VKauXpQtoji1jQHiOzxSILQy6pFDLxx
QVPkrmMyQAWMjrmHlr7pj/6X0U0zE1cFygj4MT+To49iJXK/aIn4osKTWZhwsiS3
+Z+C5wnL6re5bT8KDxAZWkEpcnEM2wSKWJ3t8rGZeOoiZbv4U0F1G3mXZhoi4gw7
3LIDHAyqO2yIHegUUtpuIhvR6RaT+rExvWl1vUmD7WdgF7pT3/LM4InntLQrL0jA
RxocDzOoRWDBfBwB8V307cLNKiEy/JQ5LV6rY0114IP4NjNvjb8YENozO1wVY/Y7
e0hDJQ1rnaUm6NuaMkWWeOT7/F43evfOA0TVWXT5zhCCh1KteCwYquveb8xjhL5V
rDpyXjq/dmcudlhKARg+lVUotsVLNsI5qoKNBRrtbawpIaGVmXLqsMr+g21/IaI8
nnyTxl+BuWS/LGYAFDFeXWC+4coKWd7QPkeStjCelczSKLFUoHdN/3EwtT0aGKFw
rHFly7MyZfa+ZObZ0QegezkWUbJjrV4m9r7STba+myR+wMyS6JAD+8t7jlNgo0BI
ns2gNe+B8LutSH1FLBjHmTcy1iBTmQz68dnwpW2IDo2rfsWefqNKjWsjd95NVAWM
4Ny1BqH/IDhrXziylj4fOrHsUfCg2GAy1WquE+bm0By7rsf11potOuZ9HOspsw3E
Fn74afvcRp7flBYb2IvF7O305/x3vlQleBgBHUhF0BAwhCbjlQwVXQcg9df0tLMy
zutQppxarefq9dZhUCQBgLtY7gIz9R3nv65dPdzwbvd6cpV2rlsU6CSLJbbRR5W7
A2gn5bKiu2rqEGY5TynxK9Ri6bzJuJKb2Viq3/UePF0LbJ8+9Hz8tjDrsCXO01fj
xsNrLlomMDe39ADprLipFzd/CJz41m50Gu9r59R0yW4ALB/7zQ2wGEdbyRjMqEQB
fPdxLaCmY/92GhMBm9ti5XPRohh2BlNzr2cYGX+BE7sKHrzpc0e51LZau7TOXZ7W
8mrujHtjLUmIfIgk0FfJD6IlfL2YPVV1WHtopt383rOvVWJzmpdh1ocdrF2/YoJ5
YrJrnH+jUT3LaXfQsYavmFUS8Dxgj9yhc1XBpUomEWzUCxsFBDq8bGLJubJ9g036
wHdMCuHAArVBMkq9oBfvPMNyscevrB666Jk4rPdcviS9CBht/f4NAVROeS8of7C/
BJPylRMZtgXWzDPqDJNPQtewoRYhqm+EpUqNBcHZL0dPeRhIYP+2AfDtqG3qhIBa
WZHMGGlLf0nnD+whkuppKxhA8MWFweggLGIq5MhQm09zy1MMnJDxdf94akBblNj9
n9IFu+PBGrap17Pjy3/I80CpqlQIuA5zn8LeKL5HmXUIWelEF7mpVqhrYb4tl6er
UQfBfDYSwzGcN3rRCRGqnGptNbvsCHPQoIzJlDd0CqwTt+jLL0DDwgNpm3lPeDfs
kmCRBY0nvTCbgtnZDDMdzCycizYsOl3lZNSxR667mNXnL4xUbchu/p6b4gNWyiwB
cE8O/wf9Np2e7uHyUtGj1juH8zjF5I4+71f/e858YTPtng4KbQJSe0VM6a92fr6L
T0rLIb6zxRRTnzQHNdBvNHuIZnP0s90BXQkfENS6DYAaK7lRvuXDRFMeEK9u+zWi
4KOFpSPd8kjNYj0CNRriwQgt3ssmNmp95Oi2h1QWhiB4a1wEr9iKxxmMvaAEHKOs
m0pEXnFmfYr8cXZsqXC0Aa6YwZ0LBWFUyrEuaWrGDw+b7M3NYtoy0lOHogOMSfN6
3lg2T26UfRWC8uW5xENBuWe9qaH6snwV9+CM6LfPpzv5e+gJK7VriL2BIQy9LAr/
s4MWN6P3JAq86j7w2w0xa0fneMpx4dQDdOfOjFY9lOHOOM0zGeqvCKBMzDYwwPYI
8D54zYlUUfRji2Sqoo/FNboZD6+W0pJ8l+OZyJk3+xF+CF3d1TJnxMMS0u9dWIkM
kRatPaVXfM0zGmTXe71cZ0YJ2trZMkpye1CWo/4XM3QpoqxrYliCI+dHI7SQvXpV
+gFGcY2wuMuARBmyGZYnJ3b51+427GDSx30l4rhDM1MI9szIawsLs75k5rA2hpc7
qk5ZICDS84MIgFtDLV5j6uj5go8i8kY2Futu9oBRuB/78oJklDj/+MAHDg6YQ11B
xzyLWGBzve6/fFJG9O3uMVw2NW5CWMUOG4JMUWKRB6YLDyev5FvHGkWEVUTnd/ii
6fOjUOFdshrvAcKaKlzDFXP6PVQiseJCGu89RCp0ZRJA2KpjCWqhgTH3FHkQu4HN
dtlXgCmyQin72zD56cuE6mepvpsByypCyCZC8dEYYvsLss4m0bXwJVq4TLwV0ZWO
zxS2C0Dk2B0w8nOYLLGpE4Dkr7czIIqqu+us9HABzj3fDz0yisakCKoWAFhWbp2l
W6XPLGSYPfho3D/VNeZh1kpXqMDPfoDkoYflLDC0Pkiqpw8znSH79EdhrbLHMZS6
2mN1y6Bx/DesaMmz/xXJ6PJiRbK2v7PsVwPu//dAmw80tN6+7Uiyyggxc8mt8IdD
EtHqR8RW7aQ0MrN9P7oXuzPstovZntx/IBqr5ESOFMf4IGFFyHKVE4++61dxuxV+
FP301VPQ2lv4k+2TmuiYUtdSRwMq+4R4zthM9waH0h0YOA4u7QPXUtnhzhRApgJt
7UI3s+Z9XxH+fKYRFuyiH8trZyE3SH1B9FnwhUk3eHGfdVZrur4J67d9yGj534vc
s05Pz1Pc4pfBHcffunZBeqnGKX0fMGxjMWntUwEXTyYC6FpibbMngnWy2+v2L0sy
QOryuUZNpdXI1oBHGBV7BT6xDZBO9csuK7BAhLDnR9Dch8p6n+dgPca+SOH5YNrm
KkT1++PWnTy/NS5bw9rDSjp8Ik15HXsEh1sRFr142cq8QYE08aBAuYiWpDRQPBQx
aHZ5vASy+fS29/6HrA4ToH1L2x9PuP+2adlGctL6QxuERxgkpZjCgM1rKkBhaQZW
pIiguYGbUxGIQBR6o3lm/CKHpe0441EZMS4RHb1bcpBcHGhnO14fobNv3Bka1vi5
r3UAcl5mVWZRSSWmseHxdgXTxCoL4JkAWQ9NYU4YAEMmNtDAKgpTZyiDwGfbYp5z
YydEWK+zfTDHaneCl7zQrxk2lamRp8zwHqZZe4LCh78PSO0FWrY3FmpYjjULv7QW
VkwcL1GcyZVdUQ71EhYBapGXmcxdHDLdjTIao2aHdDJm59JYxMCBUQHpcklLoU7l
qp72xJ7MfwZ3p96qiALwlOzJMhHYtazkd/IkmSIA/VGk2KSlt4N1PYlRuInPMR5f
piU4ZeW9qkyf+LcYq6fVUCRx1yJGfWhioR9YAjI+SfXaF5jci3zsnmaQ4ivsVv2g
MfU7k9sBpDmYZ6QSJ2tzk/PmdXuy8dZX2rlRcdjEhI+5GOQu6BOf4aoj3iVL8NY7
/PbE9/SYwUO3SWHZCk9J8Lv0dV0cvANtJeTi+M9Hynny4RDHHUutFI4vtjRZGlz0
Zb77OsvhsTyGTVIwLsi+o4Gf3rFvoVrUVNgwL26Gv7NztJbMXCtwU3ayViInwgfW
5UW4CdpKJRLIf6xdK43xukZVCQR7KR6yaJii91wUzUHS6m+g198QFRzwjJVBJncP
VXte+hofg8ZtPRBoxX8v2pqYQWRSomJhYX2cfo8lYGN+rNQtNrfusrr8j7wNCn9U
LUVKjTsrOE8oojLHuGpPV3xdKsi2NU+eJIPgPeY5LInPpeqefiecPHnySG0BPCqb
OrVDs9NilxJ8k2fKmEVtwPCGKYxEfpJgvlu3zWtdpj6TdAFvl2yTi3q6v6Pk7Afm
9U59kXBtPlwNz4bLz6RwUWfXycmmjTTyM+pBvPpus+oo1+ZhC1zARNrv7jSJGRNL
zsVTI+Dtv6cMw/CYt090idpBKhtaGQDsxHTCODDvi2RQke6wUDXO0Olk8a0nwJEm
HfxuwzCxQmDhykwQXwQNP9LOwNQykMRYFrgBIc4T5g4Ns4rDkBe1uqEGrWjxLeU0
6EAJGJM1iGtJeDcFiZJEJwAoO3BtEdqMcPrQeK+rIwBTMyGxus3TmxUPVFUtoJp8
vyfnT+ppCT0xnOMjFL/MKmDmzldui4oPkgviZOTKbxUylQ/LPo8Spmvr6vBbRhjt
7mUXCB9vRL14/wZDTnrS47QF0M8HAk5oCzFnGqONQnctAV0Y25hALU1lXUKKun63
OmCZDtlCDi0Tqls9AOLPRxwQXeFyaxrjVrVKou6X7dYbS5GrXrp9A4qAm5VLdBeO
ZqnZqtKGwkgi1EEcPwIXDHRSDcfqgPg6whQxtUqO6PIQB5r/yeiCyuO9ygbKEzsH
CFkJVuL2AYmsEG5dg7UQmX+h8R3sDpsDJrdzJ7bMe6VQUEl/ZdnKv050b47f551x
P0uPGdGvrrZhIb4NMhVqk8BXwXqRIVzjAw3MrlnhyfhUGnL3tUy/c+0/n/Acywnd
VF5WPG3KC6A5JfQjKL/BxAMBY2DvIS0lgruptlzm6ZZM2UBhqGfx99b5BI4onyvh
/wLYYXYTmG/GE1CvXcsNumI3C5Yy0ZQ3f+JwNH6YPCh5HGWE+rnjSf56du3EH+wQ
fD9IYrbyxcddNaxE+UCcLYc/8YsqC0cXc1FKGz9W6E5sAQzEPPmF1c8gLJ8gg5MW
lyas3BPryO2VCQTqwZwLnSdfOBr+7eXTU2RcSOiJBDKLKk7nZRfUKVD8qLZEU+Od
HPRH396kayArdeAPpAIsf/xoN4Yy2LOr0gzhx4U/hCqAXkUFAKvda6itu/9QBnBb
komXOKs5R/V0w/EUpsP9beUIBKgE0KKoVtKzGMhDcwXm9OG7Wcd5projw5vLKN+C
QzO7mtt3zlB4OyGd81xf9GFFl6+eK5jw73a53w+l6KPYi156Y3O++J2Sp/CKjiuW
GZ0RQtgDK20JMVYGOUuAkTRqWxD2eos2WgavoAQe0XUqGysxIjDe0K3uMNOSHYl0
EFYLkHs2m3Sk2LOtNCjsyxPDYIFTIxIJJQpxtix41a5B5knzlB8Pma2Pvi2If/GF
e41NY8WPT42dpn1mubcjBjkO2Wb2wjhGg/qLZ/63Z9WdZAHAXir9S8WvvK6zxkkc
lf+9QbPzWdd9XgzWkm9D1YBZAwRla58sqwbKqXtPrt57cQEtwI2CQql5AKQw1KrB
5EfRH9/6swUG2xwy05VxCsbp18gpURcHoEux5eTyeqC8alDf0sWzq+cef1dRb7nK
z+OCJTYAO+EcIEo1b4eW1TEJwkgC10dIDJzkfD9Ce2gTT8CakXqd2Gz5LHiF4qNL
7h+Ys0EKe/98MnLGU9vPeZB32JvqCY3RXdTJO2IhDkzJDhEs64VK1dvPFXcFyBRf
CCB9I7GXleRf7evJcjtl4JGtNdZ6xoe9gGYA2mXpRAVdGd1yvLj/T2TGacCcOu4T
Hax0TSVDi2lVObnEvI7vj8G75NMRM3E7wR6u/GPLfN5K3UaydcmkmaXkgt5MG/j/
MuPevU4vD28z07SPsLl2pOgirfMzLer1fN7HDYNqtIc6NR8ICo94v55ONGM4qorf
2l7RioQrYjRl13G0WNuImLGxWTyO0nS4BB4Zxu1csezlSdINGh33oRrI1r0SM9cm
GpFaivyXnThDPfttasVATq88VymBIBpSJKbui9VXDCkBQ107JYdRh71f7gtIV+b+
9IDPSLnQyA3nKyT2ajMYnfnoxSHGwBarXn9TpgcbJC2INCB8OAuux1c4e74VP/Za
9YpvHHkGR3eUVg0yjcUQKiBnyhpMTNdGk987AByOyvGhP6qswOER5NPjbSoFnLK8
vAUP5ULo9Gsi/WDCxGJn43jJ6gr0NJVE0vYcoTg6FUyEfwz7EouqeAsZzU9NDyAP
aSZBNCvg+4+s3kQizDuZB+hyJD8iI+w+pzsobqR/DDW8AoW6qpss/ZA36r+bcGdy
dwGg2mDavFOCVPcKbNRGr2liWw4xy41Ch+CicNlrWdycaFQ0hmA78hTuy/WehS9E
ijzVPjrI3p4t2vWhDfoolNmDd5Wn9UMfLh7ztDnRfKG6nn8INwPsePgvlf81p94E
kl+B02P2ukDKPs6by70l4ELOGRf4D2DctyGT4P7dF1RC6xUEUsQLrs6+nHQ+g0Tc
uXBFSB+erM53fA6Hvjc/dTtirVCeFuc4ghO6j2+YZCcxVW9vhEBSVzCHmVxc1ZH7
9fgQX9maO18rSp4pwvIAD2CI/fddl3mXYTdlg8zEdN/QK764Ril2KVWHH5eyMRIF
EzpAbIEVTwwcOFw4vtQe32FhD2I5ToJ0EQNiXvE+Z9VtgAqatJXiIhMHSZ/m/7CM
BlJLV44CYUVGjQZjc+kpaoKfVdw1WPYbVSiSpxXLMIgodEFE7OQEukasQFhkTvnb
rfX7TujdPHMY6MVLOLBaQqe29YSDSDUFuMSvZK80WIACmEXf/8W+WppI65p/lg7g
7bnAG/sAYCIC/VKv2589JSBGgqJ+8rEnNF7zGgjavQ5ZAOuazhU32rvwT2ak2v4x
gt2I9HXcW8OEwObUjJIay/8XcsrDiKjXD8jOU9pKAZ1LGzyenFfjFpnL2j75tROf
djVSCtCNdYDdYzTio86rRxP9EGZ3YabWrv0qVhjunSFH0EQl06OdgP8UOhgmqIy/
9Bc5zgBx7ZqtH/Lq9jisM5xphykOxLN7Wg/7ug7Invl82tZvILPkKaW7RS2li7ll
TWg4gK2qHuS30Uwv8DHQNBiDdZjsmuiH89m6gfJ4wS/xkyehROOT5nzaqEsRIjP3
U0KwLKmpNG1JfQY9tPb5Jaa7DYGywhMa+817vZ8D0etCyKgHQsXX2dREevHNJ9oi
N3XubOnu7tpUOpB1yaGrhoxvUMKCQ2CNM2NxxRXVXSUoqnbuF0UB4h4vdXngsWMg
LbI9pQ6D0LVGGfaBL0RKXKz988bsH1CZmWjP3MqozbMTskdAflLOOe5w60Zm7930
dX0zifkBPoepm9mRo4UlOVHy01Qq0JuIyiMe+iGj36yCbIsL4si3qHtc00LsMCuk
C1W+JdsZgjQghhsY8WD6scSVMbk/r4C5xejHuvPjAUlUfV+ULTtTpsUPlEvdLQSC
mEfRs85PE9as1c2LqOg6kplKQ2TB6gsRC7ZMArRAEpFmOSMW1lMSBr/HnFcI2PkM
eMagFyLvekvsrvNJKvdUhD+NaFqScZqXs8oXQVvIYyvbV+s0Tm3iob0L3iu3r7TT
BQc5SlzcMKaoz1UMKjp2Im7qFXkT9vNIRX5c51tltvFWDka2Kxh8sdyLBvW2/Qb+
RK7/8JaisbrAQkDlGAAHkiiUP6iHhQry0grtFHZ9IF8uoFvHEC74d4aLY8m37cHd
U9poCJ5sOEsi5FTskc18AHfUpdz8aOSF62uGG071M0hd2U0kofxuHvHOjezbV+Kv
ZMPJCFsiCX/Aq0FKv1sgYVP+5oC9hre6b4zNvBKiXY/7NDhOqYiWCn3ie/Khyuyp
zhqnaOZ6c5v3e77Z/bKvhowFw4O8Ftgw33QwrUMr5kAQauRtw62D3HLCh0GymNmF
J5v2aIf5fAKPW2TS8GDDcfdl9LG7t+CQXlY90UWeQcZqX4ZqR0JIa2sn+R2G2TX1
7gcOV7hif5HNawlGHpcxhtMhk/gD+FS576f6NZK54tZ7KXUtB93g5mt66Ll0qJyK
ZIPRxViHchUZAxST15xID52F2sfo9BETDOHp4xWut2ubjg1K3Sz48kXNxrUBp7Gr
520tDq3JJefaWeOtoz/qgYq3U5hGvWCJv11V/4mNyNUGJT0VT71zwAXtM7lqG+go
Yjj8ne6r37EJgsZatlyEi8Xa5/3Ah8FBuDICOpr7CrpzRHnfs8KBarq0AHUz0tgE
caFuNA7iLtzU4L8fQGNFRkDdoOYNlMKgskFOHjRQrSeivTEZg5ZvS8dRxBkdqRiS
o/B6EWhO2vEwXIq9ekAXoQSl5E/EnM7Op7KGtwhxczItxxWzR/8szORJGD4Mb4VN
ooNZ9m3kM0nqyBU23lALAcmGK4y4jSJpVadslMSfbBOOAv0SzYoS2zgpD0BI0PU1
P4EXsvFiVpZOZbfqzGmXkilAmDHX+e1cGxBmihHOdrogZsXemBSrFmi+H/yscJBT
YTQ6TB8RhRCu3Bl3RHWL1bPlTz4oUFvYz2IzlKOYd5d7x9LShuqq4UiODiCZXzSa
8wJDWd8eh+2fzXRQGay/A6/fIFfaZ6EwmW9S6LnAiyYdxF83MlS7E9uOoMFbBoBk
P5T7f0lERf3uCscebc9Dgf2OcDM9g5GPZ7E0KLX8iceatdpHqSAf6I0IqSZ/U360
bkNygWYryckLC6G4wXv8O6s0dUVhxaTpYzTM4VhDqNJdliM7Ok/rZvVFJt3e4CuU
D/U0BeuCNJB63wSjtlY4hikNrkIyqZVbQx3/e8K5dNbN6ToOtx47I/3wjKOe0ajB
DxxAMUsDV1hwR65KmZ8Jbtr50gZZ2NAjYTSmg7Vh2O2KrxtVJQKgyqrR+0y7fT1v
hJdTqtiCLbNkAqlDtNDqjCftdOvhkond0ob3/HcjXSymEvXccqLmMCg2Mnx53aHu
PkuaJdN6gvQW5BYS3kG3osiYwILNwpFelespfDEOdEDwyBAJ1gI9mAQJ36kIES/2
Ba0aZEnPEGwexBeJlgffRcYYmYMRb0DJT33W2qBbAWhaxscpr4azvLgZCpuqDZIT
mBSVzxsvDNElw/a3XJ8Z6N4k6NB3D8osLpMnvgKHzkuuWD5Zpm1z5ei5saMmpgyw
QM7lWroHsk0kDlGZkzxJSAKZmKH8h5lAkHhXmMgdIWjiFw4VaalRf5cTcflMNvuH
5+A5CNmcNh9AajLDr9MmiZD5egxXc2hRlQc9kMVB8jkrbR73DuVoAGn8Q1g2QsUb
pmtbYvhaKNMye7fiWjpIC+A0ky5WhSa75fbVx29P2gPO0a3E9HYmHuGbAV98+w1M
v7TNKgMvF95OG0jdr/e1s64FXgBTVrbkT3gtrh1cfB5URkSk+EBYukfjTt7WsNNz
R2R7CbE5iwRSyZpfFLwJfmpB4GaCf9wl5wAiaii4HaX9Pn7VJLbvio4jIrFBeUZr
IBPKiCGIk8NviJnMLniM08pivoVYaGi7CNoT7qvtHdkSjI+xoMurZpGjzv3+2dt+
TKgskNUvXPadF3p0rVINzMxF64me4OmWfgzahHqS0cwIjfkVhVqe13WZ/mapMbpC
jc3cqif8ADYxb763YS9BvhgzdH21oD2TKk4OcLuoGhYx+bUHEkctdKmlXVBU46Nh
6kWe9du7FLRbXtKakTBmmJY3Q6woIHJY8DfbJNx2rowSCxRP1lmym+ZRtFCXIuIh
J75LfGm2pkVpRjJkdeMAdPzgz//A4uMXJOJ4XUaL29syCprYhhHGosyH3tszpMTO
6pVw5CBmqspMH8bDS5TGL6qMDmthEYCmVfeaN0Ou16G2dO3ThAM47YV1uB9qEJTz
iUYAwPq93CEf4ffPWb1w2Y0AJ6jt/IL3g7ODYLEN1RQgKrUNAs0Kwo4Dv8JJEpoK
if7+ATcQtmp3F8rISPvFqYrvpX+ziSYtEYtNV81tINlex5MsxUEfP7eBuefGbkyC
rmOe3T59iSEMXeUqY2Y8jFulZLttOXWm3syak01mApnDEvOMr/3NqaOZyhy76/OP
VT6N4PdFIgMU87yN41RePkfmOYWtkOTQc/V7BscEAJ6cWjMCIMTEUuhpBNtcKFeI
CmgwOUZXZfWASFFfNeuoTKRJcQI7sBhARWaRZcOsUTn1qZga5iQgft6RtYwYGSp3
GeJVQqNPHgd2l51Xto4abrLDmjJ/kYhII/JQNqU9Z7dOwMp9v8oBA1R+wg2GDBEf
bYQkhiBm/9gXvXgK/aMAhif2kiShuDpowkK7jXezysRhTpvvKN2A+ARRu4sbVCVt
bPcl+0RvcIst8XjXpsaodhh0ou9Yjx9gy/uTuL/FALlNwl1PIJ0pO88sDz8BkeHA
qpiMsV25iUDoaxo1t7sfkNlJSzhAqMsxyggn50K37aZOHlaD3AikiuDmQAkbsLBO
awOgorWX5/i1ESoELPHxHz7HxURWh6bOm1IsvLRfAWmsIsqcqc5wtZN+C0pAFz0j
va+TbMWYmGHN0h14iVPPchuxYdBmHYp+BsCtodUHk/zoIJoTQqrnsw1ZM+Qtz9Tn
ZWexoy42kI9ML0smSSKEnr5c6PAK6HrojnlwJWQxXscICjxJOkMBmTf2joShNszA
1+dQd1x5xu5Bv0UoiJDjQT+dJfTQLw0HZGf+QEnQeWEX6tc40wBDcUkw4Yj1nCq+
D7pxEWVoEIgKySCu80MMtBCaGa5wI+t5SosDSPSAVtekMEkItpql+cfwVLhZyX4r
Pod7dx2g/WfemgU5SAAN+UxnUMmqEd3oJbfQQ9yp8xlvNYTud4iqkBEtGItuyGtB
Tc5pTCV3tcHZBvFDYxHjHW/Cu2rDzP92TTo2uTSjfwAsFLbzGdtcFpNm6su2wjwh
WHFFW5zNo6IQTt8TJzR1MdQlp+lUhmcDhtonRmhbx16UFPxf+Or20MW5A3NycwgP
aYADbYioYFy5EYaLk3wxFyekyLobuagNe5Px1qnKvlOibPZ2+QtYqAZFFkxrzOzP
yYN2CFEmqandA4eFPExINp9ec790nFKw1bHJPATuqivv4meWg1uxIlX/zFq/latr
73Rd8vdfqHkSVvRCI5H6CRocdvBVvne06V2nV+k5y8NNkwTQRt46/81PGRrGNofZ
JDp6bpWZ9YWzs2pi7TfPYhirGVuA3QSqs1eLyuVLSMB4d8KjFC0IvKcB3StS/Dcz
wctIy9p25m8wSuWpWVg06ZYQctlRbnqFfdJVGmkt5l1Xolv0mj1KZajcb+RlCaGC
W8lvjLmr5gvUxzZV2GpdQYogd7s/lm/TqcdFESNRJupJo3um1TXoYdH9175m0l2p
44o5XsCripnfPtxHYZEer8JOE87N8A1Ld8YgCXmedWq28h7rAKFODpixtfpMQKZm
0FoH3/mrYltS+NRTNbWbVJl4nY26tTulI6Q+7QYI40knx/wXuWBEG45QpNOlIYUN
64hqVmrngRqSlazX3UQ8R2Bc2RzL9yRvSW/Ecnbn0AsVf5lhFjhcVP9NiW0QGmMg
40WkvkjD9002Gy5ao1WOPX52sARMVWV5XO393d4a99ysio+dtm3UlRORi0hk28fu
o9bvbN1X5dwzL2XveupHQKjjqvukoRbRvigREDJOsOe7xkdaeuaVwcobgPEYwQGC
a2iOF2aNtSgXklCy1Bp1DPs1QEUZcPZpeO5T7at89A4LHr9zKg3N+agfN+uuIQBu
aIp0Y//7jLMDPuS1x667EQerXMr3C8ERXNPUDnFEIC6TEvt3r3BorMO5J834w088
ugNzzx8YUyQt5z8EuqlTtkFpfaFZz++d/e7LNa0hA0c6uyQXC5QEv4KKRKFfEZyO
pVUoyK3uTxN2ip6KmmuDlsgSq7dj3BMpTo3aJDoduOl9O+VcUO2XTpPiUrFiEiv6
e7mJUoxkEKxwF+L/m1fZ7RrbPHcQ1vKx+yEbBgZPGVXh+QEIkmXJBcvVW3SM2mXM
N7iSZptpFvZM+kjYBpfzMxlUbppaMkCdkUs0RrXrpfzMAbyWBoaS6+pDYs8GVWsu
RjaSWo7liEhtDKEcJ4QOzWHss4DzNi+xpcPpEBtwrt4JS3CPE+fE85vC0C0W+LiF
JMU16Ih2Lldxobvgx/Se8aqo9KibKkwn+efloWQAwsEmAsEoHLxOfKK3tZzllDPK
kZ/dyT6fhOLpwOEa3EHeJBGMJGoD/F62fEXCMdJIDehg79agmgAGnbF34/IJiFMX
Dcwk7k7CnzoRIg40Ejl+fRrz9YxYEH9MoGvVHlDL2kunIA15XR0r8bNTi5n6YQa7
44e+Kw0A+O1Tkz6c37gWJI31jTufce4XgZF5GikzZZDHP6ju7cv/srqOz19aqU3a
afj6lngbR2N4R32T45eeMZ8bw2cro+Sb4f/ciu8cwVKH0MPw9W73ddKdiOhKHUGd
d4PNi9vnarbpCdO8mJnVgx7dEldSqlVPYACEosaCJMeuhKdIgB5hc0iY3sPkTeY1
l60fYzTG1pybz2fS80LJdUCQp76AlGahpNZVN+M61aYri0w42Jn9JEK2EyfEe9Rz
xOdNuOH/BWXeLhdGnBDdru8ePJvRoYTSSwziaHBshrEhyA2sAzV6xDBBDqKyX0MW
3Nw0Pfc+gqqLX+qQqNmFSYV3uOEjPcxBgLCoKEYh9PGpspOkZUnYo1Lhp6DlTlWl
xhW4Dx9QRh2Kzh245vFV7+Os+K0tWSxcSTZCM+YimgGDBr5kpf+1NyW+XwuRzuCY
edeJkHwb+qdg43cA/uSv8hNiIOTdkIAm1kFkYuqNJwnkwTVI7EDV0AVobt4RVAVh
Jip5YJPQeY5zMuBtxJSfedhjeDQQ+wPeE+gbebj/i/iUtnqOoJh+XVpiNdmeK/Mq
BJfoK5k42DShzz9oJo8+LhUo7XR5iMJgHVVi87FoEkT2mbetEhyuT42h4Q3LRTqJ
KrPCMuCSBoh/dF+B98SYzxCabpFNAblSGyLEOyoAreDEzA/kTj0PP+rqgv8Uu9hW
M++bItZz8VwY9zvog5vMh8tIhhey7M0OrsZqFaRjxTkEkgvMwBtaqW1a04moh1px
IMmjgfh2BRg878P39QvHYvFOJp/FX+WtEF9ojVHaAoqTSCnNVt8eTdBjiTHNI2jX
CUhWYRPH7VGGQTWwHWavDeTzS6i936vMLnQdk1Z6okpU4855nbBcg5NNCNCnOkI3
9ey4sbHHQ4f06gkSAdSQGbRzOHk+5U4mQXJ/AUF+d7md7rtisi8Zslo9LX2vexZZ
lzZcnA0z/esUHaOSj+xqN12i8vE0YM+4NfJgX2ON/U4plJrjwKZ0OVYT17urZ/KY
1ZzwFXfWBBuY9AlTb+xniHw+YcnqrR92Gt6sSiBwi31pWiO4S9ebhl1HpayTp0uX
V2zlyDJEj5DQqmhMr+En0beIVXpF9vr9pxdPzAmR+ABDwuTzYV1Nee5buMbYKJtG
Z+Nx68Ji/knIpGJzF14sQQzawGfXWaogDPSsWQ1kp+us0zqZGkEZDUIEH7sYD6B/
zKQxwjwvpEdqomdetRwQvtpPfKqSgs7yCXCJl1opFhBXNH1mnhZehx5m3ui+vt+P
ppFXFuSKhqUH8WH/5AjbgtT26clnDuttXqc+M9ni1F32/YYT9Fz14sOmbbZiU6fS
ShV4+cM6XCUFfqk2KB51cIheu+n9VTUP2+ottkHx9lmXezftkyAGDX5pFd5eZbWq
7DkTI8mw55sKVGv4NZONXSXL/YPiOAd7lLvGtcVNQeAEm+Wa+V6HOAd8danGHQRX
5uKZdbcEnjnd2+rSr3OcesZllgVsRjFJ+igUHSrT5BrRhu/ybT5Rm+tHxm6iCEGS
CSVyW7tWizeU64ca1X4jKVZyYxlm6CTS1oBWKhsA4plxTqHQtJA/GDRemdugAj0Q
18qLaG5q/P+xSeT/wn6qy78+Pl149q1kGqDQPFpyInV/ObGiedtjU7tu+XD9aKwg
5SqG96YJVtX69aDNqX7VVi08IXcRC34cG8JByf0KQbVogE0JAsJSLREEP6TbuNYK
hbOWFuUhjwUuQOIoE/XrrFV4Evg2Q4sxK2V/N9aInOxkbs7jvYyNk4h3gMbANIUr
qmKqb98X/hr/IcdcbsJEbkCxpar0rsLU9Pqa0har8SOb/Ikxzb5Qz5RNgPpeQWDx
32VMFCcZzj27ZsI0ZW/+QbOCImiDxBrx2Dhw8FOZODaVIif7ccv50jYPF6eMoXrT
w2Gu0gdjMJA+76BFYI1LGfqzfvKeDqaq0Dd1GciCwoiYgsOD4348EiRC57E5jZp2
xkLPHxWnItcUzZy+LGyjIFrHNR/HAq461XZ3RVEfiw/NJtlkjjqlHGFNMEXJK9NW
dYl0nLfraPXa4QweTracsNjJrbLvSrMn91qf2K1XY5qeimDX9e7YFODRHDnq1ddy
UbLbQdlw+yBF+WcrMNSwknupZWsIe57fhLLTmhZTyS91v9m2SVMbG6J/SP/cOmCk
jhlagoXzzo26pTuOiPcJmsoc0TrVc6jkxR+WYzv/hXm3u721D5VXYQGC0/EOoC0Q
UsbfNwmccFX2eBCpvRFbF2QQWJME2YV5LWUU91ewq7UewWZ8wD//goyjHRF0kwKA
t/FqBMxmzxqAiFN8ly/F3OGZsKwi3PS7ZJFS23aAlpnJtNqV2xXAsjMe4Ye8UvZP
9raN4+xxegSGpm4jjmk+q9VGOCvGkaqz04GR0E84OixaJbFW4TwgXEASV0fdixjX
Xkf6Iv45XdYxL3h+7f12PbvNXJDMpGt6OXKa2xFMFecOXXf8ZiQq6LEBErP6qhxb
TwE90SgQeZPtLj83aTR2qbOzu+wyrzwLQxZqXtruJZQxFjuhycQy5MEv1FjjpOQH
Y04C7LugGMjmcWp+nTP94shVN+34MlfA+MlypHQbSqH+80bdObbtLslexrsKuKTt
vrpdHoNagTsuxfvTHk1DgCq96GCfdLnkNjAEk9MeH7U4x/g6qGsUUhoG2EPwcT6B
AtBPQ/1V8bxocw/q5pC1gVnXvkcqHo9xVmrb1I4NckXtDHStVirvzjnrc557mxYo
PCEeVBJkEIMqaHA9ngC6Hakc0ng4K8NPdhJQkSzTbN+pcYBEjL0Kxs3jhAAdbVAV
QhUN7I9frFmS+BVWdDX38VE7hfxP/s6JJDZGsQ9mEEyxDPJGE7gLIKrMg2dwiWIM
sfBeTus1kV46R56J7iEqlmKOg8iAOqGn/CKIY6bIDb8Hij6DqGw19FUS8nITOE/t
ardbHP+MdauyGKGBh55R9BsBkaUSyLi2XWVIQNcAGByDdfqMIxe6ajJBRJ9e5dDN
fgihz3flT06EHk4R2pJSk7A8eF+we7Hz3UwuePhwN8sRZU7RZfxqTXHrCUTQatxB
LdtUeIsYb5CVDFcf/PyGP2dfblkp30eSDXfOo/8m4lpVzxodXJXhYJ3k05fgQGfe
zi5Nms7be8XvvxLWcFbNvCtaMnU9M7OgNDRT0NqHR+03sbSS6rwOTda9syay/It7
GIjuEF/R5B1qqBV0TMuzhw6NMQNAM5/c779Z2lifc2fPRpyGtzpNIXEy57pwLJ3a
reyiCVUvsdGzbg0jKfjzQh+RNvaJ0sre8rg8Qbzw0WJ1qxsGZy1ppqoitX+5iY4x
AoG9fxEZXECFwirC+Qkfh4WFfh9RBrnbqUYiOkA3lCQrP/RyW/Z3OTRENZewOUzV
PeSgtDV5qQFe7zlwz572XhPMMf5jB5mbkwyJ+7u33F2w8+alfjMJ7UtT3K3ItWM4
UD7H8ZpgzKc9sIbyoXbt0uMRILnlYBhy+zKI++CPAaPpGTqubceUlrxv3760uVKE
TZ9ddZD29umyEZjtpsg8YZ4ldjs9m8N4WmzECbRF1VXVlGNPH9HhoOaCq2lFpp0x
XbdZDqPYQR3c0u279agnjirroAm3mXchQsRnek6CinZKRGfuLZxy7R8ppyGo1bxv
n4hBsMxibYwRmNEGNNpYt2yZffDE+/u4eahufrfQcfRcoKNARDIHHBmoHC30xnQF
yDCEYz+6HjQxMteNzKSRQQD1uubYWnv9lk/tioVi+h0hoOXnSWuFsg+nMDQfw2mG
UkMsz2RbLgNzk1QRi5TWf2mPkiiE1/YeUk7mLaFUUdxVFwHowSsj2r+ji3oKjQsS
O4GXgiVj9prHblis31zfSGvTz1BWmUNwq/qpWC0/Eh6qrcGbhlD7IVmjYKwm8YHi
SRnt2MlIbigvrHFuI1k//oLGs9R2piVmWx2BfhECCuM6IJqDx1A/QEJUCOS1PQEb
yYZMU/JRyWRE9cmOJi0cSCua8lO9g/FmTQQ/O4TdHLajhPpaAh7bt6VTlqs9es9K
8txGb/MROjTxZyhuJj5xMJ++KLIlqSjH72/Wxo5Yec/ErW4hyJJSq86N7octHo5n
doj7uYS/c6mSF9k5ZSgEFXfLd/+y76/EKFU9qTIPMdx2GU0oUSr85Qn6FDE8Anq1
1Hp+wSN4g8mcphSfQofXjmfz/yHHTB4pGqSum0UG9PpvXClleMu1EDVBh7BHF4VR
M1K93P4VRHBQeT5lNa6IniCsVJoeWLrSW+CdOhMA6ozqSbab+jQ6yKiapVplwkDG
Yyh6NN1UbuJjGlf/wZBg/wubcHxxyqW5jkfbFZSf7T2GU/0QvrENmHjvLPAu6+bF
rK13TC9ZihSMqsb56Zx3Qdwtr3p/9503K2ycstXz/UHMk+Ll1Sr4eurey/t6W8kc
qnMFDvs6C+L7NuSPu90gmcKD2kezYN14y6UR1Zv6vGSwpawK+aDYjPcod4LLn4I2
5BJheG8CNURhuMlNLmWIRuf8EBPG59G8ZUyFPHB+c1cmnb+SfrWTTp4fj9xa8qPZ
+RGckl5/153znZlnW/nitEm78K5gyrUqcBgH/U4FAzY9nSyrffuBx/XH77mZxE8I
rb0PcaznQD7EG43BGBmP84Wjul+ZqndjO4xkjx4JwXazbrAjXH8lZJuXzt1HZaHx
7q4lbxFcPUpTXgAZjOZfdh56zlkOuWS+/SMO46XyeBvF3aC+yOuyybcza8g0W0N7
LLl0GWvZSTbK68db9XlYKynrdxsmLDw2g4zfil1Yz3PhanLGmSa+jdrY6IT/s5Ey
+eMjnQfSUwuwGOsEA6skTCSbR+Umtpgq/fXmdeXYnEpwXuY3fQvvP6qKw64F9rFQ
dhxnXrwDYoO12G4Rtt4Torca9Cf1g5dunHQmKNw/57Q/Vp/5vxRi8N5FpiaM/LCd
3jQGWSoaSlcrOyCOBAS2Gq4L1//APUKrwROE/3r35UgghxfyXnz2/NoplqsHq3qf
rmJx/bv7YjkY432PGMZJ1YojWnY23y/4fdxHbizxrZN9Vkdja0gDE+ATnCeAMkMJ
382rv3VojZDzdMwKTic9imI5jWN6f07te5yCpBozD56jpjyyoUuCQ+6h0w3sbIx2
5Jzv4Gmy4AZHfDr36f+S5JoP1MkPO6XWYYFI6qOcNFMss4RGuobTCn+sohu4hOBX
0LTlD0HOtUf7Hwl0iAWXRx8Z1kbHyM6ZuD8wHpECbME7wNwItQtlQa4NdRQp9E9q
BE/xpPJDqQHI+QtKnaXHLhwT8MELQofNTG3Hn74mJEyzy9Q0UTsKjzYaqnoe7u0i
TukrxUv75mEVGx2uc2c2iYJkeMAj3vJfps1lFkPsv3LFJWes5QMscLlNWMjxugDs
Ssiblpp/1YAC2NIs7YT1FA2EMxWyku9xlp5ZKkTXd/0QIC6UMqBtdD16V38X4doJ
7kBABIsx3Rqcz8F6eFLnw4QGPT0e9xgK8ckiNgjxZt/8aIydO2lX5UrkCXRIj4LP
2gwBh6bdprsuHqdZkwVgMs0JRosuAL5pVWzOYJCccx00JFXwpSvKdhZpoWpixz2y
VgBmzqJqdfcOdXmX6/ozJGzftHAHx6KFWldavWNvDDi7Siwvrs2QfvsH///i/Iro
NAA0L5nNE84GLxmtH7BXtIR0ddiPQWazont56OsDqWAe0ilBKZBeCrFUEwzgDxaO
cbb5bZ59AntgSgIZyrDSxi+FLKol1JoHrlY/nR4TGspd4V9NOrl2xyQiuw62Fh70
xLolLjTLMWzOi/R5gf9Efwl1UC8q3NEPgDoWy+jrdU9A3PF5UTzGdGIjQdTZNEOG
NXzx8ijAN0Ce+6TkIRbt6malqqVIBmYx/T/biv25MbEXuQc5sKyJlNOy2b0d4vS9
CiGT+3Dn4gUsj5wDHA1FyW6MoMSlm2VoMxje2Pif4xWdjR86Ip8pU4jODhypkaq5
mzkE9z85PhniflL0tunwNcDE+eFLZFq6Z8krloU9KD5YijvYF4VrgA9qMP9iMcgV
jgZeQovO8RoYQPeiTW7N7pVM5WLvnQplnyaTpHqYcvcaJuZz6BOlxh3ZJQaJCxCr
dFNOctcs2BOFupQy+WQV2fsXCFqX+b7qBWp1PUbSJnMQRPlISEa2lfpcQ4ihrzSJ
f5sUIJ2itQQTHYSw2qHssxA6SoPGUhyzhKMNDerJATAEmIAT9rzSaKKxDFsn5dhs
+e2+yNZopfQRGPdlfTAPOPHRQLeuDK7vkHdJG6iGsRvUryjtI39ers6XLBJu19FH
gZJQQfKrpS9OZoFV2JvKq/5PTCo6O2JIAJCvJScOuiUCVZdozNlTwkZhuIirk5b7
DcZOPSs0oaIZ4S0f4PEiJDBeaMK8JrYt7mhFs18ITl3dOCf4hJQnpKlgctDZayNH
CFL9YABC/opipTgGWGGpOv6KVs+wHi1OZF8khIvEcZc43E/Kd3iV5q30UVXZ7nui
5G7V6xySb5TT4ZgIaYW2NAjB6eRilOIFPT8VbgmNUrP+GAHF+Ojt9fYM0xM8ypU+
uE+c7uVByNGYJL6RNzWhgeg4FIWqQPZhZ8lIF58d94bHyHuRPhiWLxTRkMBH/guC
iurm6jrP8eIBou27tdC8NwmpIyJ+R5IBIHYii0yrJkDPBwNhzGuxSDZjVEfNr3Sf
dNG2x7uixLFakX/ZagavTvymXAJbzj0uxaTXspQ48pB+M+JKRE+nVHuqOO+GENsH
buiw1GmSilHV0ivq/X6WywfoX3t8kS5mSf9PF9qzmovibMpqLPotZNoxhO/ttF0g
6q9dtWKvMp7QyMYKNyUKj5KMmuvzReqkph6cGOQdNlmgRNAPPM6fp+P6lbOVrKt8
s0eSNcYE75lVuY7O+39JDFk6mr31L3p8DcRLIF2v4G8K2rfjlInLwdfx9OXDVUnZ
ABVL6ZiT5q5ERH5/XyJlCIqIj8jasQPYKkyMnQhPevguGR9Qxf3T/u0pkz5JApFN
UrchSUw8ju3Pew5OuUK+iK7f1hWJs22eosmjWeEIYWTaeHf8/LRvye7Wh/bs8Q0f
qL8wLQGfDjeTNEiafe3oKRegQsoydMKdEWkF33XcJBP8oqpdlAzxZyAcD7tnuqv6
X42QPLMeOOV36G/ACa/BNnsLo0GuDjKY1lz7/sTaPzj0hrm5bj+3g3p09oWmoPFY
truU74llo5K94y2DsewDAIyQRAU+TIDXR9rxRah1xmAsrKz2HSW9oOu5QH+w9AQC
+kWnpzULncq6RyiIZtM1Wa89jtPs+bdKP0KIDitGaA20bfSgpa0WsAW4FUd9EWg1
74wfmXnnphT6gUXY8qnGi1kKpiqthdzZM9Rd5d2UExyMcVtgD00Coaxdwvgvisau
qCR5HqOugUAHi1ixehX3hW2VSNNxnaKJDyTNZGMGiAk5pC5fQ98mi9rik1mApixI
mgFYHdCHhWzg2AlJ9XBT6zqE2DaHknBKHzFkIz1T67XDcTzcKN/edwtsfjHS3z5i
abKW7vLPSa5F+lwP+BNKXlbbVbjsDuy6EeNs1asnWKNehMD1Yh0vg/aXbRTqUtq+
4Iqtoa5jseL+3bX5R/JBoSCKe4V+RL5UJqsskw+CJpX67spabMgwvfKuGfkkuqgU
qYFt8Lb3EdtwWh1M4ulRR8M9JobBrD9Cks6KVbbr4NVgrWKbhpxhIkNRL3h13tRB
Q1lW66TNAQyAak7YTKrD51YQaBim6dbWfXSbQ5RflVYO0eCEjkH7FW1u3JnnRLxk
4EXdEWN2ts8NOktLnWj6XYRWptWyL0+Rt+EJrTG82D5y231KJxLDI9sS/9JojoN9
QZORxTWKk5dlZfi1TXDbOeB6BAqFNd5oGV0DTVBiP2nNe4QZm963hnC9GcCuqjeh
thfUUX6yXFfQY9LjZBI4m6WZXuxAobFajJkhBYHOxA1YWEp21QNy1VO1B2CEbA6j
iMC2bAZs/eN85kj7ROWRZGa353oipgEsTafhcg8dcfs3CMcbuLcvbFm7usaiJvOE
LVvCE2GEd3X/SKFSj8Z4hMQge0Xk32xbPmR4yzksgVAN/XiZdpMv8wQ1ywKngFIo
slhbC5BXRmiAMBB3MtwuAzSdKU7XbwXmPkYLtS5UEYjZIjrYftFAEYUQDCrq4iQH
hGrJzjA1BFMCvoMSfkPzHUugz22JO12NPxsprZJL5kCer1M0GZet5NR1dsqHc5Xs
wY4Wu2K5408Yyo4Spf5mZ2qgBWjPI1Cn+PLqDYjAWdQqMZUwuyp7cFRloMj/b5xK
aKTN5/5+o4G/ur9tRC4Vk0VNJp7N/eCcqMGp9gij5FdTRnhk+5lI56O5WyFeE0+0
/oaTwz0UfmseZwDksfh7yq7Gr8BZe13H4UCGpaCsEE6Ji2MKJsoBsL4sfMVgdrND
8pFElv1DZSYx9vH4st38QdBZqStqTOL+rE5gT5xHkSRVDHgOvCjBBzLrh8nbpzJB
cMiYnAvaOOIDwNEjkFGFP9mSrL0D9LVYPjADvIyBsdcHtL5Rk6mWIWAwBB/gZiJb
KgkGsO3FEVniqtNLAmBCS0Af/Jo0B+30+YqZnj+sPmHAEd+KDek4j9UI/9gqNWc0
XHStCNAzu1DN3/Zut1fITpnM9h0udw4Cee0sJQ5e1/b8uFJionaILvTTIv6H/6P7
CuZn5wjKj06dSljzecKdp9kdtwlw6CmgNxO1v4CUQpRR8j3qG/4/unZXofl35fPr
5jx1E/Rl8PQdUMl7aBMdDtIcPJTwLPv62K7GjiIQwsC+OcENDmXIAkcQjW8K4LR5
oHMW4JYxKQYfeux4cRT2gW9Zh9ZLFl4NjlJsUtCRytcvHHwr+YOGf7sYDavuvoVS
MUpgZ05i12ccHACfMKqJ0wRCWQUuiink2opfP6FSqOCn6YVZcBOXuwMPGLH4GSxu
rPP64/LNvK5owRJD1zRQnXxED3loNwAW04Ls0OhbfgkGeddJ9AuR4IpbC8isjCx+
m1+8xlu1o95g02VXOmFtYyyx0asm7lXVbpz0qcfmS0r5KO63Eyx2XzG7t63KP7LP
RFiP2QVXIX/vpGYBs8oFMPTmp3m702BNdePYc/CuQY5JVt4oXGZKylY6yYgn901v
dhkL6Z7o2H/aZOOQKE/cj8Wb+pjxF805mAslzU0z0sLmvC7IggdKASk6KokBzk2J
iwUM9HMjODm6Jwfgr3D+HJO9LuuKnTv4QlQYQwKdEHtEI/lb8yzHvcBqFpsnYOMo
woy+FAJVHl+zMqzPolG5X/bJxOR2FYOp1yPGKC/Y/6aa7vsWxX4m1D2hw0ApHEqB
9cYMi8RXuIZqwZgg9LkWQq6ZKx8D8pLQSOFL5Izve1a4rKCxn2E4C3/WO+RyRlvQ
2v81g3I1RcyoUfhz3Pg3op6+p2njFzsbrKvB2qqEO5JsqXdwXJdDFwuUfNSFwMYQ
QuUQQRlw4kEzHrOBjQViuvdATHzaKu/gP/PwrOtpLoFJN87heZcPU7ij8oG9RNLl
lgcTR1okqxFTt4kXnuIDFZ9akzw48UaSOTETVLkLzbLR68adgTdL3lqDH+yMfP3b
J8gvCfEmnfL4Qsn3+AakxXzN0rzVqAAl/dS28fX/P98PXw5ZVB3QmpBdHp9SajR6
JPMNICFMf6g1RLF/HquaMSinAvwX+di/Eru+GNzIKBqozyjXikrojZw3RrHd7E6t
z6KWdH/eCLigRAhAw0qkEq6uzwbCcrSbssLEooO6BVbXdwULvL56EBjEvfmNlx20
OEnBRksLL6jwg1XKYi0WVY0i5IRmu8ptBmXK16AGC6MfHkpsfL6REoNZJkg0Zn6V
6IUvRKCjbtiQkggjZ0g2Q4iITEnxxOt8j+9dA+B78wxBxzK8IiQK5MCfN93erKWl
9nJveLrlWGGmLScV/XtM+BprfVSuvTemXM7XXppoPUm0lc+f9XdNUXL45ZvU0X+1
l8P+kIoysODTdK3O3t6UTnbzs8ZLbgSCgrUq8XzhjMDEOWmDozsfDaYAza7UU/op
7TGE72bq/3B6zeTGrLbIPLbGLvAoy/VvNAOcNCQbz1jYYKYBAgZ2Ifg5A4e/fE/J
olzKdb7NO/0jL1Qrk+6JOTU7DJhwPBceLjAr4r+PVzARE0HPTQsX3wZfPRn4Sq2M
P8qyBdjkkO1XTqtbNTbHVr1Pc+OT+PKI1UTS9UUZVoyE43FFxRmy2QfeEKaBhIwI
UZMt+SY6grsNjlX6ZgJ8aLSFpmOOmCLmRCuW2ROo5npJWP6AV5BwPrbBHb9Yg8i4
Xs3MTJmx3z3zWBIcizQ+7w2MGsYTToyZY/cP+iexP5hbUjkm/xK9Z80c4ZTfnzub
wBdAzBIBC4Na+OLs4r+e+NiP3k1Ik2DMuKIMnJaVtTrnrJ9Y5uQo5vSGvhGYXHE2
a9Rqni0GKxTdlA7F4jIgE1AjNRU82Hk36oVb7no5Aoo5Hkz2Nn2elxySLEIj0iTO
j3UXqzLOB5O4lmyFH5bFaD4bKwhSD7AiFC/r4UiX5uvBKfH+SOSNaZ0VasmEr/5p
ipqqQn3yoqfwiGjkC3nRxFDaTsbUalcR8lekoi3YtxqecPcOFijZJXBWuaoBHQMa
k3pzMEcvKiPLu7MoPf/KXN0FFmB0VgXrCgt9LPJon5rnZ6B/2xY2FAR62L3quE4P
cscBH3QCLmlwqegTfjnWHLc2ukCzcGvmxNCDT/32j1ZP7cana3bEpGF8b0yf3aEO
zcJGHqRoz6dCwR8O7aj8wFnRZiTl1QxNfDGQPol5WpEwLgdOaWt+Mo/a7qqiZaUb
UgBixbpw0R6LXeYOubsslZQDvRKDx0EWH9XFl1dKhLZIp6mlBR9AqC+RPuwv4ApH
TPuQbCUMR8FBP7CbQeeiKMSjfVqXkFrKGGELJ8vt6DljTOWOvwXlQu6PO3BcCEKt
QZNqsdGwmqYoY27CHKRk8w5HYzZK6DsUNrh1GS1kg4rh7WqhwwqzWUkYXBj4z4Db
yeRmRVerEU0bUGLkMWckVBhmQC9/AZGypLK1tDPBzvsZfrBUoIPqQ6QgvTucJ91Z
p4yEUUVsP1OzoU0xwwoxbFKiGWFIgy3wmRIY+jlP2CNYC0ENxUn2z+AJHTvCofIo
7eZ10+G9NtP6u08ITaTrkU62DPh6lSeUxgFXlrXMD/OuSUYvTAL1pEiDvfD32DTI
5aHywFs3FwqScT4duI1Cqe+sIEEAsxJSEoa/7Kr5RC4Ktn4pQ1BNtIgX5aHfSkLX
WUImyw/bWs1LSJlIqWhpoQEGaB5MrrAijF4bhMnnksa47ywNV78w2AgUwekKeA+S
tq4gnRo5wTaCoFrCUcppZg1YAhfLUst8NpATXZi3U8il5u+Bx/1uI7VZKQO0WQVr
atHQMZe+rVXlyWKpHbeaDR1CXO58XIj+DTRTasgCnZMWhGzQRTJKa0e1Cb40RyMf
jxLQyhADqEXSH9w2JEx/nNPTpExJGq30OuksGCUUzi8TsfIeyJLT+lpGNT9QrI++
yp++EACMJUy7fOt2eUoL5J+y4oRdoh+D00/jfh3601CSjNtnXPUfFltB9yYCCZKS
pLIaifazxp90XzKNU0YgmLcy50umi6G+ClWCkJpXW5F31MUrzDSDiXLDZjB2FZsF
ST7rbjRu6RYZWxH2TsdJTFRROr8ygGpCxy93GY4GIndLK4A4a6gEDAjuajsklE2l
N3A0zXDanvgnA0YqXoe3BPDfJgy73oztKkxCQlXDf1+gWrKPfvugjV8B9/iPL4RG
EsD7Bc7Y7OsCdjttSRu4nY6qnbHNgx1eX1J/l2GP/Rge02M1SNCn/xeZ9LoVU7mV
Y317yW9B0YxYtvFVRKz7ekqlbd08f0ufx86cSqz7DSKbKlSWmvuovKqDR6FFKTIx
rK/f1LkL6IEmzHk887ELC1iznDSCbGHBDzt2vE+RL/t16CMOenSys5t1h6Ba3zkE
XuxFthiPkxw9ZiBCf0zbHtrTqZUP6lypzrF7i/zL/5e90OLlBNPC4eSS4xHXsutC
4smTeAEFzrOW+jy2Q/Qqofw/MGN23IHPE1EuLDSod8t4BSGbfmLBsJeRDf9y6rRz
AlMaH0i6aMqSlpKw7eVIc7d7Ncuvxjxh/7nEyTkTmDl1zCB+x2OzJaZbQkTL4n+G
H4aM7wQhbZ9uDKyIFsPianYGr2eWHvhKyH5UZ1byhFp4+yfFfed08wcurZrH/MA9
+avW8BDNstmYD1IRbyV4mhIUbI+kRQJQ4hu5b7GwtiRXy7H6ph7hquxVer1kV3Dt
2eU3mqbbHpTHf/M2c0eHNoqOzNhw7ik5B+v7dGfgKV96mmHBvYYXCsyz1BCpMzgp
Kv+1KCULITofVPbZ+fWTUH4gsr+DBLtI5yLDbzoKBYD01d/sW+lnu6xyLZ7PejOJ
wFgtJGKM7wTTs/GIBWgkntw7lNxaioXxKvOXfouMaYYjox/1e8W8hHfRuBGUSUsR
c2BQt2v3Egzi2xBft4TyIN8aP+yKo60DWQxRFaREfvKAqUxRL5dmjtrXHaikzL0E
HBvFR97m3t+HArCE2RP2YQdrz2U2f9Gu1JXM1Ce7hJmXQkjiwae5PKQNrmL55gzR
e1jmVWpuH/A0KTNcazhUx1NdV0ZUikUFs7mqs1CZpp/H36ttf9h2TKnM8waNkfqs
x90t28Y/6mzgDRFlY/h7OsuzATjyMc06XUxQlFMyAZVYbLXvq2IslAj0qPGva/oo
Aqe1jLeBq49WOLXHGcu3mZpoHO7EHqeqnq+EQGV7H+t7PBmSmxqzqa6PDdB6PMOG
+S5EPcj/1RJzVz6h9YT0Ph9EYpSgyQNkkCi/l9w2ODgAtmSMKv2z1iRVXOLKG/iO
wYpXsLi34tmpa4sHzPKQsNwPxW5WeM//OgbhW4uk11yVVsBFfSErViHQsjArz5Gb
KrOxooGZHYH0psRpvKj34lX/MBRGuTin/E2hgC5mZ6QCEWVMV0H8t5829g31oP1g
S56jlZX4tKQifi6Xhbw4rZL33JmFO9L26DzwfAaoYcoJaC/W9hfOwEKb4z1aNMv/
dy2cecAf7L2XFRQFdigysvdHVpXfcwflkDV0MBMkEwHnjUI3xsCtl6oDgzw8NEyD
UR7s7Z+d+UsIlHSLF2qYcssEq7eMXfDPr598adtGWQXV5hc7v7jU8053lhL99iHi
F0+174UPmll6NJADQAnGFJUAWuJBBk1hf5Ctt9sH30gmYpABJq/1G3TmzizQ2ADm
wn/a/VKaPNr6cCepe4gVG24dtUTFS9pBfLOXqIfvAFusAWD8rY3F+M3SjbX7FJu1
kaYiz9f12ItK3q9LcJJQzo/vk7eVrkbCfxa2w1V91OZekYhLqFwCoinz09gM72vm
Ccz3b9M4ihq1fjMrhyxO6i5xynJQFC2sMjMgm7zkJTblr07nkCjIZoKyR8NWdZrF
cR730kMn1F8pHWGhICaY5OVyku3pszMOPLRBBjwmLP5on646SndTQtUiG0x4M4b3
kV4qaQuh0KpOMdR1yn9ZhOOn7OYnbveY5WRyTlagsMBN7KYwCghRbz3fg12aDgNN
FEp+nvsyByCqFoX55sdQn1tpnKPlmj1JgdHLimOr6gOJEjZ0Ugkv/9YAKeEDcJVx
SLlHYIy30mjpYkulqJ74HYFz4Cx/ELxkyPrt6RDozGCxD1JU2Mm8clxxDRvK5RCT
p4MttcTOKtZ/+19byd8vQOyNk72ks6QkKNilenI7ZlBYBIOLg+CKGSeSfuZ8yrD9
BP3n0eBY89brPQguJVjMYqkJ6AXLt5pfmTa8REQr9rGT+SoPmOhkOkRSrjvRBf4a
HdTzrhj7O6KAujK+H3dY9QzYvmOLUynJqY5N345pigTJO55Do8EV9tfU2NAwegZ8
nDBnwePUMXkbBsnEb/WaQ5kxjmjd81L7QkMPfuY2M3BoXjQcA9hQlddXWuV0SY7j
4zt0Dy3EklLEWGXxMbuEFfCCRRsrwV1kdl313FzzcOqjt6Fr3B0qNYi2o1kjLoy6
TZsIptiNHwThwFe0WuQcgspn2GcrH5JPzmy2xoGCUjhVzWcysyz2QZgMpTvHq5kZ
J85jToWDRW90uYk0REkBYvQfUS0/kRQ+8NQd+uF58YrvUpzAfc5xFjwSXmVHs1Ew
ZQ8mNLJlVBMANmO2M18TWS855zjBOxiilki1nqKk13PaBV8PEcuEKBM7dYL5gnNm
LXvJ3b4NIaRJ0NZTQpcWsQzfsKC+vHdR2u8Nk2DAOGykIRURAI2Gdh9pQx9hBRBu
5gn9qur6vx8y5Lb1l42f/tFn0qp62NSsXXOiv0uCD8ZLM7mVi89sdav63LD/uRzb
5e4SbwX0kglxdzEmhx9XZ1AQnxio+iMB4MUQFZpnyGeoznMpYWFau7jNUdmh+6J1
nkrXsJ2FYIOE/1q/wbgx2YaCYEobLYHdaaM5vCdO9rZUdtzxO3kRH2y69EDIlQ6L
jC22WQVVvKmZukFDkTuSza2ayQxvyFxF1+nIHQ2dR4kXVKVJB+P67ZWNVkceOaeK
igVB/bz8RMdz13KanMJfVYQczhX5eX5r33+cAJ3cz82m2qQNfrlPlbX093ekz1NZ
jIIyUQ7X7eIrwglpWcpENtvOXbSMijkrvQrq8YpOR1DH1cTREUH/xM6PfURJvX4B
OqCWlfXzlK5f9mnErSDbgGdbaJVJfXLklpIlZ4fI5iF6y4P+D/uhlBMVY/7ZMxZP
RywHS80ApvR/DDPBstlTVKyvkEXiXgBekFmEYbCK6XFSXpbQobO1ZQL+TMjYCC38
wEZylLJeKbZgdh/+xPWvgc3V1avLoP/nOiR4GoeTomxGLcIrZwwjWZBLJSGfXvr4
BfpAzJIG2O/GxwnldzgBHW48NBNxExDc5M83xv7zX4BW/+QNSPm42v9fYd0Ki4zL
MY2q/A5r+m1804NVigBtNQONEQl8XD8ltfrUrkrKpdizsrdbg+y5IvYRnCWgTp67
I9/3dx2TY3L9X1pH9bebUaqA1qP2hNO2QW/pr2HITf0Tua6qzmMW90Kh+LbYeKk0
XdqX2lBXgq5vVQAr/2LIOKSzhDikc0Si7wM3Q6v44EIg1XyVzZztj/tJI8D+rRAE
cZFfL5H+rrpZg2TsMA75bAI23Xkf/EHOrZOSoWTYjjheuDGZeyyH8XUMy6shZ0wA
ORi5QctFZrqeWXlJK9X2wq3gUPCFeMOZOjZIVWi30jG4vmhZamVwjIcV0F90DN4z
3TUKG7G/rCUUvWy0r28Yn7gGgfPf6AzTlVmIzsXbnCSd0jGGJyWnOdQr1+ascXVN
pXHTHiKAMjsNEL14Ap8zdZ547elR/E/lHbKoxeCB/RGdz3DAfzrynIsyAJ/YyEiq
+Yzu9m9ETAelRcS3xnEYio6u4mxNwYtIo8RvcBQNNmm86O6M/71EIUokEIX1+S9G
KK2jluHGcZlpzkso+E/u5NkuQPCySiV6R3M4AfTQH4CadzX5yZ5eBHGhUN6QoevX
mp8In79wmHvu/1oeAmXpQasnVELCatvZSeJz+sKyiRjsC28cuXpH7xyrJHCtNQY5
cvWRrGExh5STYIuHZ+KDNoOF2vF3S7UInxh9ocm33Nm5H4w7YScOVGw39Pm7ZWj8
P73yDCBhuSuaNgyuNJjA0eQzloHbq12zbL6LZ1fOZNYMCLad7iEt4B7LSzcy2KtK
JlLa5eNiZltARj68UcFtVAjswX4QvgKmTodq4wzgggWadqL06Q5dNBTZWxJCHHHS
gU1nHkeEkll6NV6hIhST34ZynA7JAJirkGCwcbtjZTkQUbesqSIdYRl9CduVK+CW
/jBdnLMxTOszI0J2Tsnain7SgAKS+XwYIYS4O6ppH0EFYq9M5SLv65z2QxEj4JOZ
pM97sqC4x8YGSuDbujyLqbokPjgob0ZdVTPP4pfhaEt+bhdz7wVYWYZEqPlrcpj2
Mgwx5ESqW8vkJddIMnTGbs6K0cNz/mYrHXRrYOPxu+HwGZghXQHLOHJl3wORs6fa
UCWnZpB6+sVMNJZvOPdDb82wgBVACBIqJmsvBKg82M/3lnWIhAyCuXl0HZJ0q57d
JRqW3+VuEvSKq9nalPTUn2BL5zSucXhKOneeRh18WbylT96tshhIYreTGMg2aX2m
0ap1fKrGQu2xyHoRaqT/zREpoNWmzSQ4yv2p8Qpcb82rlsK6HIxt1SsipLul5hrE
AY23rczzfSO2U1J8CJL6RPZudsBZ8izimMja0aO4+ba4IGsORz/NdD196B8JZx6q
C10S0Mpmtt9klOFQzsec/5wEPlO6oQbbnAzkFXQAYH7DY6DNFz2sf2bgI4wzfCGA
UVnlCHOXCpm4iLkEKaPD7j2P6PhaeC78dxfafDrWLZlc4T8GNp2BjWgtAjx7XlzV
firMLxaNah2BEzHuWCeFsscpw4Dwq+4XlQ+ogB+a/vIg0OTM5K0dJk5FhKqeKd1l
xHa3xQNqzkmjBnmmscRLbGW8UfRRgLJAxq7z8D0E5/fSXECviwEZGnkPLuOmfPRq
H7Rln7xlaHkyy+ZpD7+XaAXJvRPe7vaGlGk1AjM0JLkRldWE+8JWdU4wneRT5k/4
1Tc/ZYLwBD9LIG0foRE0YnmdIZF6Kkn4pjpt1EubGP13jv1AGKMUQ8eKuZq1LgPb
vXbFDrqfAXwsMdhd+4PtcIKpyvzwFYal3Jy6gDRQjMpcUR83ceKcYvxSzWIOsmVl
3JfsVHeWzn991tzEmYy+SfagNquCDzA5zogyO8H4zP2HVyyPLohVu5erhGA60F04
4wAthW93gcOdDG3hUNNe7HNlsslHlXzIq7EdgvcZbp79woPeVIMxpL6XTEoeeX6e
dVFcBoqErgWKvYWy/1YliXw/5ZZYuFR32LPsccNGFDs3W+Kp5rqyE8Ahz/pYouJf
Cp5+M41aOAfGzdyACa+iFEDatNCbv7Wcvd8y6JD4omcsFWCdXTnnEGdjhHUt5WFw
MIfAmjbfWFxOs9c3+wXrUK1GRyFjuePpKiLfsUSHrVpfpIPT5dIfYn6SCOx9U4+n
XxCZREMcZspTgZajgFrvl48kND6Z5BDVhNqpi7AP3LyK4YBK/mHKrSUKGor+jFAZ
VKqU2aHUaM4cAqI/jlCr2Haj2++VT0p+IDZ1WCkmEyEF2kRXV5IXbeJ7/CnSNu5a
tRJBOQXq1gOeyXub9SncyreoXFChE4nDiVUduDJQkvq/PtKnHML7RnvnfJBNcl4o
iR6NawwDQ5f/qm8crvM1GgRapU/mijDLKaDW+QeAWjaYm0XyFLyRStD8GjDEGSCA
GhELa53LEEztVJ/xG2Ur/OF194isZMs9SBz/NsovB0FlfwOTnQmZndUO8I1Ma9u2
P7CDs0mdj3ay2cIOOYCrbGrrbN7VuXG7o7TocvLphYCtaSSo+K0SfEghh7zpqXXn
xD/c58QX1+Qo58cOPZHnqIK7628ddEaXHTa/56Fo5XSS38sRINs9po7ygtQf4/eq
jRWWlkwaEvjyfG17cH44ieEN6MWNhHPsq9wGCSVLGPS6hJ02gHQpPPm/k6u06VVk
3ZIg8ZlRmk0YhPcQDNilw+IVkGttKenP7752VwfLUSqxbS9+MxpubtRs2Xiz2b91
dKPkUEfUVj3LZ+VFk12MWgmN+0gy6/l02E711bq9y73Fps/vb5sEZBbW1RSmcf12
1yNI4GWN9jSRPSMX2hBaXOJPKU3vyjaV5YAemhz40pz7PZlRIYTL0neMk56nLKyD
cLzX9A9ycdLbDtvOIPDjmMfmz7ehLVlx0b8T3xMygEV0Lcv8D9toTJAflUNEHwtX
bNEhsYW5t51DKY9M1ijOq+90YIEXQ0xAu12e19wAXPJ3k9PqvNFFeIKJXtDYQHQG
JFJYmmurIiv+5ZuSTDRn9Qn0P/SjpQ9d2/oyS45SoMVUbta7oAbnzkqf+fhXlxkr
YLwkkGvcHxMWO1OmJk3KUH96ek6EJwHysZ5vCE1r4qIljeQyhtg9ypmoV4nCJci3
GMtSxA6heV+w5cfW7NrS0UBG6K/bUM9MmaU9IP36WoI0VIQBaJC2r16Y1LmuIh87
ZNpgRelNsfUAdmOkzAXaj4Q7fDkdEkM13GBY0WJiKZ4ig5K22dwr0rcu+g6eQxCO
TRGqzbvqso63YpQItOYE1TcJ9/80d8S1OsZfTk5zPzjeU2IgA2Ae+oVUh3MWRaUV
Ryvfy4jbrFJu3YfevESaWQUWcJ99wT+5RltzdaDjUeHl5Lgp0R97bFCYQKYTdj1k
Ib5Ywr/D8Ua04V8SyIUvv2WnjKzKMFm3jd+dEj/LgyHJq0G6adplt6hewJsOOCkT
NSNsElXJQjZw114NN/8zP/T+UCtgWabd36Icg9qet6er0YG4DtBMUzrEiE9YvTWR
0OmNbQlCaDqWCd1MePPDFm7Ywju5QIyNlObybjOZj8bZx5eSoQa2yWfBp7z4GUFZ
eoCWElg8smeuP4EB+BEXx8P/Id1kW5F9BBRLTf1rcgfeXNCheaNTRBaWBJcw4IsZ
qv3I/X3urNTOm/InfjwVRZJccp3KxVxPWYMuXDII3jMnAv97BVcneRt+8tepeOFL
1z9sg4yg11+af9veENcWYZym257w+J8pTetFfUJGDZy9I8hW8mgfZSrQCL9XA8cy
rNCIQmFHMi74gFl7xprqEBB0G1wipjGgeQVTJXXQjAJITNELFbJaOaIT6Zh/blKU
xfys2g4FfUzKL3mf7PTejRmrWldra4AyqavNSOhLJDefN2VZy+sybd1GulrNM3M2
k2TR5Koj7ysb764CZRvkIDdgtF54EVbpZIg1QrzFZtneC0Ek9BvDoGB2Ly/CEeY/
Z35OV6Q4ssMW1qSDDCi0b04slWX0c8cCetuW12i0AuZtHCSSLRfoVs3KnoDIidx9
PJcUxVxFLl5YTy4PjiEUlnvhVvN2H+sEm+jr4fWkC3z1yzWQm5JmqnrdgNJFNmky
SZBZfgmmOfSICFQHXCLKnwqrkCTFMURaQyHtw/gPFs0FhWrMOvPCykl+dVw2SaVM
EOSLYWk8hnbCr3zIriiHwdi2LjWaoWN+sC3VRWWday8nYTeRxOncKWaeSB3OpiSM
ygXiF9THCd7q87g2yUsDvcmFbvh3npSW9MrqAP36ksQxFZIttb13kpZktgUvy2sw
WhnKChD9TmiDD8mZAPOe96ry59ncLtetOsr7y4VnBVXpSRkEoa3REkACW6czgfD0
fAg4hYq6uGZxnN+cD02KALNgj5qjNo0d/XZsB764EDjFGyPOG9TJ7JGKPC34MQ73
UF/XX0Qaz8Spimv+2imEUmOvCSFcfS+Sj5e/hX4TRJzZC3plbxAhT9UNL0VsJeBr
FDfZydZmfwVwO8bIZ5is13LPZIBMlCA88wXbc+jWjkLJdwDRielCu2hZ+SBR7MD1
zHOo+3m5EMxmKoNT/rERsCCFFd3NrYHgX85/s7Gu8LtEKlf5cJq0dpFNz8ENGByU
Ji0uiEV+LjEX8y2ck8fBtUcO9g0p24PrELh37BKccuEEQBpl8XhYaVCoaGF+K7c4
zsRADyusZ84nhQqN58Qami2ijddDNaenEeD69X4xktCxeO3g42Lc6+lAOiJOpWMC
NGx2dedsjyHCTD/fZPb+5/LUdp3oJWXO2BAUBueY9/q/BfXMg46nQEV0Q6S4czDL
lnIiLOPmbCNL6oARRck0sAGXZl1YrhmD6Xttcjk1kWckHcCdhLRs2Y/kgOh7FUqb
Bu7341f50YQVPw2nG6K/IBSfnAE0rqjgDW9jNOsH5XekvpV4fuVVr4nKU30uYrrV
vm9PvMp9/lX8570C4hHZpzfmdiQQ+TJChVlkAuj1MfT9Gd7xLsJtg+WSbpy04ypx
VwrwtM+nwv0NFUiYq1V0eiRAkILw/vKDnI7Lot7GLmxYQ9DfB6V0B4XvOvpEe4Tf
5K5vFzNTPm7EkrAUfwZn3H20CjvgMINp2/TGXOCpjqgmr26O+6JmG1ttia6kGcbm
zpKJDQ3J/+fK8u+MtM0rr91oHq4gH2c2q3QZj6CTcMEOA/4prYVJbnvi7H+ZD9T2
TLY9tqjcbg87qa/T+NWTEKXGd2YgumFWTx91u9/kjpXIHu1G16yTcjvPddwwI0iE
OPhCJUGq0yTqIClJzJmnqZQGREMNgriXKritZIeU94Iy1pY7EV8cFJmj5AeCn4c5
m/FGay/WOnvP4AilJYLD9gASpR8pIQLPVyN8+y8PeLnYhXxBapnJLAmX6+VKrZ7N
ow0vLW84V2UQLGsJr/aTgLUYxqAPGu02qoVbPN6uvreN90dOAYnNv3vE12/1Tjjf
4ptWe9iiCscp9gaQVL8VphnNTVNu0qcmXq0tv8KMlXvn/UDEANW48dohMrE4q/em
k2/39Yufqv8hwkFXaxy+cU2PT2RRtixcJOpMSfE/+yrs9XPq7gmirOUHraeQBuQ0
30+9DwXq7gExmz37XG99HOjEYA9QsoRE1KqoxBZpmx1HguJOPv9pFmSIuZB+RLEM
MBYWsQRGX5UrTPhtVBBaT+0krnFa+gD00Num0Q9e68DuEDJ16lxvElYtvguz+HML
NPbB8wZA9FngDGVvLwcay6a86iW+YHZEIeCJLfr4LHH9+XD4yGDvx77ciARXYIUu
TUgOInz0gA6FEPxlxcCmHL70vWevWuc4IQsZwme81zi3FGA1If9l2oC+4pnzAYUS
KtuQg/leGruntWsHAIFEx+sunUkZciT7SmeX9fajicHxO6QcJx/dICzE3Yatj9gE
o9DLzmSijLsyrQaNVdKVmSuSOzKu/SZRFUICJQYqJISvLf+zZlN0KaYJkxrRcNCQ
0h4UTL0FX/pNuyzO0d+gS9ayiQ3341XcVaHK90IlrIZO9oHCMH5NCDI5qituaMZa
8AV/AWoCj0aByRSGPZCVaweDnI5MI3EiWEhIqFvbA6990i7iWIoyGtrVjULEXXxG
nq9Ep0J2qowyUF5hTV1u0+0HrYyWF5Icp3EHPgDxVQyhjhY7G888Oq8KSoW4NGIp
E7MAbFTL3tsK9knT1UNo/mpwOPyPQnl7ImopgEIH1nJaOEyWGD3W7hDGmmTA7jca
eg0UQgaWIiBW70GLtExz3iepwiXdHgUesBHa2dzsdcT/CdcfTJW4VnoZeNIb/LSk
zhtNgyjpoUZYrjqt67iHEJfgYz6bGon66dNlx0Xa4BtLwkrKTxpO1y1DGjmHZsjR
10jBxiIMakLLa8Q1povLL6ihw/fCDfiYWNZ2jwGhOijg/YV8TzOWtlvYTxdA2ncf
vX6XsXhdHCHFhJb9zk89Px1nacxSd7+s7Dj9XyLn1O1ZXP6UxMR9E1mFtNP41Ude
O+aY7yWTR2HMN/ajr0o3n8VK7QlTqs0OSpuGiqfo/Iua+gvQmiZnfjq+ayPfZ6CA
uqFcCz3zFVvtxTziNL8ZeNtQnmc1oZdevoG1YziK7w/fNFa6ye0HrrC1zrFz7Blm
7pVn2deaVgEetrSgvoeqlU0LqaCZGywbUwmWXHdE/swSu8zSUrDYc3G0TBUd4lvy
jZJjcgul1gM0ii2FtjoEDGj3dCfND4pbf2rXtu344TPbsLE9WO61q7Upz1Nr7pxS
etD7PFEG2x49FXOwnDdsWy9cPzupPO32MYGnApCcJ2TSWbMKG8U5BB8g5/x1X8Hg
StzaETFEWp39JXZCQ27jSGm2bOuOgb0ovAJTrH4TYVODfGI3AcN4eoEEcliaJk75
1v4W8/nq7Ln4vLF1D0MKddnhHrZKi7BYuJhwfhpTBlZCnY0+s5M/7DFqbdz0uIy3
vSgLOKZTXkXvaP+ubq0ikIeFyu9HPj+sfp+UFh4KoMUvxY9tAMad+u5OFmJL4+lW
/9sjS/rG6loO1jexTBwYBm8G6oLH2m9Mtq8YZkrkTepsj3l8u6/qg6LDbsBZ1sWj
KPrCzhLRiBXxV5kwewu4/8glduKfoDePO0UQCeJ/WCHdQZTrOuikPve2LS4/tfbe
KpxlSJZHukyxpX0sY0+F7lsGphVEhODbXg33AlVYly18mbB/OPUqUl5swuED0GwS
qEKObdnxjU/w2/DOJQ7y7ws0KIoHcDd8YPBubd+fw/YMB2c1eJN8eh9lRk7kVXiG
X2sLjKwhfZojmFW7wD30gwVrucGgynaHX+S2R8JyBGzHHkR0Woj/sl0CuUb/g6y6
p0uLzda3jQjAV2kE8MsZ8bso90Y002sW7Sa+NAwR96Ykmb+EBciFIl8n90wEsSa5
Q16X+fI1MwzAXIeiDr53g4VVUHjtF8bLa2HARJDBJpXwUFuu6pUAigL5J1FjvCwi
VsC0AUH+5cGqx55crL5FQ0eOI61XLoXXhNvnRblFFMX/iS8enwH+3+p0XTzOetCn
kWstWZGt9GC0F11wzqEcb8Gn5snvY//uPGEfO4Z5MTz2yRWjF38T+Y5qywfrA5n2
BRvfXpP31KVUiv6m0ONOFgpP/34lq9qcng0uSzNJOmiZH+UE2YSI+ASXYjGgLx0V
DlRYPh13xDRSvjhEzk7F+zkzUt3i+fWZtInRwe/wnKKoXsfTsZYtWF8VSZAG6yop
KAYAeqOJhG8uhaXzanL5mCPX8uAfnmFEtvJQOX3nt6eS6smcKbHmcftycPR9N37t
067v8vytd/ly5hUin3H+GV2KLZN1FafWdbU6/AINecyE0JnQ1Nax0S/ibT7zIpWH
gGxxDI0JkWybPBHKFzRXsYDqPVIqWar0iRG5Goon8+1V3kIH9aSns97ouHD3oX8n
U8S9Xrs7c2wXVa3xq7eQ3XkfZ/tCxBFe3SdQHbQyf2ajHXRoC0zRqXpc9I6XtYSm
89Y4lOTtsprahX1pt8YXvKv7eADLoiScvU4jrW0Vfai1d9P9hrBOBz9pchuo+x27
402W8YhgDiCfE5OjpCnWIDftZNx7XfoTvoYoBfN42Unk+BfSz2JWXW8zzhrFfYiZ
WMneiJpaj+XigHvyDtilLQ9Imd5d74nbAO2npEk5qdS8o0V8Kmb+H8TN72CdmyFB
EEWUs4J3Qms/CN2M+A/q1c+4fhN88QszCYcfqaH4rYhVdkFHahHXXqPlSLXX+p4N
lI9j1oJod5WpMg38AjUSRuUIh6hdtnfwozfXYQyfLkz5l0LSjl5gTpFx5gTa9Re6
BXRsZ4jfXCHponMna1uFp5/9o0+HGN4OLi9xPr3/sTLR73DKYcca9zlRdoK7DBXK
TyQmKo6/hqqSoboKhwvJm35DPcSilQYR4ODdQuetL4KxT+b/oIzLbwd7KMzJlkBd
vm/MyDe0apn9E44x0J4y1L03cObip3bwgXGoMS4SVZFfygiL/aUx6Tt5aliWYjW5
Vqjk6XThr1vPzJM4Zq1QrKQiYGryBub586/nJJW0FQlxZAhPu/h9vfxsMKW9MkQ4
k857llEnecj0Yone8TGECchanzdk0LlDDiB7dUx4yHN0Soow06xcuDJdTzqnaCeC
lW44+TKWAsb0IBG7rqUckskp9ATkBYdMZU/MvnIoMIo/+ltZWezS1upJ10wlKnMN
ZjBN+4cFiN9oU2DpG6tGg3Yb+4ALkXzTBBuElwmnpDHMGd6R+CcfgW/OKqxLZW+x
CFfYTssf4wkRoOw19sx271uvddO8BxCI8D4cmgqHZyjkBCHAFtFnq73UXuUVcimJ
LVYFRwnOoXnWW/AyOyAXnW1XWR7ArbIFoSFbWYrZKBG5dQIh0Emhx8hZcv9DK2/w
PMNK017AFYlz/zAkQCVR/AHaEZBzYgrIekqTlJvtek36vSK/NYBLPkdWWqCkrfmy
BuSLKMbSvEpcE+8pCow2fPFsz2/PsrVSZ0wPcyi1uib+ImSYF8I4lx7v4h6UdkcO
dxmVtI8t6Qqttg5wn0kLVOkUpwgFZqGKQ1RujzBiZQuK40Hrm4s6k7al7o3RjIOq
MJeCnksy/MViSFKuq5X5zAmat0OdpAWFDu9WBNtkrTtlyHt2K30Xv/p/OcFkgPYI
n7jYTkOOua7N8t10wPxN8Wh9xoUcyqlLUkuP+rwr/9BQ6aWSO5UEKHAeinAQnUQt
NhMiE5oLYrfeYLIzv31cQf6TvdBiKG2Qzh7sbR5Lng0o3cLRj2vX3DKGp23uoyzn
6Z6e+6f7ib1lYV3G38meCnGc+QtBd9jhawx8GcBKtC95lqYvWiVlyUx0wOmNNIQQ
tx6Ivj3rKx3Rg2e07541FWlYmARaSxuGK4oF5n/EFz0ZYDtCAhcW3+B1cFdg8HjQ
y0DAGG82OnlNJBsmJwdVc8FoM07ujgD5ocqGcCSMnWlzfdyHHmNGlY94c9l6eUiv
GLPx1vb1922FM2j4TCSKCLYYgXV/AesIrt5dvmDXJJiMe/0fAv+ZDJ1Lt+2sLEva
/93V1PiSW8IDZVCgHHfZEhQIs5aNvvG0xY8rXU5+Usv5E+qH30LGfDUH+tyYJhHt
Ftkq3/Ejb5Ps+A6ljRRs1LedJrwxLANSDJyC1+fsN5hIRdWW9pFQet0mUD8oGWB2
O9EJimo2BTVMVteFL6duPO5tBxNGGqGDG2DwhyK046FvvkF+9VFW5HREj2rBSwAJ
MkeDuRqo3243pHKHgYquEQZG7V1DAEVMr+2c9F+6awG1i+WOy76LoMcXIFPt9FXz
mKCG5yCZAxNHswwzaO5UZ+pygi3JupzePCGoN6oNVzdaqd2+4rtLNmRjK/V3tHfq
7/7d655qr/CeiVElSCdMcXwtNb3STVeOLEoOTcHSC9lJU+W8N1nPOZN6Q7dRBys1
PTYmLCUm7hXFZv482DRO5dzYp0rq4C4PZqiFPLW3HZWfkJORqJh9wK05K0Btc58W
gEAvFzVBWMfuzQTcgLxkqfszVIGxlNdjhuUUXjZMfCSifgRyTw47EqJif7KPxb4w
29jR7zOxi1qU+JuXd2VclQFmJdMop8sm3xVklysDxCkAdokddBzeZM7k2hALxQ7U
aMvRii0ewpNjwXaPu1Vb8PsvE7vCafSKVx6bHNn6WeiWYR8/RWB0Y8x8txDH4qVV
JTCsJSOPTh8c3kxHAOy1sD1uLCHK7RrSbJFqhsR/z/pLFtapzjacH6XWPyUME75N
GS2LOn6XGZos3pIlclIvknn0KAf7CZToAR5uUiGRVbT3wNtyR9oZlfnH7t+9GmFR
9Cif3NBCbsqRPjcTrH6/th87t9sPVv8wB+meNn14kACYrLGzFb1eO9WLf+YkvgIY
6X4gJsd2NKX8h7iPcmsxM7Uqavi8jpAS1Vshd9xSug4zc2bOUAlVn5vr0NdSYZ+3
Dzx4YlCghhtRNd8vD3NlNO6riDjZA4Wh255ZlX2vO/1uvqufFgV2NRtRECafR+kG
AlsWqICPoRhvj1l8dZTTjScE1a2ebrA0dXaXUXKbLb9C0IEmIbe3NDGa4SRJhYJ8
hxU6JEbkKudrVKbV0P5OQn346wh1xEidD63xQkAl5cpQbEy0wc05nACgXc0DLKcR
EibGpzNulmnwdWdAGgD2Vt16NrdjS43bYy7JZ8zT05Uv5RomPgZScNbMYSoCHW/h
LpKkpTRJPZ2ROxjP0+hk+sk3WaE7Oa2M7iFuo7pmDqfcyc2P4HTB8Nj4LOKCY6Wf
0aHBOp+y/F6BAYPDxbJr7baH1jCK2iD5b0g1TgH4yBvvKoZ/uR/9u6vdFNOztTzd
TubIXNma/rEnC/2SEN5B3aseSv50zxmeKuYrYZ91onDISmt7ImQ+YXLA6/Fq+DhL
qCO5DMkuNAvgm5kgs1/EeR6n/NI889QetIztSbXrPC7Fm1uNIDOJGBXMbr3MEZba
AG9ld6dYjTAX+s2bAPWRmUzePc218q865IdmHtECr/tzqCsqUhzMKZxHdaJg/T8T
mfzAqyBHIqCoBksCN8XPvIqqGD5ZzoW+kUWaLz1mskutK7lxWGk4V7MuXwp2TmSe
aopIyaoeG7hsicOoLLmIyEnBomrb68LDigswlbEE5qAY3uUVWPr/fxtYVObD/q40
O+gsRX+NwUrAGN14hB6GDBhSeUyoe8tsuGsRRfePD7T88E3TEID8A2pUzA1+QEpD
LHswjyZV7RHFquCM15QCu/b1FZg8Hnqfg8m+x8hIYa4Z7z98pOZ8HkLOMGs6LkzM
lwYSHadAdfBzKEN7FrzLBkG7rZ+IIUqIOu65wsN1IriCtQbxfKzqhQT7c5cEsfAp
UMRRccWiVhaMZv1fQfy+D6cldhR6eUOfEV8A4RsH8++DvMSEIqIqi0g/SD442JZV
SfyIojKCdOelAprfrAZbI/i5WKEJ1/qiW2D36gcJ7IulARdGbCV+7JCoyF71JLdR
Qkafs09p6GC2sA2z2tFCzHuUnpXDnEdK9yFRznIpJrBDnctYGIbvYAr+XfHrDy2N
YN/eSOCodERlXe7xHuiEGJ0tBZYz2qq+7j8YKre04bdWqIoGux9EQv5AQEnoPwVY
9cxqjzPhA505KqHY4ENN6xvq8gdGZA//1kvNBvgjH+D/THUMNe1vDZiXKNzjhUYG
Ykf3kgLTwj8S7Gr87I2lDe3K+2+reK18K2ZMGI6np4bxsJrrQRlsmronrwH/hlhr
Jn7mQZmXX1t/8UoWQaNnxqaIAtZD1xCfzrc/VGoUvC6955nxb2knQfcg2Mj2s+AO
X9UCqK2IDb6qxNbcMG0FN7Mi/HP5xb6A1+FhHY1eVLVL+00EWn1h6e3OaZ/RyqIx
T3oss5tWMXBXCRC47sxpQVBnXZBEjJ8UCxOPe3216cDtKRc5Z3i+EKvDNP14e1kH
04n4Z305f7fHf9DrBd6qyfqs4HGwzd9WNRiQRqDrx8RBygENse1SpUQrD1jGNpdy
70snvDTqACOEuWSCvfkgh393ndiKIaFcUktMGLrphxtkqsRBOQblN6tukxhUuGLO
eotUQgtLzqGUEnvdo/Y7dYCGU283BZyohgi/p1h3AciQdZArWPmBE7WA4akccsWI
Dg9qp8KuqWEMh23UKw5QTjMSk2xjlr8vGsPrHJg0j+1uxB7aGjgpJqXACYyfxpbx
PRmAQAtevWsvSXQopMdiOiYz/8UQIhOFfX4SgWshrTZF8vkB6zpnlsXu99Gz02Rv
WQaQzQS2rl0NhnWrcnRwgJEn+nwDnJnBuvaHrkzAS1f1ofdA7wb+7aMkAjcTHqGr
kFP7yhtWNtSBTWPdvM52z4lbMCGQp2WD+OtWqPnq5HyQuSnd5t6rFMNmV+839po/
0mmX2pAQU2GggtncVhFOCyqK71c1r8GaSPIFQHtFMqeLw7fQ7R+6Hy3FKtpKKR7+
Bd+bH+X22tyZhvRvb/O3KE3LhbOcs5shPuR9ptEv25dpsdgjTLdcrQlq53kenPwh
oPmvqE/sX8w9Qbz1LpEpyON4ayly2C68G7vSdhHCDAWK79hBsZVWSopSUuqTeldN
BMYV3zN67YVQKf7vl3Rfu/Rjv/t3DRT+Y2y3zajeZM28Ue7FdxzZD5EEOBJIZEcG
jJJbH5COZLM5fPy2ARWWuT1i1kUMqiWPr3EBOtzYLxKgVMJ4DDCekSFamEBw7DDu
K8RnggIbtx/GDAT+rijzb67nsdoe8zQhF7pbnIenfFH5/GyYg1Ha8V5O+3+gM8Be
W84CJ6wzeRncnR0dV/A16loNHPJNYQqvKOfAtD1WXFFdQg94i68EDZDI+/8nT06n
qO7HDu0guh9M4GTuMmXc9ssWbzaop5zIE5hm2iOjekYP5y53HLguJ08XQ/ji/t2w
UfbswkWQGTBg2dLW3hQ1JsRcjZRryP5iq0l+CiIPB0WPKhvidBtLck1b3TXtyZIu
NaU1VP3WYMkrTUVCWaSRFz3q+k0xjpxtSycS/dydebpYAt47+EKT4GNtJ97n9uED
Kug5ScTJBZ8uI9f8ndoa9bzy+/Dhclxdc5rvFdgJu1O75annQcWEfFzPSnIyQHRq
xK2YUlJK8jYwLffcR/OoAtZTDV1Xv/e1DE+h7JKUOqWT+6W0wVNszD+u174UfnGL
hjo0cN+VR6teB26cElleYCce6gg+94rf70MLMoky9Lq0j6Fq7/YrR8YfZs8k4ciB
8pbu/OnYfhSgwIuTKeA0jCtzqQcqLPSi5PCEouj9jBShd0SJhhs05Ufcc/E3nhpJ
NG1JCMwiiSA475lfe+HHnEZxifighmlI7kefWM1vz38MUleFY40jcWOyFjC7hnU8
L+pls5uuqLEqLuhUD2r8rdrk6VFVdjHbcyVsoH5IG0xOZTaxgiQ1SfhLh1Z7Vhxb
UHRcLCrBesl9z9Fpqq+b/t56LPa9epTO791niB2NhJjsNs9SiIZB00f3Hv/oub9S
C/rMGKLElbnvh8vciN8JheLwnETyf53s7mJZ9G7x0Ca/yjp+lUFNylXoF4xFk6Zh
xNUeDbeaMjL+iOtiR318WWlrySJt/bq1+mZ2u7ng/5bTKzTTY/CciO8CySevx/CA
8Fn1+QD4yknHlC8hw00gZyc2qKUIHbco7uEXtlihtnViIGAQzHhc70meQaYM3hsW
KL+9BMmZ8UOSnKcuQn+aU56dOVvfoXJIxc+U2ia66o662VtoksVH09NmtN4Q5Jxy
6mpoU4GD/tHsuIE/81g2kHknzOmjXs4sYpJCUbGpnR0pEvnS/DkH8dVY3L8JG9Gp
GD8O4Vc7xKSq873vHpjWp68lb6oMhQiPxWkJXyBwpk+56hJpeDVMrv+eSmHdt1OX
bWSGr2wvi9D4W5ztv7JDnQ3rdaRNVd3/XH3XJschpln0z7+9jG9BSA7D4a1Q5BnN
fps78nk6q1VCsGtjw0YudB/GcT+22bpbHhemcl2uO12OoyTgnFIlWwjvq7KQaLNb
4pYLjSl/SQEhi9m0FojyDfG3ORdUmOzlry4WiA21+yR65KbR6TW+d91nQNRQofhj
l9jw0edZRkVkGwUalGmWcAZzql/AnBqdR7uLbw6pZ3ppbU60VBwO2/dmLi0tkEqN
bj6+QyOAPDTkOJz5Oe0iWe2LYwzsiBsp2/94PPJTbR7QF1tqYPVEwJ8L8fJ7a5iy
UpjF1b763LEcmAEI4n4VQig/bC2YmTZePGm9x44VzBbrT4je93TH1jNrWyJjNt51
IS9PfE8xZhbpgiJw8UeIILuGjpe8oWMcwcXqkDFIgR/TkjuRTvMBQioeckIbgTVz
ed83oXHhoRrrHbWuOFmVJS+MHRWLQkIM8P5ZFL8j6uCSBkTGTZhBbqxketYC//aZ
/7oPfvJnrvSipaQzIGgUXt5pDkJPOzTM7fNGCXJZe/gh8Zg9SqwxFIwrujfylbKc
OAhFwPwTGNYAywYOexIyVsp323L6wzKTlWl3tFwZViLIDNvROMcrLnS6EBW3uSLP
mNSeu590H1wm7PqOBH45lrsSz/d7oNXYlPSLNbfh21b5H6NMD5ZalNa2N7wvrkJ1
sd3xzvWbWhd8/BAd+4vQUwUyg+XegSF2Fctd0+nvnKlbtycoL7db/f9rLosyHSQn
DYILX46HoQFsnxWKy3rjhLrzF1gYsB8TMBfHTYmBfkTQuFK0lBt0zIpsYLiUeavQ
avtIFQeefqWF7060vPf7GiveBuF/Dt8cuJ+oAQOPrTDlPd5stoO6f+dOoSlE14I5
73L2/hUYpbeTpmd5yLXqZuU9vu/zyR8BI4RyGviKxbHM7UIf7w49yXjfgfkIfbnU
Wo3rxcwdDz4evajdc7RZ+RreTIFdnevDPhr21WvctCq/enVJ4ftbibhXdBWly5FT
K8e3cUOfEy5yXaj5V8NYvIOo2U3wd+PHii4xtLoafa1Gdl2FqWLs4armgoyc2mZT
WnvyvT2qq9lwVKYK9dgtSpRkDylM+sNJgK7WIjKkQEWsKAXrlry3iMvNcmlMYBHX
gMnxzLHqJ878wpDqEQCKagyh3C4cbYuU9nylQZ2PTERMimmH4BbAgi2gpvdLo3AK
Ul3O7Q6YLkD9/72/ME30UY92eMERwhrfIA/CZqHXX/mO9iH/aAvY26Y95KzWjd8W
B2Ropw4RbUOL4vBbinXEIqio5rZ31bxRPUo32OJP74qLYiZjbecQzZxjnFqKYjx/
IavEUY11nXTl0zXp/iciTOYrQ10NTkepTqD03DcAjm9oYmnNmcUsB08KDvRv3TY5
PsDGHDAxQDLwlDL7nGjPuay93zUiveBvO5P1dbrljYzlcwDGjOnWgP15A0+GjCHm
sh9FJCIN6sz/ok3TfmNEtkYSxk2/51Br7XceObOwbwpNgAbH9cDfznsPbeLTMl5p
ltgGNiEdq1pDF+Tq+sxC0bBok0YB18p6amSU+cZp5OOlUGBYtwqX1V7mfIpfo81v
uNeD/XsMWMZ7oIQfCNgdENOeyoRtXgIk3nubxVHMYGELtLtXMkbcVYKKpfFCksEB
wC1wpYrhascipdoML1B40TsMByhvoteUUdM3xn0XTtXx9SKHfZWi6qwLvk3DDJgV
UOD/B/sCLgd7H92eBAqWF3pfRyamlzdKZ0DolRqHWxaEPZxzhoWFh6+uUaScSxzX
Ki9EDiQ8YsOXQ3isY6itEk5WAUka/t0xBtXDDvQVB3yJWPfoHKp+gQnqOQIqhQvN
Oyze3hFkNlKcIPmapYnJZPPLTXG78lmXrQx+SsFOped7kAONbbQIsMCVIJfc6knP
ahpsHZg/1E0NvZV5uibSQn8O/9pknWp2FZDaJqq3xgxqvzSLJFy/SSncoTdUZsM6
Ta79//WTUcyMLiNKZeZz0mKQPBHFXJ0IQpa4BiLZCBMzynLw3Ffod39Z7gBnjMZp
nr5srQ7A4Y5HgMT4Kkou0glZDOtsvkDNhwvE8hkzDoWi9q2e1gxc+kujIt9h5y6J
f3DDtGAV8Biszei7RWzYNwjHNiwYdS+C8avFZDEVinFmmzM+5fp23eq8xj/sGQyZ
a2txaceEuIYOBVRTdcKMq4Zu68aD2DE8sHyi5FAFtJJpB8bmb6LDSYC5dwxDWFy3
sZQ02L6hd9xMIUK48vfRBUcuT+Bk9kre3rj16ugdekU8RUvD1AbSX+YSK54mCdPv
rn4X7L1P/fcM1fpkVAwJHsS3Bh40z2oyXhTySIxnnf5Y+SHuoNjolD41RhoG7P1a
L/0YljTMiNXOY8dcmOOXrN12cF/46Nm5rnhZ0/trAOsaH+kpRfEbNH+rY19d7Ocf
ZEfpK4jTGHXF3gxu2kUmveh0MvEMplujqcCHPvbAiq7N5JRmn7w3SP5DeU8MJaLh
Oecw9mDsfxHR6yvBMa+fPwAvDGotUnkHdVBwcwoFmw3Q5npm+WD/4dpphcuWaxPQ
Xk1TIJDgeuTb0KXkX8MEinNFzeVgRI+vS1W3vMy7PoIDxmbq2tyLhkRu6b8OWf65
KQ+i5RN8Wdz8SPEC/koqH7umFKL6nNeQsvaPDAF/zemyO1Jy/9kaHeAXGPrXqb8a
RmzOVCMNVO/q3/PIzoJz4S435A4+swvjqTeK2Ixh3rTJTsgBr+9WqEgzbbl/HzS5
7ZHjFE4VnpbMBSmU71XQdDdooFBe1gvYl+ISZ5tG/T5fZ22JGTzB17hWbk6C22Fz
UIMdkSlEu0Xv1LKzYblpluAztgodyKLXkdodG9/mBJ6eT3ctkfPTrZzGWKuiWO9q
tZ7yEje0A7AqUGv5ssaGKBbiLLxklfZSa6bayJwNxyeumACcE/HiRHY98buIma/M
t1vp1uZ98Whqj+dmLJiMVEVBPbMLkIhWK6T1av6p1P3ixHEUwPK76SQ/3Gz4uOdx
PKVV4q5m9hW+TlH36BQ7WlpbIbeAP0uI+7sJasZyusao9q+FUq9kLXb0WXqj7Vk7
HZdBT4fgF1ArPXaxzWF+WFmLD1/NTTChvw6IQAWMMHjX8cKK2T1dq+P4pZTY4ZTl
oC1U3tuOkEcQUsglDcSAlZMCWnETE8Oj+PK6v9QCx6uPDqeJDEEhEd9exXu6jfVH
vRcv0yrbVE5RJ2A9WodjV7/mgGBN2iAF2CqupswKe8uztZXwNA6ImqoT4/TRHXu4
fQpc0Es6fQffX2/lvtPxUYSxRcf3b1LM2ulOMyuhTHSCCoLam63gMGKc/gyepb9/
tZIlceLngxkZMyoNe7JwvnvS5O5uzQ7W88XOcegOaAcQTX8ljyW0SGjGHz5iJKFD
xmYPCiyACjdaWmFgEiuwKnBDC/bJGzTyJu0b4wKMg3edalnCkRTEo5uKzKRrDqiy
tG0HcWdYasFBqr42C79arYJgv6XGBPUQI9UqKtuRVZuaFYt1OckY3OiPq391gdgc
pqWNtASNap3WnxXXacai5Ir4oI6c53Gy+JFGzijLBP8et3h3dHfhBqnVJjmS2AHL
05tLyjRTv+oHHr4Hl/Iqe4lXwMsHI3ka6zIfxqvMGYDWW/eFJITNgaC1mYqzRj3t
KfsSkhc5lIW9Gi+9sh30NF/J4AM3fieY4N1MS5GvPzDVdWlUz2HSMmzOeYrLL2Lb
Fbr0/dKTtcvEs1gIte5BDWptHNU2edK7W4bmNAURkpsu5E1SpOj/cpMRypLnntwy
Fydob8pa6ZxF9WrtX4N6rtlZgqQoBygzXwRKjrIYXMr/ZB86CG4POCI9Hl2t7Te7
ZmNBGwaDdKnX6mp0KT+v707foJBCmXFxGnVn1rBRspd9KBCcY6JfZkf9zTGvr2oc
MzmG18vh6+VM5sVzWbDQ2qhag/36O/uHFlJN6y0R89dRwxAf5LVLZFZvNmkl5i71
aXZDRsLvlbA/KHdxDt0g1K1ArFOBfLPgURG8nO/xqFVy5FOEeBDKtuPqUsjgrTDo
H9jwj7mfBeMmk9nkMEMyt9RYGO5hjR1Cx8+a/LqL7WAIa1x7hif0/3eznIujEmpZ
f2lLGzeRA8nBpeNct4y6LGlmVLxc6lUmFCHGJ+iFdX7QCdkwrrJEPeVkPy/CAu9i
cn+d1BZHOsP3gdD+/VSEdcsUyWjLiIkdLN1RfZCp10smm/aQJTFRRVwbazAl7WWp
Kfl/jNO5iSC3rLzUgwISUBsUDVBgqpV7VB9Gn7cmCVvFeo7/oo2skaDOT+r9x6DB
8CoEKWMLVLafM8EQSUB4W050YK41HS+vXyP+7cYc+KLh+AlZ6Ux+SeaT77K9QQT/
4CiPqqpf/ZibIFw2bJZjm0K43wXudtKAIEofgy1o0ISSL3p9AGarS0S/mkXO5oA9
dYq8060qkMS3trti41Hk9bUyZ7NcVzTX2IejhI/eHwfOUU+HR+XUZnDjFEeQHYHf
joEdy+sqT3dCu6wYjZ48eNnJbKD4zGMhWNQl/SkucHzir/Ubg6lCKZc3+Zl/wrTD
8tFIAWSfWsHT6OATir0nW+tIwYEKgzQWILyS+GaZOa3OlO42J/x0rIpD9oj0tTJR
2H6KtK2u9ATamU8JPbbhb7811TSLxyeu/m31zA2lZ7070ICTFaxt7xUGwLi5kW+g
Ybr1t4PHNG1YwCtqCQVXOkIrd3QR0aIx/kZxw+Wl+sR4loNOX5iu8jHLA12+cqUY
dV6pq2wFeIFD7RXOg37GifkABZe04qviCx5JAvrE4wC90tyZ+DnYta6kyFD0KWER
TeFA9UyZkXrMb1KjpIgNV2m8aeXQEGWcieO6UyVznZeVEzZGlcXEPffBqzjlJ9hW
wc6G+EipRwrMy7WRaYzFbhprN48eKtftsH5Nwoq38yAlyR6neUlQNSbbnhZNqm8z
Wg3VJx13IUN2RYlgPICFBohBy3eUvEyWtUW68qqMQ8pUk3f0MkVBljcnGSbs0bdN
FAVG9n9nhlxBMNiCmOIABeo927ZUh1f5jyxBixsmMPVUnjBRHzbH7a25mZvR0s3Y
BcaEUN0eRdOy9MaclGw/AAYFcvTNaPvb8qiGQUUIAzAiKKTPD+Q2Qsv1WMY0dS63
luOzeHk6w6bYq3S5JyPRnzEupfN0cV0j6op2BynJbfLIpCj77rriWrqVY8bxsntk
6ucA99i+/Z1AkHe6i61dvGVHA6kJStJBRDGZcDQ98KXu1nm4yDefVfJLESsepW6G
I7ocLu+8i81Y97bEt0dIWNZwe1j44kBrKsRPsLcwqQXZ9cjFOcDf2axPnijkC5Lt
Frvkb5G9AUEnEdwN157G6bV6hV53U+U/GG5Zhgiak8/Ov4mYYa10vYJ4289B2KZj
sy8oOSvYH2ETvvT2+axyOFJtQ4P2GBKk1r+kaTPkwmXNmb+HdhkJk8Qi9QJO7zUk
hzOTneHh7jBN6kiDw3G6aMgGEYVRvS13USuL/Mc442PzaklPZ+ATby6pEsi3w2FV
roLe4y4wgCz5svXp3qP9gXckreXyaJ260TaaWFq+/hWj/ui71ssbbHZfC9sVdj28
fcShyImhI0s6TNzJftHbR30stOXJlOvpMzb94BeGuG9E8D+XzFbIkW3qVVJFKUJV
bL1VEdsrQ4Gzti4J1KH0+MfysXAWyV/8NdtTZfZNe+pqMLlm2rusW400KCo+AbQm
KDqv3Gd87syjYHAz+Lyqrk1ZdzWFoqXO1EdzDnuXY0IZ0Ct2oFuaKIM9VqvQPdjC
BKdijwX9I0+gI5dezPDzn4P5ksuKa8OgXpdM4CQKB9Nwm6S4g8YthbkBYx/G2LYf
FdNPQBRifM/2n7t9kJg9bJOQNMDwGvuYfS0yvKoDvdi3EIg+OYF1il4VaaSCCTlt
j9CXaG4jlXXlVw59cF2DlcMzr1xwRoR15cDixj3Sh4wr2LRKrU4Opa303Yv2yhjD
RmyqGlw/rSQU6vBHQr5lYvxqrYi3JlkfVopG2qEr+ATX0gSHVjnVODl/lQviJh6D
OG2bARVTtC49NEhQ15jx0K+LuyiKykqPJyqY9yUf2lCCkEg70Eysnx3CGV9k42DC
VTbiC2P+AbqyIeTAZK48x0Nff0o7ZLVugziRMJFm46o/kb4Y+W2yA7M0U1MQLFK7
W9Re7aGeh8AL/7qcDV/cDy+i8IVA5YhvKr2PGCgj8x5hQo9I2tJfpxfML+5Aj6XW
4VIKAOhsTs3VaoST87uJ4uaqqD0gLQbPhbAHEWlS0Uh25eiPQ6VadMuGGjoXFHqu
9yEoeTxGVK+mT+s+pXFo5UPY/NoThXIJph9YiNtBVD6sZZSz0g2X0ZplQlrBnPCa
fyB7bl9toOtZ0qqtQ66Ur3dprNKNreA6Jq90QOroZqogWOs4Zb9gr1epHsXCNZmo
uoedd1+hQJU41uIsnZ4XhobJZu0vgHeoORZwspZgnhvPkWmMpYWTNfhayJ0nJ5Ti
pL+YFwEFEbggmaDVgteoTYeppTJG9wI7jxJmPPI/cJ6XDozlJNq/O1jj24lmGsfi
8b01FUvJ1LbZCJgjhEavtsQt6BJgEUbyUN2x9wyM4Firldb7o8vca584YHn7VvwK
V+vwzIR/q0ysst9ozp957f9aSTWlSS0IjlXfoIhYXQKZkGve0hhIQWdb3bgGkALp
r1rQwNpPGh6Zz4WYKgbbIY529bmgjb6GUQYbcNeijd8Tcd7auja8AvejDxDtjg3B
UnW2iHgLcE1zObTBMcDK7pjufE4OnbW6t6ug2kDaO5d/fc7ovGduTq51lyjTSU+J
dz36KmZi3+jXVMDZSHSLy9+wuZeBLygUd2gGZa5iTNyioNxviB+VcTS/yxVtjfko
j5IXDyXRP7fulrt89Eq7Sbk22RQBScI/s2gZLOpyE0E25Lo4XSHznRTw45RrzwVx
vADymbs92DmgwoP/LcDmJJM69adlf41JomBaEZTCMQhLw0ISFJ26Z34eyi4nHHbF
AFrFVieoPJF+qf8HsYHXpfShhheN4qiphWukPuwSRM0FZq5ZTla54CXTD/dw3axf
0rADhzr3iYSRByFwpM4N5ghONdYVkFWy36alp4q1J1dO0byRqRNI4XERNInQCeZP
7/ELiohNkxHsh+UpseN17grNIWJmZTDvg1oRgDMDNYcLsB+5abX4DxC5BYHiiYpF
Fdac7ispAg25WHF7gV2bMu/UGBNuSkwcvQ8yiXHObjpK5hPvdkAq+AbZRLPCgkBY
0tlTAuH0vZHTT3MnvH58y43tS44raOrrHlBf/tTPCRHXmBouKbXDKLmcA05n4Fef
1FJVzZvK46xhdfkb9FHra8Z1SDe9Z45avoh1HHiN8jgAX5CyoWsacs8u65VikCHn
4tDVt7cynTxpbTqNlyf7DkvoQ81SGT4ASA9L64QIbna2eEWJjt777x19AOlGfk9/
xMtTNHcqmLkBkHMi0t7DmUsMeF09u4L5gGhdD3iXE1ECrSi83K/f3MuWLTmIMbiC
YwhiSuObhGo55GOajSV3EVGB+BI6xzhrjslrJ2KVLBvFH+qWHMlANYAfc5FJKwO9
XrV7HxRNIENSoSMbn+281TRkwrzV3OXljTto2zBjosFSauKj2gHqWptoVD+TKMmX
OKky4x+Pbfk0DOJ5vqi1yjRR8TiNros7ztaNXoSaYa0t2t7bm3h54VmOzhrlcC8G
CSAOAsTs5PHUcNxSKYQ/VSRe0mhGxgmVM5RcfMA1SxJOpuy2mor7dFdUnCMGoSpP
m5kfzKgZZNIziS1xi7V39yvasMUnWGigbwsoSZJghpqh4yyrdqiBRs/DEUbSEUH7
gMewhYERGDxWuSh04im108LuxJqZ4xsS9Ehd28C61bcI06cIw8yqjzIzKTHzSHf7
mW7NizmWUx2fRjJfoz8o1jHFMSeBgC6KesoSETgNQ7Cjzk91fQGxSDjGl9DZH8eP
TrcLEMGvLqfXOpC/QjxGd3ZEBYeAsQ11pBtpruoU7tU7WNhGovJ3LSy0PFEmKqD3
7oCf6AJ8hNp2qHPed6xl20vmm/HVisNkALU+kmaG8plCMLW7euKMHAscljYdXJ8q
9jZBe0gkHb3kY5uvYCNuc8nBAMSjxlpnByKz7T6vVTD2Upd78ryAXpqAYW7M+x78
APHhytzuTf/V0c4/ny7rfm1Sze57i0ATytwPkCxpnBLz3xsb8bydPfBPLi31v8mZ
oTEGozC1p/QS7CNokC2n5FfXsuXNfqLANhDkoOIPAh8Ecgo9blrWG0Cep7+5FJfO
BBrf8Pd+6cVJ58Jgv9I9xkLyR8wH43ufF9jO1o+jdMu3EEDpMZAjsKmIjBhPaFzu
8fWPhzr7M0+udLihE4MgtxtQFwpx4fu1sLUjD7v6cAyM2axN7N8lvQy+uL8Fwa6M
YXKMf3F+c3EyY9bo/+qe3eDFHKtt0K05rf25N5EBq9DmD+8IbGD2isqAHBqmFqLM
CS3F4wwFk8R1/FZJ4cPd1eQtYVJo7f4N9JAgK9wo8eiJfqn7s05gZcnxwIvoyf0m
v2cAdTnjvHebi2oQUIz9G0xeJ/NRGssrCIBBiFfbUSbLJOUskGt1Bk+xiIVFD2MB
Ejp5KkvvLFovVsPG7/zB4VvjX8ro7ei4ZYRvor7XkKQbonEIusvI4LaI8qlVZGJ1
ER9rjvpc3HDwvqHlqvhxrs49XIVWEk/cj3S2ciYul8mEzBiypHn23/N/8JIc/UaK
E/hD/besT/DP9mcvTudtN82w9SXkSxdoeLfRCpnxSRDZF8ilQUiNSpxqWOLFuf17
culLM2ebixU+sdi+aV+d0K1F9iDDX7zUJx3ZpE2mi69jPAHEaV4pAkB0B4JtK6LR
uaDDvZMcd4nAjdGtrkOOvOwFNLHii4Zv369BMsyKbh0bqVCcWo08++dAhNfAwLfc
SScMLgw0J+q9WLbEXoG9nS0v49irvCZDEUXlfE+qNt/dcJICHK+42s92djP3U1s3
ePAI5EB7/D8PGFe7safX6YS9KGPN8/zRtP9BHPgRYIwkg0L8Xo0yniQlWLotqiAT
6qm3KAadnGqirdsCeOZswYP/URDoihUpLJkTV0aKW+zcZOR5GJFH4UVATcfJ37zt
ifhYdIGXw/2/LyDvKFuqPGnsf3fcrYgpH/AnX0dKbQAFPIzpf8R8cZaMkko3+CgM
PoZhJreDdkOHM90y10RPlA6yxt3Ng4IKIfb13LZJvQOi+yNxhq72I6JX6m4oCr+D
/orTDQJdkekW6UqFo9aoA3jNKdMR0WFvdp61QlzggkYafq7xTAKXp9zR+wIPBvKY
OilFbNn2zsqPwlmeRw1drOKpZca4LzDae4fxd/qzYpQHn/20tfqQwZwPFfxWsgDR
RSdM9aJXypAcG7Qn6xtKyOqY9qotKG1muG/33nE9zHasWvD3R/t0pdy5+zLMlg5m
OR31WijSZf2XJmiW7y2k0lAbg6TK1wOwy7IkJCH4TabdMogo5BN3t6GJVNMtnA6W
EYaQ2ZOhN6B5DZL4it9Qok5yG6Exgjv4IRWYrbU8W48FoIzH91KEIkAVCi5FdSXw
He/re0Vv603d5STv7fyDu3lQmmjqWH7B660CiWBr+pUl3+H6snbewh3kVfIdZPGV
SiwD3lliiS8PjxbxlwB6FSz8FJV78VEUC2eJ9KeQUfNcRhYYj5iav/z3X1HwoTOg
hJrkSotb+2WngFS3yXw5eJ0mMRSZT7kCrUB2jkABKLRWiEwhOpjlL9PCqz0K9xru
s1X7BSa9fa59WQn6j+yPEkGn6Lg0TvetDYJiud8clSBCECnF30fGNC3Dowpsqcxr
zqm4Xki2lPZGXsjrdVsDqX0snf93H69qgfdX5u0GD5rhE9ZDAKIi1R7j/4zuSjk1
yG/wGwneGvdS7COhTHVPJ4Me051rGrCDFdvJ/fkDsTSTgXHpiSuQwhqzDMD0iywy
A4petANZIQa+SsJ9xwx7G9nOniAcrCpMbvWCUVS/Z79SuhYm4Qe9oB2X20H0dutv
8ESh7UJ7Ikg76WLmxekVMTCWoTtoQWYjADh+aI3q+Mbt8FOn0S2VMgmvMNY0cC1p
3V6OExPfXfdyyulLZoIC9tzu4pdYY1pQ4iI37pkowvkiJyDvipVS/awJh2h/T+hY
XR6sO0Nx3knAcgXVerW5HBsl9QP7x1eJTLqEo7uSvfJlE6PDGKcekrVC8B7TWOnZ
wVkdzn6nCSN6eXcYo4kXgB3VZuXpe7lsHVNV5JdyRoewFNvLVtL8qQJvRHthfbBi
ShZgu582bqYAIltkqFWT3YuoSFEGg2OFtiCqY98nYQzEg9qeUOfhn8voDFZe3YM2
7xYx32g3pMpbFJKiuQvNb4g1+RIdLkVTb+mny8qpjukcqz5WL8tDSYnL9ZSbzIMP
LaYJIrZ3loUZe0pFRgk6x9l9tVmFJ5X5EJCaZZhOIQ6E0WyJqrojcic1hWIkqwKE
uEpWJDMT9GzcpEbPiZHQT+/Hi1CXsmcf+9SmQOsnCX+wuDLpFbw2+4a4yVUFtDpM
vIGHe5Fr3bEoQ0dagpRdePFJP1eV3BELI0sT4IqAGNUwsSr9lwUBWnZpxIS7NPVd
Nl70H8iYkDPmkc6FbVh945pfK44lb4oLbbafPtb+jzPaPK1NXWsS6zrKcMbOz0mS
UmYV2FQ9b41BFw9/wiOMuBCo9dIIiuSPjrLL+8txcrI/mZHdR4mf8g3THSL/lPqs
wv7jTF4Qrj/B9mtwWEHn58haohLoMYqJmcOA+xQAvkxSSCcm7HiaAMlnwRjHnZl2
2jkSpdPQdw0do/vM3jJZxVY9SsJnZkrSomDfZPzstmpagqtjaX4xWb+GTDIOgAKc
A8v8y/hEVXEKg5J67nfuuLoXrVpKfGTv0BvbMTdBWAm/KtRfyQuq6wxs0/E9M0Tn
vvWrK8/f8BLELYzOC+Y4gOeGr5mv8JRsJkaIfgDREE8ARJpFMURihd2CXW/Dl3z3
T5J6UwdC/0GfDLo5Sm6mIspfRWXkOjVXUXyVmpkgjbldNM+hDSEVwFj8zzS8pPHM
tGPjXC62iM1oW5eUEuZ9EjuekQvlJ5caMxDBq4Fy4Z2ZHsYqQpxwUlzp1xvUNnBt
5aBKrrNS6TpOfXC5vIa2FVP2MfcLlZmzBsoslbA9RPHQkDONMscogxFbKfg0oIl3
lXNFwbxthL/F4sBBK05pdn34gpaZygCkfELOg58DBz9ZF7iNGT67eqn0Gb1n9Jwv
f82PCSmPkN2h+MrLDc2xmxkA0hBC4vZ+i9pbwmUWvDz6MpbCBV5+d0Fpymoj+xoa
7yu6s1XQQJYTPQrFYQHPjn7kHNY4oev0nnoJGi66JaK79UX56fLf7Si3y4G2y/0A
0Bgh+EUoQ0ouibbPJk40MVaaAOSea7EVp6eznVeYweBYNATQWxvv+TdFRvn7WXw4
Jxe7VBnt0XrwllZJhM5K7SiEV6qY3Z/NFV7+aEBVP7aTwM7pulwcvB6OHRLsWvnj
R77zyiD7lMQyvogTshejDb7VIvS8VlxnwxvcHbOi2M/cN0o4I3ywS2SSQ/Y0/ipt
fkgwxYYphSI6T8f2q93NEHDBDEPaZHos0Gf1uAseCL6NIvosr3W3H64WNTEoFOvU
n+gSJPi/a6UOI5kxR6PiWctUDD/4KNAGxWgeh+NFhfB4qROzb4uiJiuKNsU/KPw3
4Ud5szIVUUzccKf+cw6ZQ1QE24fkPIRUmeHmTVFOAE3yFkOVmMtfpBkBAatYHLoa
4Rymb1YWnH4ndfByHIKo7h6GJmzRgp4cWzunDz+3GSvthMNwra1OVAw5XFRIyK4F
IDj5HN9zDFXZo1Q65uRY0nO7MTBP65XO1ZpdlwOrMECdzfTSZ8PgHz4VO+I78plk
IUY2M7bcRT9ByKjPp1JczGchCjg4ld7jEIjolRODKYzbXmMsp8/vUbVNJOoc+t6v
ChulZVRVNTdKgDRIdGQDECeipIajKilpv0SgyL94Aqc1BmlDdmQGhhh8HO7Kf8dU
fmy21UDu5dQTVtNol+quffuHguv91mQ98OZUb4Vt3dmzPANpS53jE0JfburP8/n4
e2QDXatV8Rvu0GJfkrWL0lQJmtCu+m/3ex8FUS4un2jzmiZVTZXVSkUHmnfSc9jD
+3Pyfyef+FUfTC/GOPqxkeDlgTZ1LPUFVJscAxXsWI4s4kQV+JA0BXoM2ta+yrwg
mdJrsMNL57aCOxIPXOFbbg0RAnvdQP9VsRCiIaWIOYrZvVC6UY1JQa/9I5O0OrUl
G7v1VSagps+OlI4AQqxlFGFOVwMJqnPuno1ejefm1cFVOiToppOkzZSMfdMg5yzE
qzW/FRpjUcO+qh+hI3qVSE5gQhzvTnkcz5a2kEpjW2+6747RfsRBfYTLjXVidHLc
egth/xg9jhO7pe4wBzk4ZNRZetPlsS5f49p6RRSAnhvJVxy3JaFvSydkDyv+aMtN
yZdw8G014jRT5UfhQbkQQgoW7nQjEmEnFEIfX/qKPPDeIDUMNMQj1UToOhHGZ3gL
/Cy6d4mypWM50RiH2s5F8YaNMiTMUPTZIvkJk+OJnFWkPL0XB6G5kIFjbzTmKklo
lJMkGBKZ+bteR6mIufq1B/mcJaGolRU5SHNA94W35PUKvHy5OLqHCfZBDbWCIr44
cVaYActDqXBKLruQLMQylk/IiVV/B0yX79GZrumouCMm5a82cUmdRXgsiHVCSGe6
3YYrKkkv/EheGJLhW6bR7eS4pdSSTfMxOd0vGVqhkH4T6sNECMQdA7jiSszfPO92
mlFIpOpwAlmzP9dMNcQ+vMaSsY+IL0vXEzybMkgpN4gc26RWYf4ccRxMktH3wjjn
hLd1r8HFRFC2YuW08udDXsTGtEnQD7p6aJd7illlZuf8KQUYGtTaZ+oi8ZlOMpxK
en65FV+izNtHtETHcg3xvpbgz/6wvR8RvVeSMSoEuafAq29ik/CmdXtBmHP38HYL
GKbhU7Se9u5GTAOUu1wLpTmjEMDrWaflhGWNSP5ViYrooa8BfR9ExmoskIXz5Znd
V0cpNEvAZ0McrH2L8nzEKcO98nY6grZfxQ2EWHFBTuLiujag6aadjCXQCAWr264e
GACybOZoJTdzC1Fyk9ZUkeUfXBRmOLD6qWVJMuxZWmAioNE1mZCrgPeXsmw68DFZ
rhbs2nFDzP5mpACqxF7KZDaEv3ufAJYMp+DF3LH0I4T5edb08rcLcLK2eT8u1zj6
uCtSRo7qwnxd9li1FX5cWNw08IliBPxbbm9koPMmJwobIcdsT2awkEbkAT1mw5hG
QKlz3HgR3CIiI8Dm9hOYgY7m/U6oMxyL9atbPGztGSKi6y3RdZRoz1sjBlCV6Qji
b6InW4TsfWo5pK57h4NI5wzYbCG58SiKX+u+JRHAigxpoQINULOBQxjIMPqTt5G3
PmAX2ykNMldweU+j1FK5GFPxdTyxAzX2iG+Qv35hRKRZZf4PZNaI4vCB7znzQsL6
QPXONRxSTzVcoq1bl8tx1f834pkl0UKB7hJpqH/GGVYYdBxZYB8QSxkpm/W0h22G
As72jvpPGekeN5fxiC2CKW4jDae+Zu9ssDpzlTAqJXkPsbKlFGoUdaq3PNiqvRtO
r154qTsTOd85zu2/nNvsRk6dLBwgn9uWV8C6ybnbcKDkoPq9UU0q9/kx9wE8zfQ7
34GwMB1FUq8aSbfBVY/TGUqFjEhO32l74oLBt9Cgc5189aL5l1IPdLyGs7YbNXHx
h0/c42bKBM967PR1D82KW7g0n94/pGb/R/s12I6WcuQj67fqGJcwYEJd8Uv1raQ1
NPouVFoh/QgTG17gI1I1v5j+0yvKpvsVtHoOlkaN/0ED6HqxU8IMHGLCrocAi2Uj
iu9tPCQXd6P+qdHLtEWc3FgDBWdc93uFC2FdGpY0iR/txN7YbCXPEda2OZ9IQOFU
YSVo61XnXE0b4xI8opFDof/nwHKB/6dX2XOijF6OvBJQg+CMBkXjmytiC68FkRnt
yW8ru56AlurkVIZuGfwIXpbia1wqAAi98fyeX1GzHuyKvT77ikZnVccHA9HkyoIT
g26r4vprvXqupIAW3IHhTx1vbcnBEe5EHi3w0S6uw2tKWXWA9n1XTngVOmfUnXWh
XtiaGmWbzBJBDD8S2iNp2pCyXxyHAM+J+rSZYtirurJY2LbfmIUWGGbrSAOvGU1+
YGRGfmUHIICUddHTbYDFRZpwLA7CdkeUOFYkPnGPoFsR+NSCxXVKWiYmfESh2P+D
fhY4zR/UM2fe/KWZndwpIGc0UMHOgcr3ldYQFMX7Ifqbw0cKJLgbBJbZ/8WBGW3Z
O+lAj86+oDdEcw72XGy+W/A1Bqi6iXRcsFNmnkBgZVEZgRA9tAMbWLOzVpUkNvZk
F3Erx8do9+TsWnCe1HKKacFcYqfTP+Zlw///H/VxWbgFdncLcpebEXH+iz7FRAw5
srhz9jKTwX2LBsiiS8WtfonRY0T/Xg+RmbryIWNsb1A2vEWXvbNLfOuYuMIRhJKb
jGbU8vZxZDcqn2uu/7Z6i5p509Jl3oxwPJGq3OX1GHJ0fb7v1BmbzooQzOmwjcg/
Y7V+VJVvRMMWZwFeWKaGSJbZRFMBsf6ruH5MC3Q01wnfej8kybBQM9vhiVnp00f0
hHnNasxMKnwQaO1oL3AsO8ZFlzMv1Y96GljIg1c05Kg/5aeg7QPxAgBentL8pNH1
R13+6X0Z6rCeItANOoSBm/w2Ux9rbOd+V3ePIG521Homz/IEFW2Aqbd6BsLERLiW
HzShhw4r6OxVcQZ6JOVLuk3WgN5CLbxVGVP/aKRtpSxWGyW5AoWOal56cOFO6pd6
yLZEqJ8UgTWM2dOfcZcSdxgj94yTVggKq5OWu4baH0VJNA1oBIRLSf/JJEo9YSdm
PvvqfZrgJbyDRACPViips/446870PK7W9RTeVPwvSJXumVFjNBamWvxGov8ANNnM
rE9bTiOuvxACv8jL4ckopuOR+2cxNG0U+3omdWOddgDGFJb5F3rxCA6B7uJymspO
i1qq4vZ74su6r6c8cSivuUlaiFciCSmZ0WLRIzqYL5EPU2K3gau5P6ValeBSr8/4
FaaPPQ+3oNaZkW4J3SelIlKxlWjqbBbPPmhK8btZZq2FgXLt0MrtYt2LOK1QctU0
9A8V2HOW3x/nIAvlcG236FQWyyJ0KebqKPkV9u0N5iUB78gpwEtz6aidZiqdp/HR
V/zWivyWNsQQ5SaeZrHButTFRoisU0TRUhvrdvTeWIuibJ85zuij82tl6wJ5Ny1t
uXDRZ+AbrAWKKMlUOoD74xBDPh4p1QB/b65wa2teUJZpfw04a5t4E2nyYtPPa/ng
KPmvGZeqWqs6oUKHC8i0njGFTYCPBHexMd/O01yAr/cXDM+E+8CWQC7n8WCE4pM2
7nyImBMFtHT8zqPCK08Q2V2C9Dv+TuTv4KIO6uMaNWQjr/4fQ0SbxYMRne7IiQWY
sGlWHQVcANCCa6rjHwKyXJlfrup7al5OMMX7fESlIYcGH68WQO2juI2p6dUKOTVN
Y7sncRgHbyPIHogq1Uhm8mNx1vjzck+7KfsVzo9guIkaitdhbHmLob1lhH1+3rRI
xLOl2R77NG9ipg3+aMMRBxc4rGFg/Klf4F8VPxvDMv1ieNLGn/yK06hiWllZUv6m
tcZ3ergk9AFsHRDCFibVXJ5GzWdyODnEze63EQyFY514CtlGvSEZf/MVAw03VJ4X
fGDUKuQwzHVq2jql4OlUxnOup9khPK2dv+7100+IIMCuLa6PUv/8Xk7WJ9Mx20Ox
tz3sx7059+NgeJEi4EouBVL4Xhe+Vjns7kif8E9vLKxDRSRBO47WaHgl3nGqNf3K
BmujTN3KhdCE306pNOpiVrwfJ0+HI1AGbiwmo+uZqt6/f9gpPw27TGxw7d2HRP8j
O41YmjkHDdN0LToPieNpA65ycFUM8bGm1TJBd9Cl1P1oVZmH2jtdVxh6kVHCL+m7
Z/J5xdtE5/h8ZRw7aEw/n0a3XSadMift2CmEIAMhFLhLl99I1vHRyCLoKCTF04Ug
six2Oipu5XHvKfeu6wYwZ7aEgZI/p/dq7iZrcG3dhFusYroBXuHiVb/cO2SUXUEk
WQVBrfD9WgLUV+ddAIouHzcrNM0FGDPyZVV5hO5IXLcreqaWmHBKKl1CSAOYRJBk
0Jf/b2wrtx+bkns7Ed/tmFXGEXaTRaChLH8buUOS4jMK1gCpFWRK9QB9UzMdeDF8
bu+EOBfP7vF9k3+dL331E2kUeCJpPXMyZXv73m/BImVssqTH1p2+R5tSxnMKJBUt
b/zbr4IJbk2NJIkp6ZNinjBTzTYy6Rell4plnOFXqYvMUJwDVzoiEj9SbSi5/+wT
N9YVZtYEImj6AtOVvHx1cD2gzoCW2NWE4AocU+nCuUMSHKw452+vfIFB4efjLmrF
SSf1zn6y7T91Nk/fM9QRVLDuBlUyRLjlR6aZgwXnk0Lv7ieFgZSs5zxrORL5nnoO
9e3k5ynYVOFUImhNBKM4OfUsWcp4Fq4MOckt6RcH+auKKsI3SQIIddFes0wqDI2U
HtkzJg7aHjtruuEbGUkYYwdLYleXTluZ62iBTyOwuJWhqWGTInZy63pUfjjcAseg
bc68BcvO4XzRZixRwzDM30Z67JBHdsSaS7SEgt3Bcr05z5pWr0ve5ZAb+z2yzB11
vyCU+HZcxJHFtUNYWdAdLSHzKy4B13mZoaBkzyVmCtGJfwEp2nGjkEwI+fO2fSM7
mDFeARPoVO8yXgFw+GyvYMy3oD09zoHNdfX5qOK3SQKOlFrp5XqSx/rp/dEyAPlE
SS0PZz4ttB1dxJQqkc63DVHljsKVYX3RLjzfqXlen2SGiD3+KoLzXb20A/FMB+/N
ycfau4ySDlb8do3176R3QwyITX2fg9HuAHzYvC+NaWTV9Da3kz74jiZywNEvdnW/
i/UaP40xhviY9cmaNOVL15liwDe4loeBb3ErE0gf5xZfVer3s1/i+lDwehLnAAIC
TDLh0rRQeCVU3fYbMdXgIQzGGUvH7OfsmnF3Qj61l+QmJ79ZqcbanVDHQL/00gcF
WO/Omobg+oUj3rVijQMhw9LDNlC/Puj9qgwv5KMALR2AOLtFFT+mefQGUo2M1OVR
N0vu33xNbuIifKk8vNO6+cpTSbL4W5u30jJVC34c3LmM88KDFcDSFrCg+P36BjGH
KVRBjunBEEi/ZICbzJ5v3PAA5ALCaahYHViujmL7KHwQOQDp6FPwlzcS48zFGJCI
DznLETut6XQ4QAm3714cjQJgKHzapkE3/5X44qtZDER6bmuG84VVgjFtubtaTYoE
bR6y4DnbV50UT2AYGdrmlXoQbFgMnAjmw+U5Lx4Y33UbGb0IU5t5q8LpXCroONEw
YcUFBjWXKy6SCkEv/DOX2hbqcp1LwF5Qp/iPHN1p4eae6iycQWn5Skis0oknizKi
azDMEQyiLT8Ba4vTWK/xwYaPvj3A6ofVof5AN+qWWOuoUtl+lsYbKSsXQ/GFBLW4
75KKvOCWqbvUv81ZFABsWvz9B3macXE2e/21JvPGkmnGO7OaDGQVgMtGrO4lCBww
0EIp/EeAsT45wZEsM49sYc6bs7XSLNOyjAu6TAMcNBkxJJrTCKEBDKSnUOvAzVDb
qDivZG0J1UiYa0DlG0rchv4Gg57jEuHE5uSuMR8Ai3Q1NZKL/zccI1IqbwvCNS9G
4pjvPgGnucdS09LFKEvE9ydrVC2MtQzPfi/JPWXKqKqR00eH0wxu4lH0HpqBUTp7
u0Qh+cwq09CFALtMOHynTYUrv0GYPMG2kO4mNqCGeYzT5bY8NbnGFkKhOaQjhTy+
pvKN8U9Ejk/niIs+633ED6NK3hFzDOoSgOj5q/q6lcJE8UicVPcMIPM53kT63KGu
0nW6m4yV1Z8H4a4wZwWV803TEEOJtEnCPzTE/4bhDHYAHBz1t+hg+FuQo127vKXo
2DJpbvYiMbR/QCslCNHrqpGfZuAkF18aWlaymLUmmkKg3qqnQ4NUkQqdlAY+b/Jn
yqiWWKiEeBPObP8pzmtxt95hhjHeriY/yThTv5UXvffXZ1PwrfCfhl2peAG3czaW
45Nf53KIspOawDhuwqtXSKpmIC/2oXzIdnVcmOf++2Q77loLvTngfVXHVVWk6mrc
vik9XiXn0c8qGbtvrrMBa9eMV83/ccNSJo7afoqjIFUIhLwspoZCN0PTYq5w/sA0
1bQNLQePWxxT7Emuj5b/puNo2Re9DxdS1O3tlL3IyuvkRzNTmopqUYCcIJn3dFwB
injtwwcmGFWOD/4OWS5Q8TPTzSZXBfzCElt0ng5TVa3tnm0aP1hZYSiZYO9z6IDB
ech1rdCBDxntlfy7AwvT7u+smn0bGokPZ6t+Q4YAQi7dccsBtJOxYGeegXmsaz2s
L/RrjcyGpyK0zb7f3xzCzTf1XOrtrFth7xQhReRz+RHzOzgM5lPM8tQO4/dR7ffp
r3gAjyT2rHXuWaBrD9n/kDkpqhUTBWs+X0vCM3JdEtQ4DDCGEbUgGCqjc4TwiaWT
2xwSF41KsQVZv96RdhW3w9A0CeZ0Cagh0lCDX+WGkGmDQ2uRNmdd/Vqt7ShyIkwl
Nrm/izHEnLtzTVbz0hQ2H4/9P9EmzEBqJbwcXagXQA1V3BoECochqUK2qf277PjV
LHKVFYLfLXxE2KyTue2bHEzXbJz7pwi76gYAGeSzfVqlMtIM9bvrREsOTl+f8aes
cEUJuUcE3mNU3eJVfrq1zFs6wU5wAeHEF2XYg+TXVEyhWsyvvRzh0gayiMWagF7i
g+Lhkk3YjRmrCxrT91ACCMmr4L/4AJLTmO4OTlNWvj8pMcBi/RtQNj2IAlNto1gM
Vak1JTcaWJk8KLuKzNbfYnwBT4UGtXS2lkwJwauTIpcXbqVZe4DUjiiKy5+sNY90
/TazlKFIuP3TV7rRNgr+cXD3/rF4f+tmfwY8uD/rNrdJj9TH7F5GHZxNlc3Wehsg
nWBqpK1wAObnsxq2FwXbE2tYB+Q37jLYTPAhB8rtUzHNpHJW2hoZOo/583mvliVG
rxGrkT7gygZhvYEHaOuQBUchR7GfzBlsXgfhPwIG5s0QXsYYrrqatilGQ/8m23Yp
MY5F2ZFHqmLJwQU0/4TbqcXNkfJulWuGluIJ7q4sLu+FrtPfPkEGH5HtC5qwucN0
fYeGtxGNZfuoKLflIRvjWABon7OWLFRLnWYVPFKBsYJwEy/nOFPpc1Z/k8OsqlMP
CfGhaYDjIlkDVvtdwkxODLjorqrmZR/i+YKHUSzMUfE6I89+siNqE+KfraQoIe4e
sfzlh+sMTZ05k1q9/w7p19zdK1Ytbi06BjQ7utYdWHG0TVI3aeCH0pE76y8PnAQY
kmwZ5esOxJjeNoEUTAReNJ2yi2MYTODU83MO8Q+jwzSyFl+4Dqw8CyahmGSo3W5U
ldyKpYsvvqxcNKtrverA4H8udR8CRMkijiO+dyKS0eea5ngYd09q6FM8lLeCSXs9
tHQMuuFkTxlUGwOud8T9ahrkgxmS8fqG8cmXLAPqgpgr0aCM31btAz64ZC9kKI4H
rQALDcxCnPPN8DMQ/oGEQYA7SbZ0dCH74+qy6PttdyNNLmO+c467bRm20fPFvOXI
mneVcww/XgcmKe+WY7IXYnoXwe5JbWlUFEG0q6w5535nzaWzGwAYRxNgHTLqB4dK
BSxZk8Yylzdj2NG98b90ajwEPhvtTEPfeRywmE2z1w4pI57iaOCHQUFawgnPxMqt
rfaFnUYnHBZPnv5nr0B7IgZRDDs5tYdpRL4uFhvuWsnxJRDOiRi2TKBPsNA/FnDk
XSTmzt7zJftQK9JL2/q/WqyeGKvnxNBpsaNDPYR7G3ssOuO4NLDd/7XnwTOtt2iK
9NlJdTGOMmCM80wpN2/SuizbpY0DedPaLZjTuEeMTWkvDMJXRvlO+gFLEttQxtj1
7LiwV9QxXhG3rrbfNA4QcMjueHdBrmsuXy/8FZMAmR+1Dbdwf5pRRrAYwYZBCfXk
bCkuoK7RnfXFZxb+ihO8NVS3PCC5qxqbMjtdaQXDMFiOwO0oDhJwAmarxTRFk0V0
yz0fdQWf/cKrbzyKsfMKS9qgFIWHyBuVYjYnNaGCz0BQ/eZxQNSTbu+5tsEGlc8u
6oBOb3jLP+6pSzFbi/Org8q6KarLlmriuwB2j48m/8Hgq97qSlU26sSJRmtrXjDo
OVzTrs3I2PZbVtBzqKXgqAmv8iiJoIfdJzN1lrFpTiXRAn0OjQZUL4cNp3f8zpAR
n3VlrK66BRZob+Hyx5e5bVlEgviy6TJPc3UlvU1VPdQpuofMB4NVREH4CaWZFqae
/CA21CcTR+q2qiDDBxoyQhAZ/W63ChBbWq7jIw3f20XBEiiXylzxBTkTzH958mFh
Z8aNr1ht2PvBape/5vCPAzKfFSPPWq/NlwDIDxREnALb2O0KS1wIbpkU9uGjtXYQ
j+mA4TeO1XFPfeZIgUvQ7OpFR2gTDAyqdngBSDw2Xo8hnBnT1TB3VL2EHpfcE0xp
Yfkl2+9YxsfX0b3dvV47yHNyjPHSr0P+hUSWy9IEwBaZly51Y9MUWsSYwMpDADFc
SP9bX95zT5QqURXTpax0WQDsGdH8npmFFYbMKBD2S5P5uzaJi/NDuZelaopkocWX
J+9HWng67c1H+idG29fVrZiNUcQmM2tGSxrWGYkLuty8lTZrCehjmwSonv39fJsz
LLu/Lyycy5JImhU+3/4QZQFsoK6QblRBXUgjjY/qZCn4SktiP8xvGjU05D7zBixp
CBwn1Rdf5Fc22TS1zLwbxrStryonW/Ijf6L9EchYO3Jv7JfRTW2/qhFJXTeqwaoP
rsxzvxR6E+5elDapWbcS025yZNePZ/8Qp2eW7iKFj61ry0oVgCQ+d6ExhYTRAwqG
QmhutFrraWM0F6OQawduYdEcuNcOHK3L57CxC2UUqDRZqIUQj8SpvaGoipRsjys+
vJzzcHHYrOrDFsWGL1//JniYlMdw/FOxW22Al9jqQaKe55/gHQCe0lp0U70gowAC
GHKW0OdDPEkZAcTlLpv3X0DJwP+LxwU1BIakna3EGMxdwz7FiqdaErlHv9zY2XvO
bIWazhj4GZpRmd8SpXRq2bl4Xnp4afzYsieCeUgjvlD/SCK/WVL4fep2cl+hNxPm
UvGZip+JZEFvQjz6QgPxQnqCVFoBPDuEs8cCGUOmP18OoIoQUeIs19z7rz4ajc88
EqgzU9qp0UgYMfP95FSAUqSuPyLMS/mcTZ7PN69Km4rJlZW0FnpkKfjrMnwQF0tD
YdLs069JCVhp6+TdVIDXp+kKBwITjKvpsgd8WxBPDoNxP3+hglqgEdvZN9MTkm9G
AGvimzJcSzrMRmhO5cftagNr68Z5tq8K85zJGOCkOCsGCmCbe4oLv28NlA5RGk3B
WTBPUtioBt24/WrANjJHagOg/B0W42RHx1hyh25zFNkHj5p/YnLC1xbUcgO2nDoh
uZSbwowVkUGPJgy+ExDocjnEx28HTeRgQi3s+GRFCt7BnrbJuCglmc2swB42mXqC
xefIHc/LJkzkjDswegC0VXsq341ukLsOkukwqC7JdbHLTUkMhbOGSNBpeJGXEbNR
AwRa/1KNS5LUJZU5UaEIMgm3OpkbfA/x3Z1jO1+c59HS+31w0lDjn4HhlH3apEbw
1kwr86MOdNnL8WfUwQ/hV5zQr8GN3hBBerEVhRvK9idbVv3bExMn0PS57EFCShDe
nN8LZJfyc3fC6bC6l/TvQt7qOoms8q/rGa44BaEW/ZIhzpP6vBQo2fvFfqA59ggZ
9rfOV6RUhCOGltzittstg+NUWe4tD7tiNOSRC0UT4AJlxFu91Tf8kGteMvJX+L+f
uwt64sI5P57PgG2MQQMXyaj2K3hDglAwZ8yjUOXzhAUmuIyLrQXhYzHaoFdeCsH9
q+yyUopxMe7HBM02Adh+Pgl9udTYlETN00mIKtCJsNIlvvEkdg6Abq6d2yAPB6Pr
TM+xqyIF7iB3QiK4LAJwqjDbC+QFvo9k5LWJzHfT2HXe1wEKhaQuZcU52XLUCcQO
F562q53CxGel3SyDvq0smldhStvkOehwaP7kA1uyMQgHeDCR0vTCaxplusMLMVgd
n2ueqUL56DYh3jqK6KJMyRTAVHh8sJkzcfxumoybq4xsqFD8MklIs8iIf/j725jW
7EDn/bY2aQk2plUh9ll4Uy4T3fDs1A5nzXDScK7qN1VoCgZZYlLfSKaoTfvbA2/d
TO8BABcqPkC1OBbKJJdJlg43Wft1/YR38Nr3jCk+mN3OB6DpPDeKu0xSqWzGJ3Ih
sCW3HFFlL65hgVzZkErZCf/BFVbUT2/lse3QB69sqxNKfPfck/he+5cf7Wq1FquK
UgjYbaOyztpiFR/SdlLXO4s8FfG2u7w2FRhtRTMscAQuZnx9aW11FByfQkNDg9gZ
TQm31kgL9F25FXVwdBtMozsFx3JWpYYQgz35zDU4l/Bb3BW7YE2o+HFXHasyEkFj
UlL7b6s6XvbejoteUGarOy+RjuHqBIEfq+sAW66CCVzds6wCPOzCx5+nVGbhO+Wj
VvnteFer8W6FdYDThAG56sZ9SyTOSPjfD7dECFyS6Q4RSstJWr5pLx8oMV39YimI
H6Pd9mpXOPFqEDNgL9PYMjhrGYYVsLx8PnkUnMmI/kDDgHl7Al3fdEEmqm/E/BQM
ygviQTgEYWP9qm9TDGaYmTSn6X7fvmRqXg0d/dt36rgxZGpjkom0slymkP+SWVVe
UxznbTuiJcGBfC/i+KgMUJGNJufZEbW0A0ut9FQcYemOio2iMjW2LwP3V2aRrAJL
l3TjaSEcd4y8uCYHBSAw4PZNeW2pNoFk53AQcmNj2VRwbCs/cKGFodvGYbl1ZXzx
I3UCN3ZGPW0biHDuL4misG0Y+8Hk7//fAojh15EzR++rZaomycRd9zq0fOdEfuUT
MxpCSIjCnr8YR7lxlX9BvfYVva+3JZ72dWasZopTSJOpFJzPD5sgzDD7kAfFA6bs
KEUV0/Tzjss25eFncayScDx0VVgNITlB7lYtvcWjQDs/Vm5644TOBc7E+zbyp05H
9wLakt/wKx4LiFPac3D4pretOT0ydh+P9F/dpccQXqs7Zs5iyeqJhstNidtQVqhr
DMMPMLaejmMEzFmfbldHDOBwP+l/8fkFsgeWnlc1IElsxobj813Bx7JD2piv1icb
QMOuLX9ilWD9zzxVDgwMIsJSqqTvqFn5W9GU36OfG1Yj4u/O49AslH6LNwPILLEU
HyWHnDiUkkz2T2cIQvr1Am7ZvsFha/b+BJgGBRxaUwYnD3kEVKk4mp6vAwqO8XqV
Ba7A831j5nQztMPa/7CgtXF4pnrkUN8Annoa0+09ExJcKvQYYYMFg/CHnZtjK9xL
JYtCV5V9k3i1TFX87fzp+oN/cr0u4R1aRsVyHn8zePSquXPumsIFaD2peVP6AbPY
o1XItH8xeKTAMLYAN4OrcU+YBKLNKXNarv3ybVb0PfAV+O82rmqxa+xSYTH25TCD
y49A5hsLRsepW3dMFBC2Zw0KM+7fCFMUOa8QD2GXSnAOj9bN3lMzJzFS9A59OnOk
vZXd+E1ajr/KHVaL1dktafK05LOgzT5pWnRv7dfCKyVXO/O6aJSZmIHeHj99eb/b
Ir8T0rzkfG7Nsi7SofFs+a9TUqY+aoqkilrZAxInsJKz6Du1PufYP4W/nTFeThIg
QQyYbo04FEy0SJH3beSB44nyXLQDyPRC907iS2cpYAcXdQnia6ETFx8YAxvcB9u7
A7/JRYitfoNmUZZ4AiuQOv6j+j875zZzH+NPneiMh+rfVQE1xR2T1tPpTLmMWj3b
4YfulXP2UEy4VPccgLzD9+vPhC01/ksw5tiYoq3yy2wU5BRGdxLfdYU6PGK5ZNn7
sfmgz7YKX0FON/xVu/U+uiwJ0LGSMqqMI0s0ffueI/20UN9LjJvixZJdew6T2PL2
HMYUz15c7+secPJ2XwGBF+NmSTK7UMtiaVPDkM7ZROZCMYx1JR1Yvf5Ihl+c0BAf
kMyYE6cttLOJECEZLFS+AQ0BV7AZQdIPV0RkFP9USIddN/0fE8S0wbRQpEI0e61o
EpbVlp30/N4dMhZ891CvaH73dGqjdLYoTB7WBTvIKUP12OnnD+2DHbv3jjxh+kCL
sC0ch6Bys3hjGHJZAmGiQ3MI48iSXOsr9n/RRgsg2RwZIf73HZB9L6gDI+kukui/
gC4WQWNbTEGVXKitR1IaEdV9Zm/lkd94ywXuo4Vv7+vDzEM9l90SV/qthX9veWyN
Trc8TtFv+h0EwdkS4W052XYHJUWmFWrxPpRenCx6olqdmb8nAiI+iNE9XUIROzma
1Em9cZfMBVH2cHs1bBhUxDTq0M7V0ywPlVR4H0WMfA0PFXPq82KVQrUdx6VpYiAu
wLnnqbcijeAqXlKOxMPsq6iThZIN308EaNiVRDDpKsPK9Bkih5H5mQXV/75ZrMs0
zCyGgyXrUR8wxmfz+I2TrL5QBZM81bNAKdVundmVVyCS4sTnF+JpwnUWtKhkgLx0
Wv6svLUGvKWjtAkkLU53LeO/R97O2vsgWxuSsuKNA0VlvZuAGdERc0be7btnWiT7
5GIU60hrq1dmlD0cS/YcjXMAmmlc5iC3qKVvwDF7JDRKXWTXZJrwJ7/tS6qgsi3b
qJBZ8vI7xYZAtK7rFjpl8S3PwS74S8T8FN2CUwkvPSfjclqQxudtF2aWxig1cLRo
po7LMKLDmKjy5T2xewkPdXHjUR1nXxJxOHGrk0M42O7Cs2VMnTb43XIKzJyFPcjq
pBTFQycZs/mCSwfku85VVITJ4oOOhbEH2Y8f7FtTLqA5iwuojJH5MgFzohf9RrJc
oJ5lzrhVevAdPKzhIr3UtGYjT5GnA2wQuWyMVoWgW5RQlmxrw5Bg9J0rpdO0zSYY
zO3sJc5vsZlFJzeb6crKCSy608mJhB1VsEihKWG+LkKZgbq95cjKFUOE9wAF8up/
Hri1GcdPbI3oQWMjON/hc4lw1wAtHbkpZAEKZcufdysO8tBB/4uEdicMP9KwT2Bq
NPp55gxnL+laPIXrjdechVwz1t8Qoa6D9BfViFl3z6Pz7uQrq3ERPl2Gf+rFvboB
ulIALBJ9Ciz01655POISQKhuS/Pzer/WC47wt5/QMI+7sXVL73mBdOIoVBUbijV8
DlPuI9zdQsF9byNkZLB4X6UcqOF8sVgLJ4rl8GfJAfF4XLzFukrVP1N8n7gUyoLT
lCzVv4ImHuuiMPI5kNtcFt8FuXbnzedplb9p60kVCzV5AtMjteGaGeeCei+6Opyr
nvdisRfBspO5kZu1W8E9HSJd0MBrQ9Zfs1xzq7MCRTC+fv1YwzZW/iL5WzFjUvAw
q9Tj/sLYQCRHkNRjtXf5O3EBdGN64krxv3AB6yHphx/iNqqnRoLTeeIjjWo93VbS
wyLcoOdD1CApBNzlZwBvniqkQv4s4OG3lZu6chyF9bpGJoatgBWhxVQ9pflQ34/+
dvSA1UiWbGesUMrlBaN3Yh26WpxSWIvuOfyzd0pVRa054uclksx8MX00NquBGmPg
Nl4tyn/WgOTfwm/m/SrwubfPA36l3IdX9m7RUcxqkNH77OXaBacyWyJBDpduiqYW
w/4e9YPh+NyU6xZTGi0wEuacMQYJuFgYlEGgO/hD8qARbbDwTTQHeWRmOskNhwoL
jXIBNr6qpEifh/iISkdaTpYtuvJK6ei5dyV1jEFSY+g5nCcxfRf0ZsyL1U6pdg6H
VUBytYv0TQkxKeLdR8XpGAKqrkJHSYmyPUQ6xV8mAzrzDmDmZfM/iCf+VBYjc6Ur
3M5T2DmxfSY9rx3252oBYDYF6Yd3u89wt96qi/In+yoJiLzozBV1oiRi+3fjQaBW
OpnJNdvU+lc+bT0DylmkeFNkCZuE+ZDHE1WT23xEj57HEmXn8ePvYKiCbmgA8l6L
bONEiylW8m3pU/17UHDPssYckLytpEPzR8ixiUmjz7aRWYM6IqhhNFhqE08eZX1U
vZ+fdZg6UmDPUDGSgbkdXIANXNo2ujm26Kw3dBBPcDcIxbfHvF2phrdnQzAEIW+7
NTDfZaduVO2+4XEiVY3/dG9TtOTxRJoMy1iZwcXEYC8KP6v+peuGSU/iwLILhlqg
M84qDnck+1iCif+2oZoP3bYhgmyzEIDfu3yExS+knkzty4HJRPMhAnG+VmWzc5nE
Iqc6UpLKygMydTiBTUGQirpnW/svdd5JiA5Xo945EEWVuIJQZIMWY6UyIbEatg/X
OBC/FoUHdnFm5MYG83IqO5tA9Yfrm9KEbqiSnYrmoHscnbOf+N8kCz9EqxbEq03U
b+mvNqJ6Jgb+4JHYxMR1W32HHnH9IJIRdUV4hZNOC76FkUyF00u9UbGg2qGUan58
ouhNmYcio/gvulxQHhxoEu6VPlGvymOZeOyIp6LewdnpJVRKfIiVJTATCOvDWK5W
KnD1a5n9VX55gk+QCI7pX83uU5xb1gHK3MdaW/FGL50FO4UI8+MqVZH8nEZnl0IO
UbrA3jrrJE3Q6mNbtmeiPum/Nu5H6Vv4eeNkUCHlD76uaL+yB8yRinQCKp5u1d/5
vDcD/2G19OwPvdFYXqFaFm5qwMOzd2QSq/TfJgY40kcolKEmOWYQIFVxo8IIDqQ+
IC50G2kQfPWabGxUFwuC13lGu/dNyPNTSEw3kvTimLHDfh0XcPMQ9CAS2jOoy7vR
QVWSEg7D+XkbKBg7TAEstrz/qeQXefbfnzvBR8//Ndb/WNOodb/xEQRBEvtCzhfv
oBHNj/e58nyUH/MJh6xN7TRCqt3s8UJHnkqaFlwOADs8SFAxBbMnHa/qraxkH18I
mdj5jfw713hQRw/ZbRvbTtLJugkAoYkj5PHWFmkxyPDByVEQ52MFOs8fNgC5vdu4
H/sPpHhna/g/MwiEvPZn5F/9NFGAUBYUkzWx8xLxU3YFWLf8S4TwMIk6ijd6HLKJ
xnkw5gx+ej4wuUIjrtBVKtUx/w4u1McW01zEg77ulIF/zShm8ZCixyi9MVjlImcZ
o+hZioq9+i65rZ/swyooSKsNxmGBDW/qtvfgqjbHzdTvEC0CcwvyWxpevYWh9Klb
mOCxK0BWN1PgyJm6aTDKTgpKgfTW8VdRT5LNjy3VvlGrZcflZWXl2oapIYcosN5N
mF4UKbsS7cQSNPrprjlyEkEho1SFzkDlC1iYC4UbbmNdIDJnxV+Ll95UvoQnGTH5
iiAHC+PxuD205rwNFA6vWro4r+RWzvwkIxOqdnIBHenvmMQ9TG0im3npJufdTw1x
2L+jeQR+EZPFOrk4Ly8KEpdVSLmTHhCHRPe8VPMz6C6OJJwA6BjIVb4PIjpCxxxs
X0C6Od7UnRWvtZsiUL2yx1GTQYHytQkpoLGqJj+LSHNWCilB5SiHbi0cm3mBKcN+
FVkDsSWUObb0/Qpqk7E7YbgSPBV3wEUMEeha2LWgCZhgYSm7+Q4AHqyCZangunpk
bJNME5b0c3soc0HoAGKGlSGo+wrmadOBkFNT/0RIX7ooF9MsKd0/NIZ0D/3UY/uw
5O2u1q6fZiAsygnVvRTN25e9t83r1nLQ9JXicpAtHWmMzfoKZ5Hp/AI12Drkj8lf
nFKQ5rDNjwFjh1XsUHijrF6dF9Umy2rBTSn6e5h6prugPfYNq/R5pLHOu66Os3b+
uy8WboIHJ/lApHSUqzXW/l0ITtcQPVvNyZ9jb2HPZ9Dj7JpWXrKIM/t5SUCNctNK
xeiTSMqRpKtcgmMYnzpSDGejIXw8OBmxEoV4v7abNfmtTBRe3cXJzUCNlEUutb3M
BaZd03LLjhP4SF09gQT+x7edZzJ01Mgtwcz1RUDM561qmGZNIFjhciorrnJt181i
R7nVOwPil+cNVm5FHiEbyXlZriZyBSI4b4meYWIudt2N7Xp/3bINMgTEKLKCOp7F
s1eX9QiNRZtDUjqgXsvXRekJVylW+aOvGYaTNTrZ2XS0itvKM2pKQjBEx8MIcXeE
pilvmAR4JP1Jt/5kZVj2GEAuLHehryC+5LCsk21w8XFKX/jLVaeU7CrqtSIxfF5Z
5M6zhDLy7ijRqQuGFvBQUOVBqIpzFzfT/i4ARY1YXuZ3N0mNjIGKM5GCzRdbhqkc
pACgkzv851XKImMYgjnpT75/Y4VgKpEJbuDciYX01oLwuBeurbKaCsbg3OCuSR1i
/faZABMLhF64aUyUKCsVCTBggBYWbkzB6Ha0YGsrSQv5FK/lpl/RJzwgKUH2f3Xn
u45xmmWEb/+YBcYc2uEWaQ4goXMKIOvbIHAsPMXoCjfASf/M+1SzUm/qcjsdFKC8
TZFwfY9alo5NOdsqWGT3WHHJ/1vyM4AqPmQjB8+HNDUjrvPu8TmWsBiKERM34qLA
rYQIWocP+M8OcsG/CSde+JEErOFePl28UPWwoiVVjN+2JrUQsbbkc636BTJPV8ZR
ja6ZQ0mWhgKdw2ILpvq5aC7xG+pSKaGDV0EcQxeNQVZhNGJvPyejNGLCcQ4TQL/C
FFiRV4AFxwDexKxlknHedEGV4ahY1ajZSncJb3ACeOkATeBXkIuU1LFsVL6KIQEj
bsdBx3OM5VMN31N2CqpCE5gm0OoNG5AZHZmjRnXUDVsPb7QxBAl/rTthhKJhxQn+
zpwxpvaWRNjCqMk1WsK/A/MRPsCOn3wHHXVIJeEmF5TDzBZqFg7H2pCk4MsrLNLR
bsTC5iBlVw1Rs81l2li3xCSaKLD4dGbo5zaERxMfWyuNMbS4DWzUuUSgFkTwJ+20
1KsyR4wCJcbvlfPDUjdfd5d1rwVdPI6SvDg+r8f4YyIiUw7by+FCxz7whT8dXBtT
YbV9cfol8PFVsvrCebnQdHqi8DUieJEzwvQEqqPrvepsu0leTfqadcQap0iw7b/j
K7iq/Px3SB4kHJqGS11TO4OXSCUWexysf+QuyXSZMu5FeDhLGQDQOVeUwA9BBAmQ
m9TE2xAiPaAmkB+axqxaislUPnbw7LwopJrcOdQxRcxvNXJe8/5GTthH85SGgYs5
bK94eYL688tyJ0qQKVzy4S3Huec/MO89ZG4hwgkKFUUZq6ReCdQreCu2Sp1NEWeC
LfqPNZo+Gi1jrLrD9akmf7VPmFCtJFh0SS+YvCehaxY5qYzGBhaW44kRypVSFdEj
VU5HLwWAnzW33MIPjZp37Hk5IqN8Sv5SITW6XQIjw4jg7ANk2aSgNhlndZaX6ojx
842ynTSXQ95VAyUYSz/PwuO1mSLUZjn415Tnf1nDYAivm0limlRsKM5P9c/L3Lik
brUVouuKjoOnHGwKTtAMNm1QcdxLbWykYRhPj9S4oTMEqup5sjBoisVthaPleRbs
juVg+L6E0BHXmLv4RhHdL0Cocd3o0npWPdpMmkJyG0gp0jQ125920av+yQHVXxSM
jkOQyOe3505mZb7p67/i6C4+TfKrdkORKarskvuvCIcYbM7MshNm/blO+f8QdXlC
K32cQADLebWSrKh5kALuUlPyibC1AdkhT2xFtBx4ORAIRKEqWd6TXLX+a+yXcJQh
EuVQs/hpOoOSjRcFBkjLiE5LUYnYdSXhD0HOE9d1EvPqJTbJ2tH19U9DbFMbeERx
XNBfyXPm/s/yJviy+Q1UT9tTyuZZCozuG/xbPHukhW1l4aUEioEdkIq0WybtHRUg
5wekvmGZpkGY++qFBzVEaC5/+rgGMB5NzsF8Y2AcnSXGRkJMypYGqFH+zyVp/Y3f
MWQR6KSA1IM2fqiZ+/oResBbxmlvicmEQeUpkvQzBSUVbwl7xXUlUGlAbuUSlnXy
I9juujx4U/Q5p0/yyYEVK2iCvJP+dds+ThH9fIWw/LKMVfb03aiuBXvGhFSxzUNb
httv4hyuPsfRhWOLj7YM3nOfg3vO5bVOK4oUCnkAUjQfqwtB/+teou+X3cwhoR4S
qtQ5I0NBlEWf/N6wQiqLr/bnE9W1NzVQOzTUt0q6T76sIa1VMjioSIYol0kn8Rw0
NbziTgtq8rTq8RyFGVUuSz3mGx/NL8CqNEbfaf1ZvP/h+jR8AwVsZxUTHxDmqoER
IEXcRZnSvdaarDkniZZZmFUsXedWfWwaS5BepJI/7Jv7PLfreSRbkkHkhh1oo8Uq
MM2b1p92rjWysAyflrUT68p/BoXq2KMHrRadobICf6Frp3sanIGI5dTP1mjhutny
peG9yzC/cGQBVN0/C/Wm94ileYDI21+XN1fZxDAUxDX/9Pc50Fode/rhXGsn/tME
N0ogn0uCgsXuDrKB8UDDzsoMAAsCrbFAQP2Elyif+GAwFodc9TZUaFOB4ryaNaoN
v5K1RfIKZPW+TGxuyzNli36P4xYMnwLA1nWOxk2sD9IpqaJU6D5HHg8CHicfmZ4V
caBciWjjeLZIzAa2bcyvHAVU6cQM+Qf58kcU6OZaphL98bKFi0h0TiDJmWqbhukp
q54v0eVL7cXv4t1m+PVCu7jLvB7tc56P7EdVhhv/+FOW65UlDqY27FaJt6EVqu8m
uOyeb76oBxjXo6IpaEfDnfGRz1Vq+gg4FuAvi0o4M5TRWtiA6IFT7Ko5KLexY2Pi
d3GcgJhZUVsb7MMhxihqovr41657dMqAMyIMXYfbOd2k5f66e3yatrTxCURU6+PU
xDdNtnubIhh9uhDQnx9bWemDjaTWEDdyQ7sM3kAh03TmfmlYo+cy/BRR4xXPoAoq
w6aW3q/5pMlHDQd08ueDp9J6c9tbI8Iub28XVyLyNIKtCq6ehzv4NANv+lNn/iT0
p5Jvoqw51/TO0jgwJgUWzZnHTdZMirlqEY1UBMLqSc5ZePzbZyLBECIb2Hei95jz
RgLCnmRMn7FBACgAbJiWp6WDxWdt0+tgLXdDRnDSYstO4XfFo/67Vzme1ndCE3LL
P5D838Z+grj5cM6qbOOdVGZYeJw8x+7x5BCc0e6/owrME0ET+8jotT6kjpl7wjMW
6OYRx6EnthrjMFSnQTb/Z/hIjtXKLGQiUU6cnD4qRGDD/C52UFHu17mLZwjf/QL5
mXJDu1S2haVMwlKJSH/uW13zZQAILj/oFS7ZhBniTnNirDKFbnx9v2uhZ87Rv0pp
dir39O+X2sYbkliywCXjThxZ/TjKbebNU7ROfsH0boc1KVbudaKkT1Hnd3pAZWND
dd9US54kKEtn2jYbi/qpmhJwVbthg5SjiIf7V8Nmmm4wjBC6MrZPpR8UIy6r1BRh
3noCch6nU/qv5453eUHLJYKIcacYJFPAX3qryi2WmN9Xp5K29M58ZBMRtEH7Qe1J
oAnX89bmuPZ0vf4cUXJVnuuAfgYT7Z3sm3YNztwIv6rSXe7795VFu6R1G1Wo8xBq
UMihnKRdw5e3dB8i//NyGC8ThdXva6DU4Tn8oDBznhwzXH7zktitExQkwymgLTgq
tsF27SDQBosTAF6+xUKfFqvbK6JjXKHtypaj9+5IFWtsrRNtNlAsn53rtTO/wRvZ
WLDNttAEX7d4MOSCjQlhaZzW2qM6W5P8DRBvPmD/vfnzlWwjl3f4mEljjDufMWzp
YigJhqjcnPhJNesTCm1uqTg0HKtaaC06Z3jyWlBsdqop/WwUp5SkeOMYHRKFbqSY
0JnU4JKIDJKRYRkNXgp8d6B+XkPrjkz2zUlV4+YdN9uII5ufm6FCSUPbiQeANvvY
2LMOaCi/K7vJFpWayHtiw+dWlJAQ3/+FhYLMxXqM0T74uJ1cMI2sy/vDifdYBEf0
/q4wl0C7aBKdRD5RyHzn73ePS7f1Uj9e0hyQG6+DCuDkbC5jsYe0+QBD0QWECsF9
ebHP0/EjL8yGywDf60NLKDvzZP2uIx1xGLffVPU9Yoq+8aO/tzPVI6YOQz0Pw+hU
sj/YTB5sfzdZbeSBSACKobs6munIsIHXyyEUbzYgRSfbGbiotsgI+f+sMV9qdKW6
u1juKWuWKqAyQEzilNCCCpcNFmqTiWvzq/ED/yP2sl0h+qz2W+l/GMPJsUqHvLzb
RXrl1qeeYT/XWW8zYekR9ZYKgUuydM984ucbn8bJsIMO9+5OTVLqRoTsWXK/P6A4
kZ4SmLPLL5a+KUzqhiEu/v7QT4PD+c0hJJB2oVt+x0WrJLUE0ukqC0lBwwhIGXLY
4aDoZwYLw5SCK+lCvVKfUk+k+ylMC0Awqxif3nXEkyCF6SHjrg1msIUqUIvwKxdh
UREe+Y8QBP7ii/uGW5Oo3U0Pmq0UDKyz6m+wTm4vZK6RCrJYiFPGWFJQmo0oNmCk
iDtuCDAHc372L2e+/hOoa0notaCuBn//UWxYndhlefNHuYBRhgWXTkgwtd5JSz0D
EeuxZG5MlxSywlG8RIf2fH68sczuxd59jIAPHU6RXaCsGkVFDGCyjIRNm4AHGXCO
5hmwX5jJI0nZHlx7oqcq6cIdJ8OggaPCXaT+suUkMO5NAG52XDbo/CCwV3gpiSvh
FtSbp+dBstnsf1t0U+qvBSz/8/7pKJdByzZwTS/q84jlIb1Sigdl1HCk8fDtdxwN
JOtb6t2TxX5PABhXypzeydc9TAF96UypL+6hxWbVm8CDgUKjFG1F9FteyvaCA8ba
Hk0+6tuYTLZELMtqFFa068BKJIqiezZGA9XlO92zdAZna6xEWmbE61sVp8ZCJLm/
Dy93iCuHjFEpYo81CmbsxGdRD1Dct4crW3owrIiDiaynOD5mnOW8KzsypfEaPAws
iQqnpnFm3mWPr79p1WH3qVtI/tgu3Njt5kprlhaSjEpBpIPuk6OQM/HBJlI6Ya9/
8rCS4GCIzpPTF+CvkOnxagnpnyynpmn5USKl+OPgjBULO0VqZuowZe9Dpu3ylgy2
XdPdfr+44rO13EGDI0JdU5xDpBdzYV1BxBdcXAEqn/D68+8YgG+AdmYveN0Yzr9m
N2XZCMk6CrfR3R1uE853JOxJDmS2oLdmmA//e4ITv/OrpFkI8FLd1/KTwNS0kItq
nVjSKIC6WbldoN1stdBENhx8nVchpqrN6PjGSPbatZCBlsE3XQ4ByynY2PvwCq5O
nqE+eKmHaZ+5u7mfWIk8jwg3QiZMiID4W1iZW4Zx76HEIQbL2Ym3YbIarY38e6lf
BfjqrqodVHHlQb+0YKCOl+YhcOrFOufYc3u3DYS4aHVhjXLGoQQ2kf+B2lbxGYpO
EEhVGzU3sh1qNASqyHBm+qZ+4AUFv1dQWCQqpYoBgeWV1AqUMTClJkupowdPcNsS
Wgkf0eX/5z5Tri0zFpqhLaIETMu0Z7u3Mp5LrvP35xuIup6YN3xd3al8Jod7oeBq
EBOBNjN3eBsPH5KeBrDXUZiGf4U88t1prHY7hrFVoeXvS2wbLbjVJXRDvw62X7Gr
XXcsf950f9W/Som5bHTQaji95dT41S1LuxYaVHRQPKv7NPRyhhNqiFT/HlCZl/fC
v6t5ITMOy2NcYfM0e/igYQSe0U1Rkd4bYJ5fiNU7weVyd7ZflqAIZmSSjgcYvthv
2CSamipwTD94Wemsg5x/ZCwLjO/AowrGOxz7x5gQMsmc3wXf0HdZ53Qef7eIWHhK
ZyJn/EE7WAH/zipaw/2IdIGaw6S7v/97FaQeF1WUsPSuXfGUGX2QWLO1hoI7RnH+
Ra2BiKxmKC0HJt2QphBmyBaeFQ57u71KbFdT4bcPQkCLRdHX5rW8Ef7i1egLTH35
HZ1wJqyvj6DtBzPumFRSC3101YvD3Fg1oHvuKUowdL/QWD8Qy8bSfk+C6yAjcAa3
3hO9cV0N2HBFVgtH1Tn7EH4iBULSofXR3lebYV1a6IV7cCcE1A4OXJPRxtw8/js2
yRoeFLhOiPUkXhepSHFZ43cgJ1Zg6Hq/g/SEkKFBrYiPNfs6D3Nq0wqh+GTs68+X
tICNfSgTQkPf1yaFxJBtb4g6SA9bVxRfbSKWtrGXiGUnUAp4WM3kPwCmvVIUgIWC
XM2tvCkfEU2s3iQgukUlbBq4oTsElCKBZ6QWkLEx5Qg9d1tnkR+s5a3TLDGAob+b
tCKGY6t9thrrKaTTYLOp/LJbUAR7tVWgwCghKYEhE511/UtpW84aWO1DWOsPuoke
oFUA1A+uTuoq4TBrlxFiW8YEliCS3THMW0HzqbzWFVjsmcgbUE79fYe3doqhVBIE
SSHNjLcWIqI8ehEhBP61u05gugWQT4NXqTf8uccqPCdsXMJXCMcIGr/lowESU4vo
r+KSPDPMV8fN+IBu/6EhdZ6MGxE7UIHBC2C8F6idedVSP3LZCVpjB9n9+bdtBXKA
9wwpD44M07Fb9gqW04QRVgOiijTnuxaLxeWOzI9CZ473CRsuB8CG3eK4jWkm7dqs
gJU7eiXpYVlWra2tUOptjSlLQ8WEX5Ri9yoyOMYKudp55FuevfPIgfmMvnxC0nTO
7ay9AXUob44tD9Yr3iMFBCVAJiAY86gAF0Zn8wW3kYwOw/FNklfxjU7mJWZcJlQi
SBAsn3CBR3Fmr7/z5p+CkLKYWIhrvv3WvYG9m1TEbd/N2ThiNyTIIpqoNY2EXUOx
nvxo5qOxA7CupRnTfXiKvxQZaRyx+AfFItzoMpUbU7wko8R4tDL1nu/wFkYshWhg
a3uX1Uo9I/h2A1vJu9EAjzvR4iwDcuc1bpnv3rcUUq461cfnYyLhgMa5Jff4wl0d
M4IxFgfjoB2Q+rz1a6uR2Bnbf5Hvg1SMBqHR2wkWc7dyDDFjSvGXLOc5MIWRLxlP
bcF8M03OQMwOQxhd8tete6Zia9Z++uh2el/gzlW/h1uVwt4tLL6s8EdmL82vh1cZ
TYddqcozxk09KyIYiL9yR1te8PUnnW4Du9dlQ3EriuNt+2fklCJR4hjUInFuZfnm
EahcXoHUq22cjnmAZi7LOxcXibPE1G59X7RI00C+nNb6jeKV8631W+bVEwY6goCw
yQ1tsfzMPQsuc/LDYOwjrwMJ/iPYlbxlYZu0YO2P+y0WT7QPJqeanH57M0xZAz+2
LV2Q1uH9US24LJfElArvqm30G4SrGFKAjBJyCYpm07x0/oU7cKn1elc4tZJ69JAy
Fk8aVjYLink7B5o5yKhAo5Gb40YEogNHhbFv9edbLPbsojOzuGoZ2fc7K1vel7sK
qHhpcep2R78Yknso8G5XZVKmaZjV58hs9HJaRZ7Jdhe//cMZUDk9+5SN38ZnmkLe
RwjJ+iIfzKqtC+c3ISVspT3WKrYMJ77tq25pps5PlFlzoajhwNhThM1gFZGG9RVo
TJMb0U9W7t6+5Anu26w8hiJzuIJtXr99SxbtJrz/JtmPCDUGes0G41aOkms/0bNS
KU66RzHb5PD5HN/JM6i7RQlIc2HBgPcR1xrsKj3TUvRs+kNLx6LU2zd6uGMxHkS/
knyxhyQ8CHh5Fm7+9A+HfMr5sYjXOxHccmDRmxW4qYy2ZwPAT/24V2s1v8K+3ajs
C/HrPzpq7fnv4+b79earu70h01qmQRrS2u2Ev/tELGMMrtZH1pZt4HcA7q1vD5Qm
SiqF9/0aGnwFoEFqLLBLJJjCEcueB9Qm1mzXMMGUH//tRNMpm5xjE9+oVUbf1pcV
EmNtN+r57gX+6HWgYxT3z1KBppMh13EziLpYxDbHfm0Yk4aXuqiF8HiaTRvaSjCL
ep5q/pVR/4Q/wiIw09hSDmt664XIhtvAh47q4p6pTVx3PptoQ8VOq5Amo7Ov+QTq
cpVxvDkX6cii72duG+kjd1Ye4w8LXZQ8miCx5Hs8f5swqTZK12Jm9KOMswrVdzSl
uPUJKZm7W+jVRZnRAYFhL092nrX7oZVEjcca1NIE/TD3Fvk3uNWepFm5lr/Wwhaj
zPPoC+7mnJcPdzJiiRBdlpRLmhPb2Q/3Y5X2Uo4YkQGfWTXUNbS0aya8ixJvzjkR
f0V2vvBMo/lwWxXlYuzPsy+7Vo2mshsZLCQEa/gEJGbmECR4C3KC3WwbKABBvHGm
AfN76T4vVA21y53gLLiTMy531vKEsTbt7gL2xAqw8ZGbGchyJhoARwEi4h/MJbuM
DBLwjwG7SVTT8SB0ZHPm8FmCg+b/HGZXIY8D5c67bMEJkpPLYSQYqkxVC8v6hnad
PewuOTD09EGdfFVE4py/uCGD7Y1jlyC520wMui/IR6dKsC1igt76G7kfwWpScdCq
Z7jIHqzKqOhylV83j9DUKdvY+rsCSA4+gKCmVhDeRkYUEe8dnKgCJM71TSxDb5ke
3K433MyRKgPPviwg8FpitS+9kL0h6hCp0vuBgUtKGYe+4OrNV3t8dpAx/0eTL92m
STOKALabi9TW8Ki/RarI/B+8jyNGZJbw6bfLvo0b2AJnGOzOtRvIqBVZN32cez9w
pawvoIye1h+XTAWqmbDugQnkjXJXmG4EwFDAwmEosaZOj/pc/Oy5Idl+iQMRUmqA
HAyUaKRWoZjCAbB8HdTwtH3cNcX0Gh1fQFtw6P6ICJUaYekl7FNd7QdIBMVW6NFt
JFWNchxiFLt1/cAZlXOQu9aJhMKuXTXAjyAxkF1Q+bxJKMS3ck4pKgcuc05HJBuw
QFrBzJhkwof/UNuFLDLCckJ0AYB8vsDjz2+01ZmlVp+WCVFpt6tMZuBRQdgEyJ5r
Y/1YgO4of8604ap63dipqxSUujf28j0DEWYu8w7svk9Hf06zZHFXgBNHfrUkEVIR
MUnviux42RnXEpSSfK9HBjvfbGKTpM8wVy1GcLsne3cUobHN7f69Y+VCZEMwjmUF
YirVfiqGqElFTdW+g9TNqqUtSOQ7hniP2d7rw9hcksKXUd5ZnrbGECjf+uF3sEsG
Nwc237uRN57rL5VQ4QpJq7hO30duT7H/OC99r7ich5wlXbSGuReYAZnd6vUNGReK
gOoLrmaEikwMwbxfr+XCdXCkal98dJi1p4m90lDBQFdb3IfVd32Knp/TutLYci2J
u7Flrr96ql5O4nVo2SqeMZFTphMwVb8cV2s0Iv5L4uY+PWg4mmMiXLOOjA5foXw2
Udca+G4y4WGYoLdCKm++9VjzoX6uK8icqRRo4aej3rk9gXMdqZAv8fKACx/hWgOE
W3739Vv0+cxT77VWxwiGZbBEALUaS2RH45ZJ2aHA1lQIjaOH2CKohb/ulvcJj/ov
GZzyx/0XkMScmBLltQFkAkBtkC3+Bswy/cO8+7Ge/+TXPQNNKls+yl5cbN2V45Sz
VvirUqNgM8gofKJLqRsz2bDaeAZJ+x6oY32CKoPUrPx0VNpjqTphbRVZ4oVlCnUS
bMR2c0mku6LQk2J86yZ6emOjM5S0p8jfEOj2nUQIQfV27X533JXc3lnTPTEOCVvP
QkzAu0Pxw0/xeXRtgcoZZBcTAhMfgCNG/YXtoI7y92qIMHHYcxbovxp3Jyj+6yNE
t7N0hcLyjymCuxO3/JS4H/3UO6643hEIg0c4PCyjuQ06pvdSM9f150QZ1A86Qcb6
5E9Q0KsUgNGCTlPxZV1GKcHgGq6tQgxNKo2/7uk94odEm/nKiBWG7DyhiOtVCN9e
XkMUvEeRnuX+lVCqq7qag9HTx1wMd3PGuFBqtwBAFBuMJjQuP97Tbm5HsXWxMxkP
wuYUim4cRDZlQ03Adnfuk3g5qAWCK/VVZqVeHdKfn5F1TbfXK2pFccn5pdlqR8e+
fecQtyImnZYr2Wx0nfcl9e2O0EIcrX/u0cOcZILT4ZHFUhGHZ/oyC756eA9qiKsH
Jht+wvLwoSthitkEMSIYBzEuQdnQYhiKY2xqzj1xXjT07+TuW1F4JYQiEQbRIBZP
9Mo8trvRfBrqMqpXTKr9cnNVUcEkPm0Lzq+t579WOsLL91+jiEge+4wtYVKfDb0d
/1ozrko0X/BxO0PIr8HAPcK8QEgzqSBMyC2VFJ73bkoB5IB603zXaog7sGmStzxo
9X8VSSRyxrt56OvTsfQxQv+othucNwIATDTk393r7N1bRY+AUmyVH+UBxKcuob+Q
yEWDy3Jm8Y03tRPY9SdVICW7ZYocEba5c0T9mU8ou6OgmdtGAI32JxZaAAyB5SH/
SanijrcZOxLWmGXgnZXkwbGKVpAjoFtL6TuwZp+DRnku51VYfUhl2ewZBoMJ7xgG
phLWjY5ezA5KIpGzR+LXG6CXP+ATwvZt61aO8WxID6shdxDY/yW9iqMJLIKZtzuH
LPOY3q1Js6qvVBHb5AOnSL5+Da7DYbqXqr445HfKneBqGAb1nSX/KOS8T8yK9YAn
EKQoVRRHeAovzCoa2wFXNZ7zT9VkOkIPpS5ivfz5TrYTs82AKrIs6BP0I3D/xmXq
PmVDLKkFt57oIhqq1QD0rHXqQX4Ywe7GGqn4Q8VwMgZpYzx5lDSROBOu1fM556fs
8uOIe8CZo0cbcb4jFXHxKeVF6iJ3Mchlk2k03BV1JVrVVx1pg6Szbsyoxsn1NEro
lFybAinXZ35PdKjxCfFraD2YiUE6xETv5XkGOsV2+9dPIraRKCRfPJ+lEFTwfMB8
lJNDXvLygJV143z6wgOD5zdTe4XgVv+YRMF4XqwQVgdr7pKl3r2j/PA1aTa7bznp
eHySD0qt7ztRhLGEn58wZ04Rd9WEhDFqDtk5f1A0qPJvIpB+YYp6dEKJyrU6eTAv
4BrtlulHCpAErq2L/qNaaPgYMOzWA/v7vHJ+Ae960y0frTzlMOKIAnWcpevIyXVq
sqPqjto3RnWWxVDM0viMMDOnbMr8gtlAwTzWM6EilZDRSWQ3QRjlbRZvmRiL/C3a
mF4VRGF/3aOtsN/pwb+X7mR5vaaLycB5/o4TN5oFwgsuW09efUWxIStSZOK/4UVk
Ng8usiE8bGkFiHh1oHtXMT8aL7KaDPdIRWTne2HboPt9UEtblfbv12CdrpGT+Agh
hZn0fLNxz9V3rtTOfECNbvRtdtzzcCeuwW488xSL4O92Lq3c6740dbTTZgGS/xtb
zIuSGXsEfpPkGyJC02P1vs8cNApQKmXYgWQxpJ9GgUwGRCltry8dyMlF39XCJdDY
eBFGy/h8Hh1j7Y+oDeVvJfiTEmOr9zcT9KWDxGikqh5g6SkMktwfgBFOmFL/UDR/
H5CD4AvkMqadx17LrjjCs78G2hXvD1zH8uY6HSh25SJ9CspfymJC/Aj2DdYPAA0p
sOwVQuxxe3GgBb6Ev07qpRhxW1l1H4mkMNpqDUL87FHUuCe0N7hYvyQoFzpfR/1N
6/Hd0GMdNdcmyW626IIIayZno3W1PDvPbVaENdOCyjB/s3ZkW1FNSz7qJi8ZcjZx
vhFMTrdR3VwvuhDz6DhVw2ET5dXGXgIGo1vP156M3ljULc056onT0gsveNZVli03
8Gu5I6hg8gSEZE5ZQqvAFPnfvReEHEVaaZK7g/cG0YlciQPDfoMFD25diVipqSfN
gGp8io5X+dC9+aSpKKfI8sQNUDcmRA7leI4mzxsHm5e6PgZqznboaRd0MlRM9Vp0
RdvFyV842VaA66cqoQx5khzBFXTNWl+4V0nMEQ9Zh2g522x1HJC8MsZ8/p5uGnoY
Wf7RUa2SA/5I49XgbP4uRcE5ANmxUlWQr+im/MJJJULYiSP+lIlkIqknxY3NkUSa
oZHJDzaZhfwVfkguGQ8RIn+lqXn/p+U8jfTUQj8Vr507yLrhKkL86VuO+TLAjsCC
U+Wm58nbQsnhWv5Av3/g09QjlIjojQiIF3slBJ5U3xZKN7HJgykKcO4tpyZdV/O0
sJwOv8L64DIM+9hKbGfqzrncULHX9kgY9le6GHlqqnwPBg1jhdVS00/MtjiMyfvG
T2VbJjvgCzlDzwFvItP56dCtS5UXYesiq1zobfHcgZYAK1nOXeOnD06dsMaYftRX
0ha6WWHgQ5rAHa9sgShA5hIjzcJNZyZyvk2kHLwPDfmUMTAIywtZhrRfX7e+WXuL
vHcCuby2ITmW7iGBqZsGEXqNg/e4iikVgsMeBSJkHqJ/WMBsRmS5TS95fJh5hA2Q
GEystyHm0F5TERLrAwkzTZS34ISUgLAA13EqgxoKw/FdjlXitgGYe5yL7a1Zh9jM
sD7Jw30xYkOWgYGcXXvrdgIAiIqNqss8GW7AUAyzEJEq0n1W1jFSVsefUGGoEx8F
TwMqG7MDiTop9yCk9zzk3ST5p8ic/xnM+n/0IQdlZnK1eD4HCLocVBUpeRKnjNqs
JE9483ztHaqfCSfpKicL7KQy1I8DXJJKnL9hXY6VNIbc72MwpvzV6XoU5c20OPwb
L7ex0FiKwd+2hnMDnnzkv/Cukxnp5JIznIdFPE4/SgwBCZ7I++4zSauYUaE30s7z
vQo3K7JLy+ySgKkyZwo5s0u4eSh+rkvVDmVr0ZBHJU0c3Ak9una3pYi+t6mcL7TV
CZ16ahKyT2I89hdqf6eCq+UcrR5iJA3EqN/TRfBJVuYGWErgF3nGptE8eU1k9G+e
v98YW72LDPtZDTiWFxalq5ioOoYc+7rFaZC9MjGLZjRp2Y5oYDWRJgTRR8gVNJcg
wqjabpSqL1lo+HGGsPTVjsH52CUiQQoEJuijqvYze8gixh6z2X7H5wQh1+UhMKYs
1Xm2BMNp28cjE8zE5J/1V+7NIKuuyeey50WmaD6B9YRtCsIRwcMZgPxI0M7x1TO3
ML+g70IrdwlJgt3QOb60dlvXmFfKuCdg9CoI8c/lGPvNtWJs8WwrRJgM9fhlQrGc
w7pujnWAM3N4aiqRUcsg0hFcADj4Q9ZfqcL41+qQAfL/aRx6MftJJOEx/wsn1C7r
kZBYqUTj5kHDt+kDBhhraPOeKhL5mKXfQDaDMRh55gx5mDjtAdiXLlbofskJOSVZ
saGeJLWfeEc1ZjnltkYJPHdrqc4AT5lzx2j/pm1eDo90FmTSwzx4YqNuoUgIkWKF
yYFugNhNjccr5pC3JaY94QS0GQofAbQEoRGGGV3FLNoZq7Qr/1Gfj+PwMGyKz2MY
TCUJ3VyMWr+PBTY5QryAsL06p1H07J150f1aAH67HU9Qy86qJSm50pxpl4vPuTB6
XDIe6eU1WsTL1rKuadhIF4EqAOOrDkRhAryLlkDCy4k2lxA9WR1nRJKGBQ2ctRYz
sl2YkEm6n34ZIu8P6Std6DbQrjqdq0MA3/JxssJ53dxMa6UpBr4IzsjcWnUbOTig
fckMmcJ5hxcsWMLnzwqmAWTxpxNKRB6aOWmUpdpuqVPFZGn8gTjVylbIAxfYbH35
BFz8feTSW0KXDdBoLPR2mEYxFF0bBkAr4fupDqywbNg8iql6GwzuVAUz247IbNtS
pX9mv+uizOaxICFu14Ns/hkK0Ur3Hd2QhGa1lQlQomTr0KDwHEKGbTkPzFF5ccDx
OlqVTIjBorcGtvWSwRFs9Pdaned666TUt4D/cMk8y69dsZOz8VeG8jpzDLL1kn7q
oirko9fChgeg9gBnnYfhcx7582j6OZsd2mFsgo9kHmq3Zb7LcoCRZNCF4a/pNloF
EH6SEMvtgvbEwoMVHLczKRcOF0RGvRAyxfZ5ApS2zDgtSbbxYONvV0t4lumbMCQd
uhaJyCoJHS+AgiDjrdlK5aZsWcoVYQBchMhyYqzT531N8Pb2DRvkh3783X4gkEUe
A9W2lKsWIId+Tf/aOidRkzJ26WhIhnWb69uxL/3QdQIi9qVt+RylFEt9ZetAYo0p
3DM+3/UZy3cUcbuWFHXuMlTZuWsq6Um95MUn2P03ZFuugMs14YaX9cGkg0YQGiMn
KHsJ1jnjD5LBZHpiUA8a5SXVnDnAHDt62mamcRp9aFWbpbD+iEhj6C0eo2pcSJ7g
KVfFEEN1FNYKEH9Ov60TlciQWc/qiVS8vaElRqlPssBBEq/GTRHJhSluj57aUTw8
Re4JwXItdHCNiwcUNaS24gcXjZSBqiHpO7fQXireIxYuHtMK3o02I0S7GOVAWKNR
APNt1u32ctE2iXQgqjAt5D8OEc+1w4opPPKuSfckFi3yWYCmvt8KJxmQWQWMQXBR
6leLwX/Cn45osmVMnL/LKsymA7jtNr7e8frp/6nC/D5gPQkluTyFQaooRGcp4S1d
RsyEL3+ASoM3XhGHp+yZ0i/hQeW4vQXbWIzMn+ZLTgUyMZY7vwwgS703JFKW/Q3a
lKLx123q+lAPpMrxgZ3QdwdUk0MRPKI4QBHhDMApXsJbyyMIXGh5zNBE/VXSBAb7
N5tYTBCo/RiTGE+zSnSO4MKE1nJ490nTp6zkFTaHLnc9bZGKmMVlYdhehCPu3/gu
3/7p9PwDPvUxKSawOErvi/ePXOgArj/UlYqA3FZhGY0PcAMGBx4oj+Bhr0RUVvyk
rdVTyAoimgpj0n52n7U6HVqndfJy1usvCRriXEuAJzZGiBs3CQmV4TOcszxFnS0t
OKZIYl6IXgayXDIcK1mREPI3zG+LzzZgfW0J5dZmjlBCvufM85GDLWYaX00fdywJ
aBnTsEKllvz7W9wOHfNZkVKquoEsa/hpay3NVp1EEwRvdF45v4Ft4RBUEUFs1AP2
v2fGZOCJD5knOYQ7Smr4DLMhVAFwRleL9QuRTpYKaTKx6RhWi5c5e6icMabSAya2
3H8uh/vFN1AdgtCBaGPtuh6XCc+FE+a+6pqlvI9wUQgWvEJv7UQvGuxi8z1PyTqG
dOA2IRKF6hEu9lTryDOkWralAp+K7Yg3+l478JnHVe4xgESY/l/lCzrIrd1FQD0f
xDblrXnHMAN8Eq5Uh7JOhJrIdZ0ve+CwXwue/cZSGP/Rlz8gd7g1T9/av1HVXu+Q
RV4hAxRQCkcyXKjQYBj/HCNZ4C4YMZ76iklsLTrSNkGiza4dAkyNI7lNV7IFjv2R
0WX2mJUFbASyMs+8bl7hFUgfOsh4O86Y9hocSaJp658QOwjJdIst9VTi27o2kgn/
1ohR7oc5XdexwQzVk8swUM/bpsCouWI0Avy/uat/ogdkZYf8kTfMK9UB8j7xIahM
HHfYXMYGOr4i0W1VyRmH/FUdxcaeuq/Bsog6iDbh4fv+uFfBIjOabko8MytyGBFy
PZVn9YwGct5kQQZldhvekX+eCzdVK/sovyzkRDxOCjfnj+5jZuxCP5kC1ElJhImZ
W3rGi1H7utqsnyHXiEvNzjosOZ72H+0ABZgdpUV0v7duznkmEUc/maxEe71NMmgC
dE4WokR8SsjEb5jxAQhfGFaXMcSQtBX9fTSUiKpF0o8x8FB5zdCpW4YbQ/Vmv/x5
QpAUfRVW+Hai4UHNsCrPfZOU7boDWKjcOQx7ThJAdQuycmSaaCAHTUdPymcqPP0m
1xOHi7ffYEhYcCHAOlkSYflRMFPD3Zjzk66/fLqt8Zb08xFLP7vSQobVzRFqLIog
E4s5UxQHr2BlxVaYeEtGg87/SciOtngj4V3EZOmtmCITZvRzuEMu/yT0kVpAwfH1
PK2YDw2UR8wz1Fo2VUmZHNd9+i4sD1Oz06K5209vwfNV4UmHS8vPDwCNFEQLReYh
pUB6I9FB2qvaFGjrrnr9G1zL25CuzIoXpguUzK+qTbBjQGgI+txK8UiWGbnQsgEb
LScl6krQahhvEsur9SfWSj87e/+EOpeiu5TzozCHXt3jdAz6CZteUtxRrQblPnYF
ZwX40cZM1/lW29zGqJaLpXvZWpUNNOK/hzJkTX5O1Hd1U+HnmFblcbqT6Mx1L0pE
wlxpktuHycq4+pxdp0ngv5WiOUxUVfZxAEbe0w4GZTHpuzpi6J51bxf7dSr7GblV
YnrLhiu+rNn/LE22LLtaQDrbwSgUhO8CeDkFmA28d5mBTTEX36RlOv9JBvjIbpqr
lO1oHovtKdrMz4DJU1jdj2mNQ8CJ5OubVTLneWgK6AzwBNRlGtzx5LB5UUwdAJ0n
OOXFmyi4/I1cWUFFtfmyAogqVd5S+Wm4iLNAnJ9LkwtXRY4NE8ysAtjj0tLgqNkt
KLcRevSJMT3DDy6xn+28lEsyr2KeEbs3DotJOZHZ5HFfPjlz7gRW5DcWVNbsHp5b
BrmHyEp7lngqaDWBCNDSz1cD5kIk1w0BIQ5rUsg7FDTIauYykkOphoOfYSPW66TN
LnYZdz7lEBfvXlnrcosAN2Rpd7GMeO7jxHmNZ2t+ah8sX5Y7XUrby8HWO4aXEx3U
0mx7GaXy+Xxs9JjB+0MrArJf0QjNbRJWe8YZcXVcKt5RtQoZlL2E2MMWkp7H4pbd
QDS1OXv7+488EtnlcU/fmdwa7XidNKrBB2XH2bwFFVc9CQCuDVAY41XZ3zLdz9Ji
xsz1m6zmNXA7PhcTjbc4xHl3EVmqaI5jS+AYUn/hJTQSIKIenbvclohnrXTyzEF3
ec44uljuELt6eKrmddGKqVMjfnczIO9MVY4TlE96G2V0BnqGfIy8Zv5DmKFd+hPg
bx0eVWonPGdieGv1Lo+6euIO0rZNbb+Q3wTdNmrdORmBgmW5N6Ug0R/MPGio04RM
CkO7B357Z600u0cPMeQiYCEj2wHT3QUbKqCr8q+OuhoBcaPjuPFf3y1FOOUnY3zw
cpEr6JyUEep5Wcm0FtvTGIaJJO2NMdXNiJDpV42UaH+/AIj7VUgTUYmYfMr3WQF0
KqMRfxRBAxFMPGsVmpHllDoEMSvZNLgVB72lmIT/EX9DyPx5a/0XqGJwcnNd7t7x
5kTpyqJO0xB87G3/OW56VEWNjpZRF/b2Ky7+G8uWCAeH/lzwSzFDmOxITfWs+6IU
XAkKYOBelNJyheoJjDUlozeaQtoDHLk1pHztbvTpGKYuD611XM2LBVvXi00PPq9q
7MgzKF+9nowmaHiQTxReOg8h7OdrFNPr3vTqpO6dpqOqD65rQq5U8vT5o/91DXGY
4ncQvEIt5V6Nqf4uUkfMHITtVANtmtYOwic9Hju/vkGj1HVmZIL1rZ204YeY4pZF
tppfFoAcp/19nj2BRw3tUaBbj+LmDmS1G9+JaN/PL2OT/AdBUvqGBNUr001tQM4M
tD8ACZF9lLC3b4l3dE98iLsTJRiVFDIDojuyyIqLwF788LkFDo6NzNwRmPq2kP5Z
zcMqs1SvcrAl5wzUIN6o25UbVQD1RU3pjqMaFhrHY6mD/qIKI1Ggz1rvvDN4N4rW
aLb70ALTlL16myE+uLE2AD2gGmG6aoLIrPblCKgWubCDyTDgWzNOtnsPI3vS58Ik
sVzt1rW5MPxgyK3riMHqK3fBVNdxXYayKMGxSKwEVmcAH7olya+DnJ0XJOE1jlLc
fppxxn7O307mw7CvkIhVCWG5m+GjMwO/tTTLVnUmLVxmDZdBfuo/HtNi8SFi0IlL
PVl/6cgfgVZMojxyqzfGwlZ5Zc26yuM2BvfHsgOePb940XZL1YUlhpDzFdObL0tl
e0VPN8M/+d/bFIXnZTR0pR3hYwhbV5hLln18AbrtosyO8G3e7eQMVacAoN9ITghF
lu7uZUqhL5pEke/Qt7E7iyPWHXdSiyrdC/nm+fumXXVe8R6iavc5717iAdO73leT
Jzb8qMSYAE52aFHkbQK/+7/79DKzCC7ZnAM0uYPg2GaaM8ss7pYNnAeEUAR5hmHr
rWlOcjs0OVTLx4TlfJGcrSN/OaK5quK0if2ukpQHw6Unup9/GGVRkIUarmObX2cn
rH9T6iPKdnmeTaMa2mT7L+6qL7V6jq+6PLtAKaARSI/stZqo3GB0R7Xhz40EEpsh
kfcr6lKsWLvIOa8Ai7Nxdbbu5/y/q6jfgNGp6ZEkdza0dXplk9oHz12UfzV5BAUd
eZRS4AvHZk77fIBUICro0630mCGJvYHAAapAPyI8Y/BXwmSqnKHPxlo7GDq2YPUk
gWNHe3FxtnHmZP7OGI4QPVe7WnjT4NTDUbNkddEvENaCzyQKHRHtNbhJYow9rXEc
2ThAz9lnFYdy+wETMBfayHfkv1cdkxdUa0bTUIl3HoLrSIxvT5Efy0gQX/Mn+pJa
rOG8FTB8NzhJD0jp8p+A5F8sJpWcXbdK+s0WCedWx9e/o7oCCJsYshY/5ynOUUpD
yE6TIrCmgSsVYF73B/g/XU9UG7NhnjVNvRpsCy1ZGT3hwx3CETRZW48ushtXipwv
aw6MQTFwWVZz2mBgskMFSikYh/XW8Ii/BjJexC+0gTLibRZR8AIALis13bpGXjCj
u/YFXG9QFCLabhr91gC5Y7CSAivg6gocMpoJeo0j70EQjK+u6huoevKoRjJC+NxF
dxQ3SSfVRV6wC3TqxoIpRufZ1njVkwxKKVrXYt2R9JPDbzqLFGNqz/jr1c04Uhf9
VpFJJrowPekoCfgqwwCWBFioI6ElyiVEEp4E66OnH4lQKDpt2NfCs4SuBveNXb7z
6nKMSPA7vJtq1huHzPzRNGd9ChZNUdvKPt+hqvNhBIkXkb7fAuhedwRu8aqoWzn5
dgbKgpIflDmoQm25MuXsZjp6UoQKX9DQ21H8WEBT+ACA2HkojuWa2LpN+x6XzKZe
jQy3GZ213H2imSoOPr8UGguJzskGaqka0/8Ah/fYR6uym0Vj4h4aQD0JJV0z5jrw
JAmM5ksgid/OLm4lZezv+Fp0/bPHC2SFuckKx934Hr7GWiOMB2e6csw8PUEMV1lp
PpwsSaw9cc8rE9yO0CUI1oUcbXYz+alkerldlk2XMPmo+ji9yFhcTyRg8dW0a2b3
X9wHG5Eque6I4ueT/FedIW5jXWp93MHMSbK7kLJhrIhyg2TshMHmXwzbAlB32AMA
s+Z7mvswBGgl+bJYlPvW5HJ+QrXycHNHHta2I57wfe8Nw6veddOF8UOXhL2qEDdq
qXXfeko4o2qsTfKoWlMAZddCLQIdkw15K67i9Fu5gdrek5VcCSDYlhtIZ+MS5HaE
WOrGjfRU+Ew8I1B/CDLv46Z8rquqQmr/atfbVDCIsJr8U3RfHg4LYC421p5xG537
MPYvc+llIumpJ+LUgfL6sCIrJUfk81bFXga/jsMrUHtY6R/LjGM9KQmlgRPQ5hx9
vF+5kgp6iCXUUlyXFNXBg9v0YFKYd9b9cBrxeFuv1kV0w5MKAEQhI2RrW5gFobul
2pB65+Pvs1o6/9STjNYZe4dkyvJyPrFhVS0uJCYS1bwRuD6zLNI2ZmhJfXLPM7rG
gvSyaiuyb0+fWS+vnZgDWYAfrhgGTYd7f37tL60Q1Je6XTcGA/dtOLYWIi+NEcav
k2Uh1e/ETC4o9j2G92Mj5h659j6ngy8phKhzVWF7xtJumFxF9QjeAr/vKsrc9p4F
4Nj2Y3kHeKGdGchvPrKsD9XbmVMY688htRqyjmxmMx8m3R0VW2hM1OatnD5txRuN
VBhQ9H1TMWdjq5Svn6xRsWL49t9PchHkxu8wsZJHou89xYUzL4ctvxIQgR2dtdDY
GDTm6JeEdsAAGZrSpshnrIqpbEs5qlq0BEgIzLY0CVZHr3ZPciX81s1/DRgKWLdJ
hPabgOVgmIfR1kR70eW1iwHePhoLwCi+81qaMdI/Yt8LJLV0mxt68OD7su3/o2uu
rqQMyeSoTHnpJqn8R7fuRzlQ+RGwlyPQ1vz+TYv1Q7Ntnx9jMlrWoIJOLOMxxTrM
/Sm5FAahz5kJXQKNSVF9HLffqSkEoSlNKEbB54j58iN8dqXMFKr1c+oa5IorJdFY
+7ziU374AUrGpJOoxgxuyuB5cafHxqmqAseY1boY/TZfvwGS42LjqpIAA/4pN/LR
KO/bOdqxsQ/LGlFV0n1pwY7v3zsxOCy9IMx02FqGWIFWN/XxkbEq+mW8j4X6lU6d
aq3/Eoor1uSqdyrfIA/MDukkdzyzNRJp1RYP8IuNFWnYCQFwkvEXz4N6VioR8M7B
AxNtWpn/euATuwBxmQGycpRif5r7EcrqVLNDpIrfgFVLWhrzhKRSJEibAMZQJso4
fvCstjP6dAAwsy3eGqABMkPTSw8Qpxm3PZ8XlJD264vFiudjktlVoe8mxdECp8bB
RNfyl8KBUYfiZcjB3K3915U3E4wEIy3ajtfaRj6wBPCeoVNy2heE8nqk1D34e20Y
93Ix0AOUGztwYKUGGXbwyfoPQTfkrdXZ9D0xPd8w9o8kN1eJtc4wrFW6Sd3AyAZz
GGjtC4yW1waPPVQrStHvKyR15lv7bMTr0aBjlxuq/c8tORhliQe4GVffa+zmIl+V
KKsVPVNTZWhH1hzSUmceZ+LFu0yqPGe1I7UGOUft6QeoWOVU0es5usx3BnhlBsWv
AKRMlT/1oYbHZpoc+nEjf55cN3FfK7ecqTDhbOVo1jXvMoAetnglVZG19lRDno6t
xbwhQRTMz5z1sd6q4irnsA6qNxCdDcFf4S2o/WVG6Gy4/HV3do3bqSG4YBUit9GS
o3xCAB2/qfR0SH6NbzGTaI5wZY3wta/5PBh4Z+TYiccReIrH0jzd4n14a+oYAV5F
aJszkngk6qUlgiaOcycS9if+t3vHWpDHD37pxXc7YnTHANZUx7xCQqaqJWFsH/8I
Jx0Q9F2wHw4FxCr4nSvAp3KA7i51c4ahAbtMrytFE2/dwQFrA+Ge83P8mw9U76Fb
38/wXnI9KIoVPuAoDKjOCaK/AGb5BkHfNqS8+gwtt5XpUdcfZByK9+X566I9rGYU
JyxfmjcNHbbrXo/AymLPD0J/Fefv259FJjwHOG3OeebDDSnz7i5DZbJjjmWyovuP
8F5h5QE/bpRGjELe2A9QUSPqLEgkoBI4L4Uz8zvDONLU0HZDlFPbNxFMHRCS/mLd
m/pjDYOBNEXHie0nrFyMFGUZjn0M7hcARUATVA8Nhve85638G/Sb/DOGCE08FSuJ
KmlW8q9GUOMeQrSiZCu87TKU80RKnXj32Ruceoa0rg6eOxdjZ4Xov5UvoM+CzZaY
ymbFm+ys7sID6wftD1BTywvDy93VQ4sGLhwAbB0PdqRwfWNxCIU1h/3NRWXgJ1Sg
Jx46WalJaYRDUn8ANAyrZzwbjd36saAjUurCRwgQTpmncRtEX2etUDN9GrQaPOV4
a52Jk72TXJOKLEWVN5z4iRvMLYdIhJBj5kkInc20DTZAN5kpIYEZ3Jj7XfD3Oz7h
fdTnx882Lt8Lh7CCIx+sqlLMAt2FIJTDdfeQrrdMveUPBaDXiDbtPXHzUWQnq7Ik
I6j9BO+N7cg28xJIIaUsGRW9gDi9JpRjHtxec3VR8sAmG/kZIlTJz2LfiKOtDvIL
3sJnyngfbczbYVXyfcI4fxIT4Ugt67+t/7BNbN5JAcmC1VUpiZDtIiWVxyRl6YRt
2awhFhVzLRFYIznCfKPKNQbsOzNGIGujHnN0koA4QILLQJE273KfEjeBI3p3y7WS
OI5UEzG1r2hPi56CMBRFxKjBYfmhHMLjq/aVXKPkcVG+mbspxEcyU8QOsdTv5U6m
fy2JKaAbmnGUaGgIJZijX2G3vs2K8ruPSBuuWKx5GqB4wg5LKRIg81QHf2WnCRR4
yHQQJz742yuxJjbjt8qKNVY8Ok8bchA7hoUA9UOnYTjbafdk98TWkelA3OabM62a
cfPRBr2HkinUyHsVq6SiuA01vjFkVjCz4snLFdHieWtpiMXOcjEpWEDWfKUdrKf+
LP3RBEMcYOYto945xf0IDkWY7WoUhwyhLi2TtO3lpZfgEzf/GNhfq/iUUTCro8WI
E/hk2Pz4oBamF6kLWGAGMTehf8r4M/6NPGFhHQjkVLt5Ue7qtFH7Oj8SDd0z/H19
X3UZN+jG+rof4GnWBWgvy1yOZ5iY5oi1XO2/EiEzLy0pORbYwdQ+1tam2R6DkJWp
ulbO9oLcY6nX5Qo6PA4xc3kZM4nPVQ9U5Z1SjDaUSkYUnHV7b8ThA2l9auvn38Xd
GkQyYZ553g+tv1Jx/m68P5USyQJW+Oia8oSL/SvLWTdOk/ISYrJgVyJnRaG+Jze6
kmv0ZnoA5RLl+5rIhL3CDc/1yFjhZ0g/V+60zCmxVANSgNgRQkZ2gBqnimZCSafq
OcEvJPG5RBsi6CGJEYhlXnmCIchAHntrDDLbZMkyqfo3mQcnmHbQdleWfYH/ahzr
En7vbC70VtqGGUoRWs9MeEMExArkw+QpuQWlFJdNDwurT9Bi6+rGJjMqppJ9Lize
wWO3VKCcT0pb8VOnhZdISBjgt0VDx+J7od7OiIsytPWYD6z5y9TZ/5/SBDwnxbQx
Ya6O2qG6pKQk2RWHsc8edbQJt0px4BBVDxpZcecRjT+m4Ofh+rDi2wiUednHuv0/
ZPAciwWDGnwJA6AiKNLyl3agIzwNXmYRHam8z0PQkaRIEPXwhN/LtLdMz5olMV49
HsoRCr45B7AFazYu9qe3j7edlJaP+04iK0e/35o8onWLS8h3D0C1YTpaz3KR4gkQ
UfHwDaNdKjlyK2lwElV3CrwAqAdtZh1jPU9t+lB2ro3Ig4NV5aEp/iEetM2KaEeI
Bj1J0ZnEOfjKnYxAdQ/cwgFOuwJBAR7/qNB3lAjmZTFQSl5hCKtEjoskyT11MP3D
XRT+3XOhe60wK/HibAAQ2OCVniygceSdDMLZ1TlogmcGcb7+JUsWc1N8byBYYkdH
y2AuNLM3w9q+55I3U+2bNtmgyxMzeKlWF+bsV5kAKJf8RRa0dspF3iKYsvom+6rQ
2FwQiKgrc8590cgfa8w/wAxdkKX3uWxWGjyXYj5vfJBWjXPAMLEaY/e+o6iec5R3
j7G5b0nGoouwEYbaO9AAN2zXzhbnDEYVJK/Mt5L3l4pt/EwYYvJIP22Ix0WYKndy
uphZ3og8ZnNETrpj+C1+MIT4KdxSFYT4QzOs+1eeY2RcuIuHEPWBenWOZdsQgLfc
rtUAVIzGuT33wNcx8ZIvNcHZ7d+155mwSg6aneEdH841F9nT7fhbtF29hm//pyIr
k6wOkku/YWfu2LHOHsrUBQgv7B6uS41mzzM2yilhqgsH42I1J2SiUgdJTY21UWHQ
HTpqpR5gM91eMU9q83zQUAP/wKlG/y00VDUTxrD8aZw0PwCB/9Sxoopa3uiOoTvx
fwWWY/NtCTDb450y3mVfpf0aBi+tLeVYxQzmiG/e8qd2T9mjY5tH/qEX0NRho9kD
sirwTiVX8s+hbe8EuGVTebpUTGK11eyBQNF3Rx21cl7X8iVVD2yxen1tuy0dx4AW
+0LNDrCoykBnDGuI2iNrZKb6AasoqazDbXrkXsQXgXdP/7Hlfn77+yiStnZORm45
Svzk8ApIIRZqdqAvqgyAWedR9YYFosfLgElen4QWGn3ECqaZ2axA+vz+1U1FfVRB
j0RVHXrzSsXCkJ/P8vYn5qsuv3DeGmZou3YLUj7m2ua6sC6YC9YY2bUpeq0Q1sMa
XM0AxdgFOI6vDmRcOq/uDyefrigUV3Ft2Q3L/l227nFMHAJlWGpUI9rlbWMOuOEN
RssF17wvU2/o+sxZ7PAGz3KPi2uW83yXyR6siY2D4zbV5dc6XAqgv9MwB/fPCCqX
4/SPsdZqBnb3s8Hg0gwJN+LCashwVxZQy0jmppYalcXE3O7fID2D49Me5iTYirk9
+QLMl5B4PDlhj/hyHJZSFHUXcVc6gbMn573tztG3tku41lRqjV9VprAnSjjo+SYM
P28ZrtcL9/XUyz+h/svOadOitB3fAtkxcfAp9GMvSXOSix+mHCD11gsyF+ktRjIy
zk+HiD9blW7dR2+8ESrfq1R7Ojy1DmFZNuGmdSNF8S4/DGNEfLRy6Cgelk4vVEcG
kj5I2+EubQL3kUKecL1ayXzI8gWhPpdyAkVdglBQAMy3pXhqSDbDyPvMvvxpGoJd
csRnMCAZa5M0gZblbTbSMLpelUzmD+VoN6BPDu1JJh21QfZHyYyVRrHb691xKr7c
jVBqdE+CBZcSppHvfqmOIiG6GMSawM++KPbCjMkN/xfC9FHPZavnqY0p3X7xXzB9
+Br4Hq3YTIVQtypicw5RVu6dcJvMohUVtPhxHqPsKBz2W2O0D7J5dVvuXDQvYPAD
rRtRaCFa+0HBAK3MBcpf7pLhE+LP/8O6Mbogn0wPOiUM/4hyaOGUCqHgFzNGkF35
ZQy69n8teGxANG1VNB0xp5UZLSDMowyveDGnwpRIQG5nP4q1ypZCL6bfBsXnXlek
tfz9xiVtIDp009109roIf+vUufAoFaqa7qonUOpv9dX6X8dOABrp7mOgyqxtNfgO
qCTYeWO5Z9HEXuL9sOilLTkSGLpPfQbIIRfcGdtEJTC0LNbU4BXVnPX5YlcT5tz4
1l6xP4t0/BPe13e+01g1k3YvWAw4Fem0qfF7WJMHmPTb9u9n7j5+zHbWh118omGl
xJ1T1GQFk8jVrAr9AOGbC8gecl0u2hM1zaLTCW7ksLI3rXK1N59E3KW6+ANcXIx+
uz62CONty6SRVMJJnP/VEBtQuRMj0P34a3T5uDICLNcU+Aob/8L7CfmAhtZ11FgE
jHIp48kVnP2PchZ+QK+TB8w23fwVpT772ZWj2LLPMHvOjcmXhIu0K6ZNe0BsYCLw
t5NehtUa3saU331NnrVHrCFBWc3/6YyTfyfdtxh6U9yxhfyOP+xnxb1qW7vdoy4G
cfB/9Oe/NNdkZansssSZBPUmp5GPlQMqoQQOubOASezn5dUT9cvPX1097zhXwbPS
3dDHF9QNpwHBqFflHFIuKm3G7KfWoS0nQI3LrSLomt6CBS9uyjmtOj/eLVsfBvly
ys4TJY58oqFUYM13+H/+GUd6P49J6qX6W0Q+ZVLW9+eOHiJAG7wFWOoB62dm4ZKb
wB4olvNBuRaIsaywPcuAhUpKwA3HGPyAVuQaJ+X/fXHa64WSyxU51213q1wq/9oC
Gk+uG+cJpHzeMFNtjIbRYD7zb+S/rZSeOQwiC3toXtzNUTxrDVuVHaxmIiw/WVJ5
HjYRz0hfT/gqEW8nBAtyytZh8Z6wY6bEk+nllHyoFyfn1yX9V3hk26wls0/6ku+F
rdKfu8NBJwT/QrKJFZ8gx44+e+95geeAVe9AhT+rQ6IPOh1INNMqIYoYpYbEIE0Z
XO4Aekdz6GSBARH/Q4qWuifywyW3LQqcxED3BsQW/XuM1VVei7uUOugXfL018TKj
jt6W0S/TSG1ntuqQvEM9pTb8kek8lJlgiC6gEmSETXJQGEJV/kR1uvHILpBo8/d9
DiWdSZqRCNB8hD72MmnELnPbbiLzZbdP0MWWNTwfOOUXAeAmQAgJnGoU9yszCfCP
8X7CSsC6XDuTf+w+Ay6/9X9tJO/JXb44s9bBT2HqMAV9ievPUzb2TRk6VMTo1hRL
ZvyRsCNyG8rcB1XL5UvRAs5wL14XXITsZ7sZTwE3DjRewTj1AW9QRnstwAAaQ7aL
D2N1rFrysTPPVFjN/N1cL7q0vIUmXAY7+/H4hrb1o2CZyHF8r34morvRadWe9eII
7tY4qJhEUTARz5UOKoEXuUBuhb5QLDCYoN4C5j23TVfqbWtD2Y2LOfp77Xye+3A+
8cCf+vtAAukOqU3dUbzoO9CGQMLlkqApYZOLM3RO03vyKK1vo15b37TWhoT1LizA
Vx6ZgA9WB9D25R7bCqIAcS/AkXex5U3556HqRzOegIadw9KFD8inuUZPTaeEpgTU
yeOGISKqhpo/w+AJaFTlWRTK1r1oiv0XBO/kuebUtZPe9BDmRZoQrb8voEOA/iK+
qNjBm/f0Dhssij4fJgjxp5QT1PRuX1Wan9jCiKccsFHyGbrJL77u0oLBsAPIcZ0X
0WNp6BVi22a3wXJVvnBZK7fRQksrHsDXlpenKtelCKMxTQcUcaH/ECSq3/Oorfb3
9RvsdIlyDiJBYJb21C4TwAcdfLi+YeAhhdhzzg5FijA3F3PAuQJZqvjYMCtv/T+5
C/nZSHpPCWg03pJwXX1JNoAJFSAqIEL5CUDlkjIJJNDqM9/RM0C6BgXS3sAKrLqw
tfkNOHJ05YWVVYqI/oWELTg2nVotBdE5NRpmRJEDzEVR7QKJf29WNRm1wUBSBlzn
CJQ6pzdiDOOUa0yG6Wu6IOWcBZPG36prAYErFgdfh7JumkM2kYlNJp3/qz4tzYs+
NnegIxBP/Xg6Bj/1CBxtv3JQVRrn9sSGhh0ap3SbSrCEiVqxF2UkMASSWPuJsHpi
ZbxtVbUKFaqWg92YdY7HHzXs404ZKRffYJxs5u1M5erMWmet9B9XcMj43rUxxuH6
aH9jqnPiAwkN6q7x3p8CEOvjXTIfoH7yMgHHp/YxvUDRWq18J8xSaysA7Ho4aign
2HRpFMn8PchJewQj7C1TUs/3gbUMxru0+N/gUNwEiuSiCIb89tjnup/HYUTVkeVe
LQylMWabhV9E2tqcDoQ8truiYSugYmAQuZWDK4le6IU07OEIrrYloMyrx9Np+Wc2
jz3Pb/OxgElWY2dpP+JMWkPePtSL2GwvAdBM9gCWAstDiQNQDPo4b/T1LVWNfmh+
t/3jY1FeE7s68YQwRJz7pHOKw57ToHXeqPZQRfyXwNIhijvycE4y/jebomOR7TMb
qXHL9dldOVDUzz7iBCbFCeueN5xWQ625fu4pcDgrnxK3Lvo5i7HpzCNzDmMVLrNA
WR5uB/6e5rJog1GZUVlVVFmmh8zhtH9CtWuIJW1TMEJ8zqnOdCq/0VpXq1raT4de
8zHHR572Yf59mTnzL2F9pkpUEwJKMM1cJv/xf2sCAIK4HvwVftSRP409jS7oY01Y
10YBZ7AxKMq2gy24VZOXG9AkSfKqUblmqnaCD7LtyE39TWibdsGe3My+GMUWzZKi
PqvL0EICuQzpyXMQYh+96f8IvKXHhfLOsMhHCjKLpAz7QE3XSJRFhsAWpxMy4Ebk
ljCjXjGRm5l/jrKDV8QJ/N4lgLKDxg8ipBfnEuI5Z5S6xZArpnN6pZkhGs8y91yt
jG0hgLCtpIUNyjM85W6TC9O3K16IAXTFhYWq1hbI4RT5IvJTnz/FnGUMwHnuShsT
VEWEImfxAE8WFYLROVMkDa75xhF67Bc9NWXt0l1ixaqhS8fz77tf3F8K4/w4wtCp
rucqEMcn8rjhyn7by9cTrsymfxo7M0/q7DoXmQtXwQC493Ti5PngPgjM3p2BvkGo
BBBlfmVJga3B3A8PXNJlvJ3wHsnCR41KaawJWjys93aR6VLC+5b0BybR+9u6xpDu
6PzxtVyI/9ZUcPxQ+NL1Z/2KttO5VYl1qIWpqfhQR40OH2YrMCFnhvTLT3DCwYxg
XMgS/iofmPqxnEalWd2+YoPAOGXAJ4LmK3xy7Ixrq6O1kI77kz105zjBazVv5qKf
deEmoPX/zXlTkrWdRxEIygSJRVt5hl4AhkRDOuFCsJoqaJ8CmKQP2E1JaRpVvpVD
iTpnjbn887AvvoJMOy9FyHej/+BMRfZlDOjvYYtm9KJhrMSA/92Jrlx6tW0UHUiX
0c11DmqgBWSWEZmbX/l09Msonjv+WHNVLy1yHTy1nKoUizbfOojjptO/mPhnzi5O
Ji2+LUxYEh0z7qFahv2SzI/61OuK/VzNpxUw49nqWBMvTvi8/KoQOdGJFkF76epX
Lf/6XL6QGfYTRHu7DDWY3VqRQQ6b+MENz3NDrhaeGiO7SJy4LJXpCN34rLf70rpC
vwDEZCBw8ARY65INVPPmEfDvjFfRRY1uwNWMXrb5XwUHCKOrQrbyyrBUt0RXRyA/
y1ErIxNSAmK9kA152Oy6e2mo5ghm+mwrUIwM4SlDvm1I8hl4YF9RYDq0AyNHJBMT
VIbRUWxsbQ+QX1zovVPB4l+1+frUAaAWcj/cG7Gk8vXtEEUDbRD1aumL+Iq9q5rF
i3n0QThok8l71oea1W8/lRWY/pDrwi9JaTvEOKF8Gr8zZUfNhNZplxjK9tnXqBL8
P9dZIapQRzLbh/dbhAg6L97lvp4g2qghDCj0QwabJsvk3RpeT1c5/Hegi5IV/lmy
cEbsagF7qqUOJiqFXv9PgQjbsDrlK4oqP3NCztU9Agki9nk2yApg+QsvHmI18mvm
V+CAp21Dhv8MLQNDAY2ql1Lb9XrB7d5ssG2LOIP3ikaWl/DEZSITLRDAWgiJ+Wnp
JAo9XMo9abbXnY5znS/0eRc4No3OoHNhzkc1l6gEg9ysBiqwnXPa5S5rpS9wb37F
++IRXR+4GePX7mSLn1EG6x2duESOw7MFMDDdhYGCCzQTai+Awn8VtL8IBIEOmwB/
ferfyR2sBIIWINUurmZW354k37o8W4TZgqc8KEzx14rVF0Tgc4KEBrz6MOkeGBsj
ccP2dHyAxKXhXp5GlEp9DNjldacw80vdOoVaYzGlsVlZ6YPb2goEbxtWVO57ul2O
lIZN9G4x7FDT9cdQfBeqU9ru1JC3bwWzVpe0LwJqq4NPkI7j45TetS970IALnZmk
9DnItkRQFujBh3VwICxLkj6KN7m6wR8nzGsCnV6s8+qKAk4QRpXneqT++tTyWbF0
g1N4+Dw9Cb+z4AqmopMxzMZQlV5mZ2/huJeQ+ZK1iKWmRfCXZ6iLX7qcQCTCALQS
zzad02qepg8Id/XTgurtEslMegvy65oYshQrhsc6KnqON8EOn+12mTgWEJkG2XOc
1gNcY5Jo6+OX8miu/5EodqlYNK/QnGWIuwJ/bArR/sWoKrrPW2L0zZAU25gzBFHZ
X1TPBmUxekfPswmGHKZZzyCbcbX6ECy6fUEpW8+NAE20YbONVMD+wivBaa3fkJ3s
wtARdvYuokuOZcncxkt+UJUFZArIcDnozWo09kpxvPim4unFbgMKQPOZ2Y2Qhy61
739Xa/VMRNrw79LiJEymOV82uGRLvv/Syh3B3mRtcEqwBCwcZcNLUPSySUSd/UT9
05DNH5ZMHdlb1YeaUJNtWEZtsI+I5Z+0bOfUq3T3ikVQHgg2+5qmqCEt2XPaHUN7
UrzjgvcA0IyCc9Lvs9X1C/WcNUk6uMr2XuAdxAHwARCOsx5EmP2lZ+myMyRCHKp+
Cp7/S3EH9bUkbfhElp4sOWLpWxyh6v1Uwi4aOvTLHMNWfs/GeLktoKdRq+bsSmlz
VWN+3SOUGgCkxnQybw2Ho3ZWUeUN/PZtkTy4hRb/vgxba02FIq9ByHp7PDJQZ0Yr
2DqBcfTUrH9eUUAKZLIIvldcTDBE/h/2Aw4hv+ahZ/StiU4LV3gaKgskAI9zhCQ0
3Be635dN5fp90Hfw+qn9OzGQYBQjTt2piQEYh4RVESoKxp8LbplAF7bYMLSWlk7+
V84DuFhYI+AQSyiyz0zd7GbQDV+yG2TLPOt+sdG7P+VcfE75Mh2zEMasWB0v8sg7
UZxIBMdEOAavpFALQUobeUqZlYuKUWumc7eiPitQhDCVFqnvSE64jwGaktoxT5PZ
M1jt/fNNEHvf5CsTfkCrHIbSaLXiBTapq+39nK2gb2Wn7gNOh5mCuyDhR2rFa8cY
TDr6EQ1+5/c9H6y0L5vUrFff4YR6K+JcM7ha0PZ0Jo7cuSGM2WlyqR6tLcrYjY2X
yhxHxHKXVslhMA/ME/U7S+oP30CVMm3+Id5FNcanBLPykHwiHbkX42jg2liU4c80
SLXFwMTCv6ZlvoHI5sfEeB35e7zkZMfR2Hg0XjUSjNGIhKukoDgTeQeFC/OhyRrn
omyHXUiC+jFxl1EnbYfB2JTUzzMT7Ts8+/tiJUpKQUH/3qJ7RenpQAem9iSN4NMe
ORETpAsiNR5oPqCYTnvoH8xsJorPisYCrebXqVLh/9nEzEgNJk70zIa+z/K7Sqh/
OKMqu0B9Gw65H5dKoB5I8P1x76K3vLNLxof+zu9RTe0OpRkNqqYeuR2xMLgj1mtp
tP+GEVyKXDEMAFoJMbNZZUfTqhKlKlVW38sX2QxBsysQ/TaBm2PrBcopXhZVBArI
19twQ7gCsDldECTH0Zexep0ckASU6QH9Z84a6dpTNTtnmn+JS57sFF8a5x2Qwnr/
CXpOPGB2d3S1cMjqndtiZxiKmriIiPZjN636QLJt3JpEMZmoI+CSjRiZxkccuHZt
0nmLcfQ8gCM6+BCE1RGLuFaVYo/WuSiYixHadu4dg2h9KGFLnt3Yk9z5HIO6+If8
lCmk1KVNUZy2UkYN1A+mpZYPzvo6kQBU6a9Mu8itmaMQk4wnEp6dOK3wu3+WF1sY
MR/fcDhXDanfCxbTnV5J7Gz9mGm+sGCMfytZt5YC87T4ed6LSFWSR6Ds4++EfwOb
beRlWDTe6f2DL5TQ3nHdGUmTaz26nP7IY35l/3iHCyVvvPIxZaY+mVntqiB4WDHX
/NOMrIbKLkWmaBl5svRUKefb6kU2nN9PQazjEEGDD3JOn1okLU5hjeWuZMwRY1W5
PDTtqFQfeUNqaapYaNXG6Y9yfyLYC5afTZQE2jXoRK1OYVq/SpzVA5bqHz+8ZlcL
3xVfGY91tGGYqGWA/F/mDtmkOD3x/vkqZphAjSrje7ayxgtk4N0EbdvhMq7maOTb
iREOLHeZvfS8f+SDvO0/RlA924h40Sgpn6GVQGOHHWwbdYH654vw1N1iKZ2sT0af
x95usu2Hnd4DrtBG8ROdhxv51cCIO8tor3gilnzYjGwPsV4SUUhWFKcv0otlTiyr
/hqN6YyIwISimLntmWxkp2Fs68W/I/JFrUHbdP92gGckvMPrJ+DH7JsGY+KUqb5k
eV5fMfSTIHxLpBXqkQtbcO1cEVKhKLPM7IGDGGMo2LjGtOe+KunUisrMUCf1iBHC
qyvI+dAzhknEl6+CpSiYSHUoEwcFCF3jGmU6FukIh27JUdw03RJJayr+RxY+haBc
XHq1/SFIHsbdGfuS/G/Ws8GsUxLr+DEbiCxdOMhVB2k0Vd6x2666fd7oDaOJzieQ
YvIxZF/s6+Cw/KvfSE4NQWy4j1xNXV00Z6a/FYrGtCrSl1uSdDJbAUBH+/3Tzmvk
n4vIkNnvE23RWJecPasi/VK325GNpSZKUypuW2Pnhk64NJfxSdbU0ID3TkxcGemU
OCdzTFl1buvJ6oGT4ciLnuJhV2EQ+JevxHqR6Ww7IV0e+3qlyJyq1Tu5Prc9fy2d
qR1MphBX+5OgQQMwqi9KqviJS4bQ0q5wLFZc/wICvLWlXE1Ll4tRJGDapDbF2Ez3
JUL2T5JW+n335hwnFe6q+nfjDysb+Oz/v9gP3MtJVvjCqpO5vXcpvgeJ86F/P2U+
Si7ckTRa3yBPgXnAfSulc+LcZQ4EneymPPQuCU7p1ZTxx1+N5kz1P/bfH/Cz8qQv
M5BHZYpVQoUAXCxUUqhA1+KO3pnCUuXU/CLNq9l+gC1GXFbuvT1VUKKoAYdVgj+I
MqR++jH/AZZskh+bUqK5EyGyEFN1XB7+PLeK7rhV1ELw36uPxqD282WdQBIXVs49
EduFSzTXpcZvow159sjJpLQnuCnSRqL6AMSVZnMxkaNfnuy2te0KI/M2OwGe0dvR
NIzqrUJryHiOoD18SXcPp74zq/Gs8/9cJyfVJRkhvlxUym2Fa1B99titVC+4FOVc
FWCob8Dy6yOtIGgokG1ubupyLty8i6g5bn7BRsrrxqYXuxPrihANT6NkJGDqPqke
dlRnMEGPrwlBi6GbYhhqayVGyg2R88uPCdNWZYnSGsUWEDV/1UK9JzsZHxW08CNV
ui/UtHZBE/ccN1qaaO39GLcI6UGexorWf3bn5i3KBS9HdZiLB+IA6VHRLOfr0f9N
kzc7q1dgTqthK96kX+9FsYchFkRh5kMQR44OQ5CDJepaKTHFQ63FA/kyLlC155Oa
8B7ppw8uIG0jAxBBS+lBcLJNxYFSLPw9SA0I53cv4rdiBR0QI6o3OcBiofc5U476
7z0Fc0cK6jZrpxkZucC74PA6kV9Djo81avj3vyahifK9S1sQtsULp3KXk6HfhmyO
5qjYqT2q6HwOAjYAp1HBqJlPMtHceiSxnDm1oy6OEXIWq7AtskAmfL2jFntA2wTp
cNEmUEg9BIcwLjiyxx+XqFjsqdDjXX/MLvxmLuKLg13RuDkQP0TvgzZypw7oNMbP
ZmVYceygePDOaC1YW2S+yzKQT0aaDN1em1fTkwRRDWRp2s8/i4agEt24YAq45RXv
nMxwjvpw+UB2dzE1jYhy4Nr43TEDfg9xiYvATH4be6oZL7y54vi/hJEC2bzPbZYw
jDPKIE2lZloFoumPtAh9aumHyQEU9LfuOun74cFJoth+7psU6hyFgeZUpVvjRUC0
x7E94xr/sYUXQw7HrIX00BfAePy7x3zXWF0tYkDEHT6MtG96IfWcvJB3cXL2VeCU
Dc3Le7fJZmoN29A47/5rVb/v7vwyy41tmgi40ZWnbXv+iT9n+9RuFCwH/G5bi7lR
WNL58qDdH5G07fFqTW0GnOiBR0h42Vyv7LqxU4AuPkiVRqhbdF7O3cc4/b4G/qpW
dc7FXrEYKBc15bMrY3SgAYXK3GZ+eccnhZY8y1m4duhKT27maR5S1X+oXrT6fjX1
OlEx8Lbw+LMeLTumfNCwVapsH+VRxMrTS2mmT0SDKXMOlnxgizpZaxIHzwr0LYp8
nd4s62QmgGfLfRcJ47Ii/GTOUYih2pSfozFLl8kNqw/82yzf6sNhZMsn20uPWOE6
i1qQ5fy3WaKt2r8gGgkEhGioPOMgBque9CQoV1ajsWMJRfoU1bBkmkZPMSlN/UHB
LdBnwNS1kP3P1HmrmerO5IQNbwjAAH9JMkSJtg/9BdF75FfHQJSGVsmuU74ZF5oo
64AlXO0NyGlkNA5iAdaeRyIgzpKleUCK7z5n+OCq2qSXC5kSvo01BerPlayoTRhe
5s57LTkYrWzi8pwM3bktp1oed5IWDbbQysPnzTOWDPdDojQnXnIUfJphVQRJhH4Q
JBjiIljHE7/bQZCO8M5lce9XqCXIxdIV4S8Uodnbk2laWd6r/5oz5GlA/zDbSGTD
8GB4HqgUiG4oKsA7VdNSD3higr6SMpyYxo4L/wq5vvPxUMFKqfSzPg02A0puHy96
0DvvYTf/oG+GCZsAIIcJO9nkh+YcVDsaKGAlEwWkg7LQ2baxiROTvVWbKrBE9NqA
64ppWtzb9rCapgyej5rLdNwqZHIfxnppbb3u5c7N17N7D/fSEOh7cFhSTPasAv3C
gtOBZSE9wrdR5sFYLRDAH4S3+iJPo6i5Axx+pTo18fAo2ao46CCfxxoR6UHkcnYe
08NVe8AQe4KFUVwVn46dvuoekTRwrlUDT80KIiDoVv6QVecPBC8i4nEnxR7lg5wj
UAVFnjW0ql+2pHIRLGfVopxFItU5HX6hHncjSaSGF5u/TuYl+ll9wbp/oDHb/fnm
wVCgKagDqHLSy54ol6u7vXQuteFRC2bBAFpuAu4S7CEckoE+2Vc+VaPDtW/7N8wF
1C7G02nNAn+RcIRzDiA2sCachtTQuMCrROHnsUM7ZaKg8T9mzer5IfHVmGBtsKJH
+iKDABOgVPxhvRbyIqpjdRPN7mwyyPkJ6AxsCBUukuyW2H1sSdAmridstbrn6YI0
UPkDJORS9Y0beW9+dfLDJyay0eCsuJKhBoDdp6vBbpy7lNjir0qWPk3J8yCUK2CM
6P9NA64gfomRMxEsQbg9kHJTecWxW7btnyQAU0sh9oFeIad2+vcPC1mFyL+LSxu0
NItRNh8LOaxHDOV4hGqF9SHqQpVeGAk2UsT6Cu0Fpsml1mMf1VrvU9mQj2Sv/qKn
5p4gLx4qqKvba0uulOBbweqz+d11xvjvbLveZHhmucMMTRpMDnqZ2XlQnOUXYf4k
t5HxArx/3waTTXYXXc/WaBTM7gemy5wXUHPyBFS2zZeMgfwvTlZXkqfcHx+nS7Wa
tC0horIWswj/fpk4b8Xx5/JeWWXNc6STRSxtLDqJlvGra6XyFBSCBnqMvoGlgpnf
7FjiUxOCAf5vcrYmUf3R4pO+HgHZlHGrK2mM91r/ODHgngyKlZ3fR9lTqMVkFL8H
1+1Ij4NN1XPgigKRUT37lWsnNSlwtI/V6alXeB3xUTUdhlUiOGvc3c0WCRNl5Keh
IKB4TJd+0s0kCwMclM0Wuxx5lk+6y2jsukaqS8aaRM2H19l0FdM4wOyF14AHmkLH
E2RK/mo56KzAUX02Cj6+Cd3xxZ9PzRPTCNM0YaKTnqNbVn6be4Sj37pdu6jjJBvn
0x3X0uxcqD3QAkFgoV75M/CHLOcO3UyWby42suJFyIP9qXIGgxU7yqnDwPKItonX
6uk4BzLmejL25iNYhWOb8n2l1tTQSXSK3gsWf4Z0v7plP3GvumsH2/f6ZWaBbzln
lIpKKCKicuJy00J+g/U5ltaP6FeTQofWJHJuRyK96TZ8kdgMT7hhDx6d7kz4JE5p
43009+MpcvS0qLceRZP82kZPIi2Yni7KGY5n+c7DK2zS+VTuVGSGtC0FOQuv8hi7
xwYwxs4OVgpbpy9O08HHfaPBCfDxyMmd272ST9OQ3FPK5hmKFXNWLa2E+iWY6WVs
VmDMI7J83Z4AFvUBvE3slDlkZsk8QuQJxnMKh4VcKU/FIIyObK54b/jx8JJLzFvA
zes5rW88ffheg9nMcktjYOgUiG2tqMsKfK4jMStYt6Cbh7EtxZ2F5nXs7ZbBzJre
eAYrFKnBKUwkly2AFpmRDfhE2bwJ7cLxFgbfRyy4uugo0j5AEpxydBYiLe2tq4Ji
QguTHQgsN8lE5mO2BKt3Kah6OkUTF/wnbvM0s+6fZPGHEHCWZA0taRJBljj4dYLs
TVIxw7eBqayfZbnt72M04lAY9I+46oWK/JgDXtSTMLR3CYNRZoUTu9y0UvYaWZ99
Zc2iRr7z76k+BmUfiRH5NTIUt9zU+SnZHIbBHT6QqY/qMydqtyXO6DCXYvOayDEt
dLTKgy4sR1cb0vKwDD/ilutRRhwwe+Xge1vTAzuFOKusOfnNeoXMpoq7snnWYg1Y
jrWO57QusQOCM28jcTj5echzOI3J2DREMyIEQsz7A3baopiD4piWM2uDpm5OgoKN
IzjEvact8D2B7kp8YZxN4LrDm0JlcUKDQFIJkDR6c5FeU4+aKSVzG6XC28E+oW2Q
+1nsGUo9QgHcAOEEpuFDESb7dbzc7NOvoquch7OQ+jF5klRIy9qMKzAFx48f3N88
ZlOa1ELdJ/jztNgMUFfSIv7VPYgKeJE9hQUYBccDRjjPkQF1+TvVx6U/r2jYz0kC
554Xqpk3jyaxXUIWPmHqJlq0fHJM9YPaXloFweFAaKH0ExlQ1EqJpuyylwPOiVXJ
qJLwL23uVm6nTU+HFP6Lgfy6xA33AEcUEgh7Zk1uHPDZs+7HWoOat8z6cr9DT4Z3
Mjy1nEnYFSgZ6nfHMOPDFbe1ktN7Mcx2HfwWo02xU9YJDFDFhhrn8LrY3t1Q0tnL
fbYmgXBunGwn3t4pAGn2ZyFZqBHfKsKWoXC3uVOKIR/T5GeLX9u4+dtoX7ZeMEaJ
RoBkptQFtemDzuzyzDOINwhEx6a8XW+Xu2q1bPxrlQKI95P0gqlAgAinMAZXfXIY
aWQSNDqu8X6h9jwgh2ff+0IDuqPrN80j20Lyl1d1Vhk8TZcfOzGqN7IXnWup4jmw
kjIidVyJzkYiMvfHz0zy4eRo+ieatM/e/Aaf7Yu6Bsfdx1BMzQ3GQa/n6sspKI0p
yG4V/8KFcZmYcyZKbsEUJMkkRBRfGTveWh3LuukeTymHtiDpY3081W70JS7jfcD3
7MDcumDagIucXAPkhf/u9QtngIle7OKlEpYfsrXKjb8M+Ncbtt+e4WXDYSxUDXtg
QHdhdkmNu66y6E+xgIPeqOqNKB53+X4pxsyPaladK9L3plDf9mQsBZID1bRz+zNX
slfRKnDb2f+1a0vjLg3+Z1tTYAjIsAYHTKib2LsdqauTRIpgWl/yCC8EwbJTlwbo
pMMiruDDfxYz2kvYq49XsqpFzbBIotyyjvG4L5Lo3NFY9xJidfZmG3Rs7Q0BGCwi
lHbrFGAxu3lhICZPiFlHElTfYUkAlYCHRNbwqiRj0G/bs1dC5Jdfv8wPjncp1ik6
9l0YUltmWvEgxIBILv2bMlv4aP72tQgjsoEoIZ75qK3icD3YlRjbXVHwzrZpB3Sh
4TaZTwXQlgPXMzzxEZkl8rx1xCeZ7jIJJ9OCkTeCGOu2IoKrbrvLLPv3InNXH9Tj
uDzAjw64lk/OGUUDVz7w2EtBx3QqLyPuyonIgddtj1qUdSFQSNHcW9W1ajdxlEbR
Nf0tdYlGio1mW/wHwSUgh+uCbvT5F8DtSGqvEjSigAzdTCTOc6caBmiwSiJM8EYs
X2KRZXjFSnoLnnTQBwAEpHpf0GxZ2mcXWOLYZUIedHgH+7+TUcILEBtR0nVt1jIl
+rXh6sxH1im4h1bBRf8zgrQe+ooKECLvznMlnpFqCXDI6y7wzFMvH/X7MtbzK1RD
lMzS/i3C9Em8JzjtmhIhDafI6uJfap8cUa+lhbH6y1ESNES77/MpgyT4tGJZ0g2F
bPmenxH0H3Sa3a67+c5Oc4a53TE9Ysfg0Jn2gztjC0ELUKWn5TnlE3HzSyGFghHa
XHQ5m98cr2zVBdS9q7kBY1Zf1iVOlxvon9LaNxc5aJsHDdTiGw8jvytS8xp7Ys5s
5l83GIuhN9bXglQXU3skYA/QuH2LRWpz8BDPZkKdEVZDV2o8kebeaCFoYrXs+gFb
Tr0VO1ng6Ws4KAMvxo3ukgSzmtyB3VTw2uwJHZ7xGNoHoWVA8yw0p6bGEZS0RYq7
n9HgKX6FEALjqmqCDALhx6I/E7mcUeF4S4LugviUDZ3MKHL3SIts9EqUpmNrBT3b
PdEVcqQ5kWDzLyR0J+ZApDCQyY51uDNVYW6CfqXaQCiMufcoEVgdTQ94XJxnwrCt
GsZfCnyR9Ko5LY50q2O9a08Knyqjv6rtRLP8rsVjD+TbOTNO/4x3q4prT1l2zYKr
HzVoE4cuUQn95z4Tiock+iHOTA1Li44e6ytOvAlRL+jMQsYNtTb3zIwbJiZLW+fn
2puQR/S8DEUUDWXNTxYAxVxi3x8oVWqSmgswVAPFYcsGcUcQ5xK9z1aO4SolZT3m
V2KKd2lZ6Znx+ssrsOmyPz5KSAdqq14/N2IyePGfhMG1sZxa8oLnZDY7cTop66K+
w8+ZdOQEtnDOgSQ6ZNJMucph3n2xslmjnCmmPj48/vID1mEaqEMOHbrNpRoQfKzr
aEOSWXeSEPhrUpZL9/AtX/k/mopCKBKXcwF4M3uHJO3hM8qZGe49X7uygUwDGbXB
RjqMidHIrcbBAyGN9PkWjKccBHFjkF7c8yCLuAGqK7cWJYHZ8h+O7l3kKaMEdCtW
9I/boHS9NSKozZI/BZ6ZuKaMduLO7EWj/0tapTL8yybe94JZSRZCdbQBjSLDGGVg
ZagBUapURUDGwM4d4sjn85zItSLBxZm3W2zaoHxbAlGTP+zDNhPr61R/hPQUaciD
kg4z83GrjTa3LQ93OfU0IwS/Y7wjw2u7fZQb1hnwu/405+qf1DS0QFlBPU85dTCP
EYjTICPpgS92N09Efsf4ayi6KpswUlBXfPOdXR8TQkZD8k7gFB1Jkf8D4FFRvyha
MnsSamQJcdbiUHaNEzbDBcan6TBv9hhF7VPxRxaKJjCIRnZ/IO37gKGjGZw460Pw
sDo6aBZL1mMonwNxQvKBBnMC7s11OdifittY6z+ZoKC3rZ99tVcvROPA3/C0IlT1
0rEwYPvBnA7p/274vt89wckyxmkN3kwIcy5WDqRrTn2AuE7q2KNi/atjghFuckvv
vFuhau3ySK6wsVgFNuTMwRTfKKv/5xHVhdEGaYuORvtHPrnExwbaT0lOpgJybps4
2YEsn+ynOPaPzLiZs4bkHTMuicopILExcgMsq0Z9Ys6AMcuovjo1jkxVaLnxH31k
ZoI76T99hSHjuN7ASH4GangitckRly3dWKKAq1D+AQZs4ii22+bVbY7rFTqULIyh
th/3We0vYwDkPPUfbanXbKIcvvB4SIoZXxF98H6BrmJnR5sJ4hhCLQPaFKetxKqc
gbyrKDOhhyOKEK9rgP/y5AmyvC8VO+ngJdl9B5yO1TlNxRFyb8U6FyDX65S/Wt/3
QzFuS7AXyMWK5CHBh766iUuEXW57swGNx2sHV9mJx5W8bL8ru50eF0gcKIvorVol
UEfUlituOI7kMUxjCKiQbMar+BWa9w9L2kC3zOVtJ6mQYvGh1VKUFSEZ7TgnDsTO
yf/jgZM2LnkWIikKFBCFB7An8JaexKJ8c6Ejsn2fU90V2UsLMw3eUGHgMncNaTRb
YFcoOj+U4QMws5QU7e/dmtzghV/VzqWnxQyUPotKxdU64896LZg1H+hwz1z7JQ+z
jM9lIjhj80AmD1LLclh82A0MfqSIX4RPBTsP62VZAKOd9HdHQcliq4xtWcdR4Ak+
FE1g7JNqSTvpsIMfSxPEpV0S7CY6yNv3Gd5Yx9UwVlFDn7DmWbf5djVzm0NfEK1b
6PAaIABbkJLlINFtIxEC4xXLDEvLPooizBSopICdKR+QWPR99rwgdIFaD9UEa8pJ
2sNeK+4FutEN1Elw6MviIzaQ1UyQkY4+TCXiNixyCw6wguEfGd01ozO/udQ2MJIj
7tMc9OxI07iEcy2IVNkZaQvl9vJUBMV9A2zmpurYelu/dsjwUtAwir7CLLwbiOtC
SPC5H6TTwD6rNC1hN0MT6vr4gJGuAcnruJ1BbzKdAz8tdgH9ScC0oCLzuta/MRlb
1fAXzkM+j9nZ6P48NeBjoK7FVFVveonCrSxWs082rsDIiK6V8zwgT9lx7kOZkKc4
YBXYsewo9mIGg9C+9xqSqEnZWaS8gHMA0Ejr5mnwf+lfHQArPdyqv6wc0eSwF+1y
yS+TqmLHK2fxdeUDoba9BDSJbDMVBVqnq7bdxYdgwUd4tTrazsARVOTM1yJXMQ2d
4iDAHBMGuG2nBb0fLcq6ERHa72niX/zoz0fZW+z9/SXA1t7j+FJmw9AAozRW87Ij
M8TvHXEseHp4k32aRUL/JArnd/wPSGsJLKbqIqL3EOPxKSFpJP4h4bq6YLTGCChn
u62zc0Zw98KPH/9DL8okLPRuR3DQws14WyGscvfzrLU+lpDoAzoqm8thxEoXZG+h
edu2xQ+kazgCuRTij5QMcTCXTlea69Jt3mvVtf8DekoJtzcMsZjydk9rqvO2vYxh
jWyBbEDHGpGdydpUGlDFWljaMRTpl8gisQv4pXkqrlfsKlPoVQLFVRwLhAR9r0iP
vg4I1Wo2uR7aAygsyozxal8AMr/PzulMjRxS7w6JaP51Tc+qw52JtDPx4v6J60t9
wZLqm3OD70L736dsxm8YGbXuuR77lWkCKJku8Ql708t1tHAc5s0LTrA7omN1e0G8
0dclXiU1qc1JxEdGqYI/GYyFjQYFZBartU9vf4xdfEebNXSENoYtPq2dfw2aAEZp
R38QKwpzTUcAU2qIPcCQQ8kRgnbfjauFioEAakiQVcxbjV5Rbsw/fGPdco4KJxpZ
qzjSQb5LER7Pg7s0g4t6pcZluHI9nog5Ce91EP1pmuOjWu/0aWeS3f/nGpKFtDy7
ZPuETee4OK+jTYHN/PiD+N2xOWWKtyR1ThqGPrZ1Rfe+YLoUtkqAkZutwUY95+Y6
YbP2iut/U1bABrCg7WHv8AIhcyzx9QJntOoEMQZeEoFbhvF4ltqc5gUgX8CdKzAm
Axy98XvF00B7bmPo0r1kX0nay8QNbBAcm0AuWl+uwBauecHWN7cCmuz53n5fnQql
LyZYO8A2STr1EDoT0X2h7ZmRJfZuC68rRB0FKk13Mi+v0a27gXZujcUQAM1n/vhj
C+4sEulPJRx2eITUmlwfWqIS0iXy9oAvjIVe61iBHV50Gn1eybBFVanKjzgu2TWd
vg7I5G1ulQJ01VqL9E2IAxJaF+CJb3bBE6Rvjwhv9tuZF1dM0eOZyOOMP8HQk3fu
ghrmUiYRs9JDSE5ywyr9Q7PxBUh5fgf+CnScHCK2YXy4PSBawBd2HiAoJz2zVkNb
4FZ6CrpCkWYUBeWsrJ15YupXhyzQUFH8egRSljQANUv2H/lS3Kv6MgnEBp8v3yTd
EPSe8qSDHVlBnFntUQLY9uVDe6uf3GhZohFtezPB4zKlJxntVPP+Bhwetb8NpEFK
TMMTQjl14iwuEFxbWRtR5guWRcdOns0fWj9FzeSWVaASFNllD7pzVrAos60L7zAl
r0tdIrnbu3jtMRSkot8H++L+I/G/rVZAx+AHQpCHl4jx7zGDJVENhD08N84ke7gM
5RmQ9JJ2J0C7CZiaWrrJCiWhnBSTARqdTumXhD1GdH267ehYTgKoSRi8ucpvOde1
3gTkw2sCLSG0n8E3p3eyYJSUIHsH+HsxlpvmOgX1kfWWyKSgFoc+3WVGCPhzuCKe
I23VoU4EdMjii55yJOzWLlQrSAiEvKfq3gRHJ3+0eEg2d4Qhq0qhYwFOCiIM3YNU
bfrAQOttOxQZOxggVRq0GlCRu7zlMqZ6N06UmRBnosnWzbVQWPnRLXdj3/GgpuCp
zkRStYuQeCWPLgdRmdB/IwuhlBFGZge7cXB48LjY0cTabdFD+eiFco7FQgOFa2I7
QIRwBAoiGznpdTCku5MSwVaehXnjqmScb0qf8BRCx3gAO5h+vvScH/zjEHIYYQD+
95KrgT/Eerh/ZBC2wnzSP0k8MWhMMGJolBj3HQuRyKFIVCearxa+vB4qim5jkXGP
hTwrwqZjxZDqDAsT02j2DPSomrWG9sZdVcWU5mNI0vCVboT3OoS65xLc9TLqVxlU
Wvol4YIcgM8c14imAu18tP5K4oDQ6XOoOL5q/3F7YrU8zVgwNuJhDPIQmKDo3J1+
1x6fsOgaOtC5CHPWoeE0ZhM+P9NbRgv8gKRmbNy2n2t1OWAlWn7sisIUIyAC3iWM
a9qGVUr2F3JHozTAZWbHCkYviElXQQ1RgE5eV8lzoFHRVD7XrA31L++YXc/NySxG
XizSqwJgk0ZrNKK2IexxHe923Q5g3er4WJlzl29Ax9ab1f3Qb3KGUxL0ElCA/anb
vF+Rt2c/vrWbr/U6SK+0cU+JF2ssS8AEvdUqU+0Wig7Rdrd3icorS+7KBR+nIaQT
/C1brGQSyzC9ZkxJap0NtZGGcViZqWKUEHtxcjziR11w7lVXO2dzO+PKs/pcjYWi
JRpqAlh06hoIWiFzTwNlU2f051f4ONYhfnD2Pa0kHqeA162DDzLSNY19aX3iCZm6
wG7YsDw2mNbjP9mGLEzg3Wl2zRwEKrMJGTBYHldfroJDTwSkJYjcDafTw7/M32dT
aUNMcqI6B/LVZts32H46ZKmQaoPi4QrNliZEYeUDmCpVW5gqobIerz0RmEx5Fbpi
H0aVRw1h1Var0B4yn2jzci97Ig+6IKLKo4PGuqJaGi2iTPjwfJdROeNMen7s5Pvv
pmVJfKPfFJwqbM3iXAAEtbmpexawSr9eM2eiK/ZzruvRDHy/QJy02aO7RmzVhDgp
WpQuhwPho3WGQwUUJMatHrmbJiQUmEnGAHsQJODX9P6MTqyq7x0KvL/AQZTXQ7y8
M3NtHCIWYaHFtONR6330ZIP2K4JPmy/999GyFP2YOxy4jKpqjh4R0v1c70NAKjLd
rWxggJvwir/92UqPHwhW0p9gSYXnVwPXg9da3tuGlaHhrr4AuILeuxCm96f8ICkW
9MAjSWUYD0mmc5tLpDmyxBASkBB9ivKJmN5HuuoVYWaQa+31l/Q5ahxjT64UeYfC
Kg2FgVBQdphzFuDix94sv7vdSUZQfXS4WqnccEjZqsJA1T+zjo9LlH+xEHw4IaC/
SGIjJvPgoQBslWnX+GqKm1ii+2fdHdsK+9mNOEvyK6axTq76/c9GAHuPsrhYhnvI
kB2Q+1E8Ll+vZnhEb3ABfA4x7k3+apUVsB1THLpmAwF2O1vQ7kZjNFeAhYi+LzSV
wCuVswugSP7XOtGyHjmPsI6kVpoWF3rID2i5Mm+GdSxKLnu1pWqXPDlu74l7Q2RV
gAeG5dHAShyho5RuL2qmEddkJHbUXzBcspVSAL0nNw2DlCrecOokKZg/VF5UdN8c
sAT7rZ9UD6dBwAODnRVUgJTcJE9BX2cLwIqa6qlFfLaxRoVO0u8cDE3ePcLlLmeY
adJG2h1ujyExB+765ypOL/WHFZYIYrDvmPl5rrQmqgUxdMvSkQfqArgWRNkD3bdj
z/qnC1XgnL+RIMSRw0/ySzj2sRpqv2cHgux6yRcuy/ZQXi87EgxzzH+82fac5ikU
YHXOt+5fbWcCWeqkMZxdLe6WZY+JXmyUaGH3T0patQMOJ4n6mybaZiVi3GmVj4Ab
/rX1wo8eSpNu7dqEg8zMzy0mUC8duwCDcqWBvCNWfBnb2xPs5dUZzZdgackhAY9G
fnEsQH5HHUsCmQ8N77Jsj4XFJ3MaUUJN+DqWtNqS+pRjZdqYxTn3pqfBPM3J89JM
ofi4q99+j09LL1x4lc1dpEa5QGhOA2lxAVHSmE+CyDszbDZOwwgQLvDVuY8lk1Tx
vGHxEzURv88+KFIThu8mnu5i2pnRqpFCgWug2bRtNs44w3zwJdSOPtRiHQ8OhaTU
4b6dK6rT/PbhUtHGjj2ZIcD4X55ZqU5PPyX67PDNbOlOlWKLXUAhhXNsAxFJ6mko
eQOwN/lJn3nWuTyKjloha7WYDie+fEpN6kD605xniVT1cOJar79ABXKIqsN83st3
cNEve47LHy5sZno82UzB8gJRMPYrIbvS2twPIEqeSQ4p1UC+Nw2F1uQQhmpUTkNF
ZEULg6BT+lDDHaPteV5tyZkjhLyLSfi6bzgTbDGXHpqC4hYRNfrthcz9thBg1p4Y
WeE2xS5IOmwlTfRTWr2yMz5mdT5DFRobGKIE+C4Aaflh1qRyS9Sp9vI7AtVYhgjE
KEyElUQ7bey9DD9Hbb4th6ShT7Dl3VRyJZe49l8aWbRWavHm/0DGwX2WjZALOMQX
YN6oABO0E/4JiPoRI2Rxmvey8mPJripTqFOWP1vHaHm9N82Xc2SngIfQ1tgw/5cu
S2YG1b0oPgRlU5ZqOQkPX659kr+ZPeRnk6zcq912WUU1RMwOT514gCUXO8jfG6WZ
FelIeeKrvs6cNcIZz9G8g77I7Vp+NmH2IQ3+H1CnM3SYX1C5QPLI2lE0P7SMqtjk
8ASStLupeKgKJ/ZVMajv6lwJRStpkWU+9hIgFd9djLHeswRwMCR3m92zT+0mltw2
nyRmRxxTw3nfJEyx07k9IUeLE8j4qsZuKz//W7EwdSUUqS9wxcYw8qUpxsaO2c4b
mPbfplGar/3jcUYJ8hPsx9H1hIDWY1d7rItVZNW0nR0kFK1Vl7pHV+TDk1T43/kO
BzC9f+8h9U2vr4gcY6w6JJkWq+Sbu2Lce5MwquTnG/OoARZyn+duL/S/6uclAkFP
Es61CnuFb1XPAThzYuLq76azBpOSD9TFBr5WqKDwhiWBBxMKGidpO2w4VdqRwQW1
5N4FHEt6j0dzj7U5VubChQxHGlgMl/0kwN/xOCiNuJuv9f33UUe6r0fWqjLKHhlE
0DaZ0Ddy7lJvjxQ+VZBbA3LETUQ8pu+ryCN6bEO6d8MNPrp7reYOlL6+OQzIb7OG
oEyecJ3LCVHFvHniB+GwBpelRNcq5r3KKAX3yCQPMKtSFl8lTB0IxDeBWdqqKhBN
w5/uJyVDvvIAXyvq9sGiBHIbQ+ZuK7FdVjbHuNh/gLzaZkz5WDGs2886z5MituMF
7N3LZQGLikBImwgVsi3Z7pBdwNyY0efz0P0A8Kq/HJDchyu9QBLPMIv2SCVFXOih
IfeKdhDe+HRzT990VBcuxCbORZc3LsAvMdPuChSFkOsnsVrY4c7l9nene0qd/wvX
KhqrGOkkwkrGlyxClEcuQHeRe1Xq5RLgb0QMlZTCj5aILwHfA6ji76M3rmkLg1gS
0Qab5rP7L7lvS6d2e/rbVXwsBzx2u3gXcK58yieoEPUtyV5gdaXAhsJ+rwn4Z63V
wh/zv4/FOfSc2bpP6Pdv67DEvWZ4z81EkIO0DJbCiF3ioSqvSKTWONXLOVAIrbAh
ghEfE2cGBYRlFQyn4U3LffMsNEsDxpIOCLMZggs5ys74rtURmIITUyl31vDrXGKM
Aw3i7+JQD1QC+8q8sYj3ZMIrAxrm8NbCAcjoCrEhXlnPJpVOK5imuMEA3zSjTx1e
UMIvez/oCldCGNQyPEyiUmzjmy0F+fn75m2eDYyoXK/o9abokyMprEanUIl+zmty
pyRv1PrGSWx69lnzspQYELeeZ9skzwaL+wciBFYbmUqrPd1CjPlobbhbWCnFpsut
NCDz09HFpI0paCYHN/fXTCgVYW+MIG4Fy0TZqLejQFqJwXdwBeHgLqVAlYVroZrH
+Zc7Bh+h3Ey56Pvk2hc/AhhSLKxAYPcxZz1+9Ojka74XIB3yRNTQK63wWwJ4Bifq
RXEBg3Lw5afsH1o1HCEnKTUYFfc+1hEDcq4zt8SU4lTPPT70JfXCHJ2ECmO3eJJz
s2/KIe7XYO5pxUEvOztqnA+74WGKsx8tirLgu2Sz/TEnQPx6DndUq4fTjfH7diKy
ay7fBhuKOV7L0V+KXNHtpbRoJnhRffn+0ENgPgsi4hVFUs4i7I+tVDGOEWcJP87Q
Y8PzSHVuY614PC1iOnlfvELgSZjO/9546dP4/cFbkw8ts5GhFMmncFrCxYlIoSQ4
R9Yn6Dkvl3aMnZtau1zJ8XFzgz+oV2bfEkvGM/WNWWtz/IRcfPDsIagCSv5y+Kst
YmlZos1QlylGCav00sd66Cafnv6sZMw+qc5n5loQbaIZ0iIH6DSGRM4WFDVPZSwX
b8FUG0BBnJOP8Bve2T3OXsrz8BJySjZ1Xs4zLgtxRjofEOo8y+jHbnpXRJnUxp21
62ftmI227nExP2n/NavYkceks1vDCpK9tUxTetkH9vq38k4KUqUDY8L/KOUFxI1r
ZG33+6AhDOSoNjI+MoTnoNNIClHRat0W8+k4L5560wAg4gKERYFQy6GHciPYIjlH
kWGfgULKImz8QEviUZlkpJ4LROji65/H2sa+yZIgnSqj8P+Y9UTaTooIPKOlttNU
TcbbMqU1cr6w4LFkx5NJ3YeOWzr5Iyd0Ae6Dz9L9m1uVGGLdi5SIjio9n8FzN1r6
yruF6wOQVQo3VeLXIjlvPF+vX+5g0nVCke2r7Uq/whDvBCEe88O27pJlpO/CJBsg
TObwcb9JI4pREsNmqGOUlQU0AAmV4i5gCJzOKjDJtBHbZ4Lom6V9Emub9MvEEzQm
vLniom1V8NKNST7ks+P8oOc2dqDLl6tLy+TdYUV/bmUIGqJLdHTBMVubsKokqwsY
t4lRAcYAtkKGApdxVsmso0DuDU4aKNvUjEcG06eH7oKglLdVsFxFYYV/6rVTo1Jt
uf+wJoHtq23vQfp6qWuueiP0cviI8SrtyOYJobJJP19ndByhoHbDWysmHT1ju0i6
Dyff9GqPQ4n2pBbyOt5HOT2lR+/XTkLxYBfJNXhWesOg4J1RoSj+SVXA9qDpnzVO
HwF9hPEUjs5hrr9d9WUovCLRceNLnsRhB89jw4Y8JceIpkJNjyaOybt3LhrhJUhD
LeP7G3neO/AYFXIRl5P8cGn6e5HsVT0p366VCS44yrvy9JGxIlp7Ahbi6GeM/HXO
7zzM60/NigWqDVO7hOzEzEvBVVGvZiLXLGekOIEso8qen0R+0pTe6/LfQbeNIagR
wDKUtf1rJ67bl4lwM3HHeYqGvZ5eWfzSqPQrTsDy53wzjA/gaSVtNk7QoUEVIKEt
MMlz+OU44fjN6zaYcVt25Rp397V9SZKxi9ZmQ4evzDtL6157cqSd6TL3t4Tk9oWp
MeiXmFr8xVPvi7rab1a+9WxPnb/Vb5VwSzf6MHKG2TlNxDTIm7eqB+r0oEvKToUl
EMC4fDOkUip8ijtun2Qto4ECPIrgHJImzsztT+R5Y79OX+ZcYlIeZg+UrnIkEA5d
fJr0aJ5FVxJjn4F3n0LaJviHuFUOAU/EINbkmXG4yPwW5LUo9qUGa4s7MDWTmXX1
DWuxBCgrW/hUTnP0elf5dU5AVD5bNu5ReS8khPPPndpshrAgm/wBByUBRmZ6dJve
8EMPUfTCw4MrPazyJcm+qgd15XHJD6Foosc9nKhOLE8zAsFO/q7pohe+V2ONXB8g
7US4E0yNCGO1PpPqj3OduMsZcRgxefEK92OERFjLaSinyreybuKcJaihyF9k8Plf
VrPG+2f56b5Sxvi05IV1P23ZA3pcSCB6g2+ge+h9YOyYcmotljJ0j8z0hP2Q1t4j
C3Ap8ZIDyzaGvXyiukjmhZud43588w0FwZO7dzN+/pDBxNRlCY/ALjSAnENCKkvk
YgweXGh1mOOPXfiwh5NXnKOBCMTwxTDNBJo+Dloi55xlZYpOA6CbHKKpAnk6FmoI
tVTUVv3e+SXNblATsPcDshCYYiG+VVlMpivIkzOoRNgLLnyyQIRH4u3ZomrIbVp0
moW3ePoiRXSdMKp8FCNf3I40GVWheJC2FyTtjic7PbCmQgV9g/8wwyBidlkj06sx
ARL7zLY8K0UWia32obZuBuqRPS+FpTCX2jAITkUrLaKMifH1a2+Txoe3JyO5Q+oM
nCBmCBJsKfDheu1Z+MAz8RR8avtWOTOAIx3VGIoF0kRM+PRoJ1Ox+H3gHF26ZeLT
vcKbtogky3UnRb60j3yrbdsrKvIlxKuEwAMvs8D2CHttKmHW8ad5Z/lTH9xqZGrH
5WD1V549TYy4keIIYlyUlpWriPubhkZ0lNl+kmv65dTDK/ZxIFiS64d+Va4vj+3A
oTE6E7+DQuqGXMjv/XPV7hJHcDitRD1tVQ4WwAo2XJuttGg9jZkem2a39iZYnnCX
O33+/GNaW56BMuqAN1yQgOj5HCZb4djet1pXo5hOUjTTeUSb13ao+CP1pTSlhxaf
dlgPaorrdXepZFx97vOgot3lqPbmECETEfe2tK5pfLd6hLPw20YyDwE/2LIVeHJc
fgGYlQVg74jm0st1Zdf0Zwu+6TvS8Fjy0aDTRiQlzho5rY9QZUus6wSsMnUJ6a4v
ECk4AZ0+rAtn2cNUGV7bFqmdphiLb4DROY66p7eBazMY9yJmrueM/8oKfhzejrlt
p7mQhHR9dcHcaYwOaaDj8Qvy3JRPtATOGBx61e6eH37EeyDhcuW4QJoELqU3IADe
aEvd5H+e7TMRJHPizJM8oOQu2eUU8GWFOWQ8pFXC6QuYuSck1bmwv0plIx+wl25j
v1iUEYwo4tONE0/kta0hnATOjMwnvo7XR4pqstys1QMIsXftkDeFkgjI6HnR1uaF
4oUKe9QNey6IxXa7N1OmX5uMh3dmJxTG4NQGQ9Jpf1eI9r74MbgwVFOSyBKUpkLd
JFRDrc54+lMqF7Sh8OMcZVxpHQDFPOH5oyCH0oVi1YXYK2Wp0E82nH8pfk5gr2JT
wdFHlTd2jHP3xB3tbqqRPjbaYfk3MC8+xJ0qP5YVziJbesrlZXmuMG1ifq8jXe4X
peaZfcOLwxr6VFtEu+rlM7BYFn0peGQGmC1jOt/qtt/t7ev6wR6wxAHAwfql21Ec
hMNTBoFOUFsTvzt1x6jlvG7tCtyME3PFEsNDoneFRhbdJIxJT8ugBRDdiC5Q6nt9
ea4UYBbC6ZkZtgh10f5L0fWTgmS6YyeW8vc1z9LUVs5HqL8FYXvh2xokAxLtg97z
jAfK1IxiX6TMKkUCYvnHuLMKa4eYt5wN8Gl0VQDIg7DtV9tpG8rFKLI3jORJdnhZ
IIXxMzmjhXMMIxSwZNOpa2/h+ZUrwYWDmCwLh9MT+Bi7oCLNmnuj7X7gFDcyl+Ul
04D3Ul8btrogemQ0CUgCJnFJsmYqZLnxQN5RTaFf8qu3b7wAUUXz5vHVH0LuCSAn
maeVNqCeHQzgGzayQws53utyqZYP2ANAXpeIfb6YHH8dgqr5n7AYfUeJYBGP7gpj
twTOYyXbCPTC08a/5AAwrABk5xqkBCifGsiDl+ni6BGvWRoahiiOrPPeijH14dtv
h0e+j+C/fDj+7tr9XFOAZXJB7sCdRBnH6Ac9xF2/FJnhz8uzCCOwi4wCJ10WWvtS
j5HEFsz5XI7mhey1axW9rP8ArElfN/ctSTadUF5LfUavAe4FSEgn+7iF7RxmWol2
9YFQOAsEvnDuyEi/WSiC8y2QuoAGYgKkoqtBF25TzUq1rC9DIYAT9bm5Lnknz2oW
VeuTooMrB+ZoI985ZrrPigP8ntFfOYg5Z6Bqg6ifO0FLAzRG0jdc4D8QBD2DSrt5
SXjiDVS+U51k7kE3DqPB8WtPw0zuDFomXO4qO0W0O6o5ULKxXMFp9RpqueNw2gKf
RMzRfsZqk9vOgeD0HTR1vwlHVZ6uVoqzUSlTb9oVLv5wDhBrNa27vCUjYnEz27rM
cXY8fC34T7S1/on/TVLvFvUGkFsLRRrFbMzZN4BR+veBY+jRlpO/Qvl3l7c1RY3x
JyIcXJERnt8lwvq9AoQCBak9AdouwEgF5qlNFkpgJdNEQlvy9csc0+7SB/Y6PQQy
TaBmVT0sVILj1tHbjok6IYQ8tIO9jleXxbgzvoMoRevezJID/jfE25mENb20ZPaE
YqGoftODM5V+1anJA4dLJrAqwHMjQ6n6wJKMa2gy0xDLYGrIdbj324W8a+VWPY5L
Igvb6h7lSQWrTDDWP5ywCsC37/hABRgoMWLfMMTNLQ3OaGA383QuLtJLycepB9CL
mU+LEpw7IZe2O8cnRX78CiXmaq6sFyhGedqjDB54xAZNExOXLK89tGWXBcR1QOnG
Ym3u7aah5vCYusVoVMe/XpshLwYYhwBAr23GHkfWIDNsGtVk0tLPP9AXFxpKS+UI
gofbxePMmP85mJ97T8F8pF/U1nK2A/mIYf3QCcyKWs4YDIAEVqdPkUPTkvZWuBUR
tUpJ2c4mhGL1nKqSEi8nIPbFjVVL/MEOOGD2BlT+pKWOHgHsBBWOFrQ8O52jp3jo
HVfSN+iGsMnwOp042JblsKVh9Jw9iaj4/es6JfIkD1RWpJZnwlgJNcIkL1MSP/hp
kQlMdWIfYLL8c3MiJuQFfBw07rK3xNF1IT+w+jg1VI4AZUC/R3EEv6ERN+OThfYo
x9HiZTMJrZKvJM+EzCKo6jiPqqp9s8hEBxknZtkQa0EUhhL17rvrbAo/PXAWs8RL
rF3Jmdr6VdPqfpJH0OaUCmrIqCxRNiljB/+A2dsHCNZMr4hYCVp+8r4FMshv4MoV
deTlksvYSh2rQzwZzvBXkzK2Pn3qBCKXEtV3F3pYS2kfVnYQXjIpICucjt2oJa3Z
acCjNEfqglFRiExX7EX6KkUIWPry9YpwbELumcNjDBZftvSa3xn2pamrjTjF15L3
dQetG0zZ9QxcYHRFECkRKDoMwf04z/np+qpvMg9FExX6ON3lH6w5+P6NcOLHn99x
PIrtMPNe7mOZ8IgsSGD61EjV1mYTGLk0vLpJwaCbLhyEESLmp+lORJeyB7Kfnpdb
2VhdGvEIJLLiKvHoEQAikcNjIMj9QWIIOUKIY1vfsIeY8nVV5CD8P+MCAhz4M584
Kvyaiyp070FpK4Pj73ReW3i58V8zUvpPZlgld7c1u9L3djY6rD6Bg3wLfltNzKDo
EKDTqaOxEfoIFTe1TTAuZsodsmpMYkDK8wLkQxyepTbKcQEUftdItDj3xt7nEQc0
1bRgzk/5YF+hffN2yW/E5F0Pi+TlVIN7GOpbxo8TLKT8jphAyO4GhAlZFMwX+OhG
VZL/NejqSb3auE78SYxsxIyewaO9Fy753sNqok6XyqGYKpQyEvIo1xSNX/DhJ2Gx
WHFTvVXRa/gouEpNthuDq1tmhx3250fCSZvMrdi/65k3en8lbb54B4Gjj1kA3VQ5
VZ1K+0inmoFUAmc6GEIQs5N1cS82Z34Gw8QiLYwoQDtykowewJlYX87JA3niK0dY
JC7Va+hxbhcxHQHCGafd+d4AGB/+fGEdPOv1RMNGcNoHEzcBAR1hAMhfRBq5y2kZ
PMVIvJeqs5mzn5IDZPbEESNANw1VXXYQYXruuucW3NGCYLz4HX6jpTutdOkaiEJO
F5I+poXtbbsfkl6U6PhU3PCPQ1IWQqzYOi26DC7wycVQ+Ezwq/OjGj5819KiousS
sxCebCfzK+8Nsr3fp+2+yo0FRW4lL9cmbrrVRa2CpzjLN/GlAXax56UKldKK8WBj
ik+GJLk0EW9VsVPSQJaoXYBncuRbK+o5vAzuQtPqeHLAj0Zv7RyZ44gPWEQdvXY/
yfVcxlW/t9kESp1oCs6oJhHn3sTaXAkPCtEya5SyujsTowP/cXwBBN53RWgzw4jq
8WOCRK9VAoUsaq+ns1gJIx3RTulhqTo0vKru9JKX9T9003YxLZGkdL5aP0zWN7il
nL4QVVzK0/SLpBbSvLk0MX50gKK4u3Dby9cvciS0s+rx/2uZNxuFLJfbiaPB54NU
r4k79eham+eDZbrXvc3XZ8aXG3CfW0PtSO80qBsj592P+LFt/c8RC9xulc/Kr9VM
XBg4jeQ8KEdEvC59vunSN8EyYO7WATtZxrkWtTzYw2o7TGh2TniUOsNE6sf4Ih9/
aKSBmKxRxBeEbbqkwovT9UfIByffp1b/c451Omb0uEuOd1vEwDiaJ6QE97LoWcD7
+QEwRwSGp7KpxT+8VNbYrWeMZWRYWipVADDPWwgKHI3rGYDkLLE0O2tid9jE7ixP
/IV2Vg/P4moKug/grhZy6nbxlrR6psfojWIWXZmn0Y+95AvtPbbeuPZsh64WsFYy
qJs8tPqK3KMEpDHqz4ibQsRMgyc4sHkfVT05JGbO95qJ8vju1z2ZZXxf4G0Whdhx
VtiZ6K9ElF+su0Z4kGJSTwQ0NOVkImYE6Y3PgSAw//WFF1GcISQ7wvWqS7EZvOtC
EqS2lHF9WpTps6R5hagTqsQ1zKU7wOvRENVYzcKyK9TkNyJrlAPDUp5msONdk3Hn
g1yIFdwwN/kA18onQg2WgtptLzU2RttmGK4pJXbmhis86A0yCwqIhB1KACvUc2oI
28nwxLxaXG8FNr2YCltpzg+Cwqpsz7y69xIVxy0N7ot/Tr3yB2Md9JZfm3bdST3u
KGHQlQcKVYUFw/H7XOn1W4XZTN9RYxiXgk+WSWN60JDbKcy40tp9yXsCeSJsQp/w
HmAuDRO1eAZ1hUDE6v2HjfRPUrr9gSEZNxphagIbnQMMojDgxAk2f2FP97qPsg64
uLqcsBna86nUTDLUgE1OXjHnY2cbpWaJ4r6VXVc00kYmCFIhUVopxAUj9IyfOEOQ
6Xl+fp8i2UBv0L0W8XneoLLVwLZLiNM75jFk0RGpYttReVNzgI2WFVbZwg22eC2n
VgDuv3ig0MneC7Q+oqAbu5dnlXhV//3AZSZdpIBGPRlq54Yc9u5z0KJHuWEeW0Mr
5CknW1LAS/n49BFF6F96dRIruGIzHJ3URzR4tVqrFsR+tkoLBybj9mDMuGnnCDZN
9dmL4dynf+pqwsPTen6P3mec22aD1+tdtnNZuQdLXPStxJx9/RHK3n8J2GOcP7ej
Glhs+HlK58q6T6CuPJc2qXAfOEkZJUwbw1SUScGO821m/5aTM2ajImIawU/u8Aiy
Ar0fphejiLY6rex3Et4dEVsETdZ4p7QRiuU4KbKY1qw235wUUBLWbSAPK9zzipil
eHhHZ9DiGKrrFWgCpP3/O/g5zYU7nujLZ8/1y7te7+IAZJZqfJT5Cx10Cd/tUeJe
29T4WLZeq6ng9WihEE3jrOTYOduLmT20WZl9tQRBK+Gq5iPyqlbEDnLiVTime9vw
5Va8k7yfEckcVlRasGWDcR57AJ6PA6MHYz99n2WvbspkdioyOC9wnrRcBkXbEIwC
HXhh5H87JYneldkrlFTGaHnt4OZb8h5oBH2E/futalEjBRjtPXxSvBKXJ01ODRFM
/u9zA+q6G9g7u7d7oWO7AFPJO99aOvjtn+cy4w2IPbrJYsgj4SgsoDfQigchQu1/
RzVlbVqo6EzbATtbPsLErnMjkD4SOEhn/T6WLed/va9XFTGst9a+22z3WsRmynYB
20/ZEnkUW5+JFKS7HWzZfEBSX2hw5136oLfWn2mtVUaI+seYeA5AQymbR8NCocgu
YfLjZZ6atC3waJkyDVrbx91EASE8C8qVbSjVhD1YZkHVO5//RDmE7UjCHX/dOkJv
0xPmxMWteLmOvzZc7GKT1anBGvoXYFqnATFgmpdtjpI9vQxQ8N1KCJt1kRfTI70K
hj7Skkivp5tx2HYCYr+hT5lruwcCbeVTUQoUqkxTtWAj1GMOrLdE9JO1j6k+SrTw
nez0jRnga5KNXoSxla8PO7e3lBUx4KQCO7totwrzBIe9sOe1xyC0frHnoeQntpm6
2r904kags1x8jzVLWTTngGD2q57ap1BbT+QH3UvLEjvkFhJi6qFpuvxzkbh0lpzl
xAEc2UK+H/HjcsMTbktROOSGAV7GeMPqiqc60P7mEn061hjsmaH8iEY3BYKZiIzD
A2lYo977zlETwteUIZt93COJ7OMAZxl9DIqlL+UZZDxpGIbusdMpDKqtakyL5WpH
1Nd7/tSZMtCXBRkeKa2KqHY+3TUoOSQvfRWX2K4fww1PpFIWRG8Sz6GMVvLuN9Gt
fPUs2puDqL6LCTs8It69ZGIf3rQ3/sOY7xETXPpY1tNgmoKdtr3vYxjFu7ESSLH5
v78+xsyC7qmev8lVbFoy8wuvwzx83RR7c9KLi76ifWOauvOMbIWjyNOPgtoScFbP
biOiY3hWssBDp/UeTDYVfXWi7i4LebhL40SXYrJUnpheKHkYaQ4JpBwtgxVO74OW
WVl1reW+F0M9JyacIfH9yGN7FrYtV/PBeU0JvXVhX4/PqbhRHnpQdfMufNrHGWlw
9xQky/ByshYCCMVmO0Rn/btF5M34GnNWakJlVBi9Z/6tnUI3Z9ezmNmeRn1Ii9Nq
PsC5NpDg75ErupsKppFcxY6A4AzMyrkErXRvinxrpckjF/pRKlUmrBczF6dcxzvU
F/q/s87bN3IYKEI0TF7bk4+laTVCs+X1pCbWCGqRXI5n6zyjEq14QOrwqCIk5N6Q
ueMQ43LGm/mtDts0ioXV6i41qKcGN94ydbch8fSQ+QO+tR3hOTOhGK+gsLUxKvYq
0vZPIuEJlXYl4eckcyGgMw8EmGPUiBej5wW63+uDymLr71+AfXg9jMDMQ66IKWFF
jPj8vWQeoBnECqe7PAGO4/89xIs+teb06Ejfi5PTZV8swoTIrz4Uh3HGD02VhOOi
aDjBZUAUyn3ZxLdSVlqCkTiyZ+BYc/xa6cJlcOKSbQxq8eDvTjg28Ps5qygzQyGS
raP8/xztyKXJu+hgbY4kzCogy1YhooOdm2BnNkSBl20eg5/eRBV40jsakfDmvPXl
AM6mQOGghII6I9k5JeBJET0AHWTiDu2RU4sksI5FUhMhdEAlEI53UbRDWkO4z1ts
/zfMB64vXy44UcE/4u7kdVNm24wEgN3LyUeq4rC9/4pu4v3j3C799ETsvXQXosx8
wzYi2qJNtpCu2DWP8Q3Q9VJlSMDgttD8W+j4FKCCOjkg0MEIp1Qlog0p7csRV/3I
4w9sCsBkyxF9M2vgVGKBSszcJ/1kYXxUPEZA7KIqsC3LEadhQUUCTH4+PrajQtN2
mXOtAydDnsyS+qiYfNkJHLENDazAE3FW2I+f5LclKcnyguZZXu1oS3zM2SxhXGrp
alKTPQ0dAu9Gz0tixVswoK45OIVkAMc6D2CJfcN49/Kik0QWu8aBRoo5NadkHvxk
rbnNq3r6bxbwO37DXhAZmWeaRHt7hnNoxjRwB7CoFfB9CD37P12oZMiAN+1CeYOU
Z5ds0oYlcj6NTR7cF7cwXJDs40TZOjUO3E+7xG4zNlA9MPiFL2NUcOwdwOOUQXZw
qh5EcrI+ibJtfpsI4C9Deag3FKeXb8R6AV5Q5mU/4G490iyOcs+eVOd23gz8vPUn
RAfG9bHMQPh77QwKYWCXvNE5c1DylIDSGqk2LvL7V7dQDZHi6hK4+6X/QM1iAJov
ayEi1tJ7pXFeObw9wPRRrK0JHSMN9Njs2cu/2PkRs7S7yNZOWiWMCAasoIdUJGkA
UC6ubQcHR4jcN1kXf2RuyhG9tu2T6vJ1kotkkBHoAA7ABQe7sWK1pzYRvC9fNWix
zyPnBBaf3ACB0+EsXOAmpOU0jC7lkrEutj8HNPkwiv7QJVIASQoLQYeVDFiTh2+T
UhSbjF1376yDuL4Q795Fs8EFJkgqspvQLpmm+PWSR9TAa71mt2pIG6YLni48Vzuh
un75Cmrv5wKRkMVWZlTI/4rGfRYZGHQ7gDYt1MwfT6+m7zOCG0+dziLcJiQ25KOe
PBymjh3vqBiyEptZka3K5jYPsbCZf1IRcmCia9W1TU/k304ZZO6TarMl499GVr1n
Wm1b14tpTGnh/A3wSxKnsQfv+HMAzhrllxdY3fbF0gesS1k8YkQyd4Ql7pmvkOTT
7YBWnRPTx2mszRFKHBknsUM2zrZhhcpiyeYX+T08QmY9CAne3xpsBvme/h8065Lf
6sqeV+ictuTvQIcMNL46lXd8++BVb7uH1QjM156O0qRi8wM1oNN+P7PKugMQgAvD
SR0Hbs2AERD1VMibX5XkcinCSwgvFIK2g7zbQ4GTmflNHRj4l3+QGYq8l73qAw2h
be8NLErM5Ceht+giGe78TdfpXXQL+/WccKwJGZiPWoLAmccj+5Q7nYyDvLfT8x51
hXJa0G8IpUHjt5f5K+L8aSLdmPCeZ5zOiKcqHG5pLNyg9vIToJMjxXeZDD4lB/3Q
ID7nJfm9sd6JjZrdfxza5oEJaKj0gCuglPuL+T781TMR542HZRiYdNIbS1AGEX5r
riT99vnyIh9GrGjYem2XSNpukhd48Aq42vaJ0hJkkquy10hsLEUspqYiaB529dao
rOVzPoz9pf30QojbgJeMvCiNpvKESIKJZ0mwO7xgpyxwgY/k3rkzlNJXmrZyIHG/
BQlbb6v/2U6nsjNjCMdvDvgcd1PrbtjLeCHHG23mmbkP8m5KIMdMserN/lnVjxpz
5Z8lKrTC5C14vi97pxlqUd2Ldv4LLlOjOqbYe5Pd+/nazxZCBjPEQXGmess7p+Y5
IL/p784VO3lp8TV/kvXLXm7Lqjm9X89soUp/QznnX/QINk1IM0Vtl8tDgcv+Fjoi
gOrBfFgEmb32pkRdMkh0WxhsxV2nSBFoQhdezYWp5P3x9+HrgeFqrQecYYbSQiCc
rWbBTuJixdHurVl07lz3ll3SIu9sxP5q79Hucqt8LiUxBAsKJ+zhHuGDzOLu1ZdG
qASFM9C4KKfYjQaA+Sud5siD8zXM0BRliIHGZs7UK6hjaIcO5PcNxz28AWJ+IjAK
xwhE9LmKJxBHntWoip9SMak70IAiTMpI0iQ4cD6Xr/azyDa7iQl2Nn3sdtJgnOJ6
WNQ+3MrChmT/wMNi2zNi/M5p9pxRmQ6+xKdQdLh9cbXOUIlS5WGzfSC07DmoUeUb
rzxZnn55D7YRtA3O5HAAb6urgzmAj7YWigUZpDuNSBscfvXIG1CzJ/FoUMfE2V1R
cj9Um85xSUMiHF7gQ2HVmRaSMWVZaXCn6sMV1WZlC33EMbdDoHxPiWrt0S9TMcV8
m1DgIQaw15WFzi6ILG2B86Ys9e/u5PMmJ3Ivzp5WaZ1iFRsDr0mobO5XCD+6ZY0T
lDjOpTrH3MoQoZcYh+7St8gjp0wKGZPV5qC1p7CrwzY+dbSYnTDpOskdHMr2xyx7
+ye5DalGBmLy9aZ/9cc+SGOoWiEAvGsFOvED/mPyZWEDhqm4iRxUuT+zmx5sQOpl
tp4rk89PrIJWvIBNPTVWCmksi9g2b5KtdglwGNN17XRbjrm+evM3EZsTiePFf+ox
gUD5L32+oIF5OC55MSDE7amAZnIwi8LN9XAvcFIhiU4LJDi5xDRqiUaYreou16T+
/vtAhveQ1xz5Ua3Ys7QnapOBWH15+U9kPJyFYK08smu7Vl7XdHWkMw0eerXRLqpx
pY1QsAxiH2mkjDppglME0ihaoyaZ/mOdAcKzjJsdbmDvkaIeUNXpLbQD2VIL8sup
J+9MQajEppKmj0rZNLrgLEvE0Uoh6IM3/H3x+u44TyojV/YO4SVQ75ZL4tx7p4zq
ytSeUeRA0N8QhS3+9YOxTpJpV5fHP9A+fHbsNPDR0lYvmNCpCILKzL7p2kMJfYiM
4hx/qWOZ1T8rk1TZWOao25g4A3DvlJkZH//JerVAhWpqRcQqeBa6/D4+MBxfKFUW
KeUrfGxjm+1EPPKOGg+PcQn2ZQ5J4DJcR8oSDwgnZIAwBFTRvdcXvKXRYvFYZZid
n5TPtRwNgK8VvMOCZqm3eCmM1vijInJmzcFMIv9IhZL7Xj7jlmAspP8YZwV6un1r
ck1sxmvUdmBj3lIwG8BN/YNZbY2wGJkAxXOp98c1Md55GuJv8AHS+6CBSbLhvnhd
uHbDXfWnoRHoUgRAaXNNHH/3XD8akrTPF6qaeCWZCed1qXPQM2nmmWcI4wZdTMXB
CFyZEKCfC5NYxmge9KpD171kfYjuoul1tAt+oXzCXVqWFxukitbq2BaGScv6nTIX
fRiNxx9l8uauqYHGqJ4SDLltL1jLO/OwgM70x8K1pB6ATNKpETidz942wRSceWNr
gfsiWsPy+uczSQQqPwTx5wgqrte9wmjhhZjGcZEqmSfC7usbrfC0cfkvCNyGrEGz
59mYDppkj0LUFMVW1uEbtru3gqa6aJ25M9EcphHJRFyd0fYADD7vXVheA32zCbQ6
FMbKVA4Aa3iR6MiyLiH/0hgmFxA1YzsNEtIb1axVv2XibzOUR8rCMIxm11qH2kEi
v+a80xOENLhXR64BhS13wh7KNkEwvO6oZxoKoHa1xXbLx/XFYyuCIUaUAHOtBSRs
Qrg+H0QowYhM4MAMrpspyfFZMi9h+SBMnfrAH5Cgl0kvPHqDAfrvC5rMcRS4QPJU
/wty5CebohnSz3UizSQoBWjpC5fU+59NLifp324GS4vU0kB7wGAo81Bts/2Rrgta
9q1s9qRnLXUsLjpELuJ0jGIttuc+zLTHYu6YoH8hrjL8QqFg5e8yMaB99i/frTFt
q8mtsdYaYVYudBuT6DXkiM6N0MHDvaJoiEOMwGOF6YQLAvy8Dlg+gRg3rAbWWBzn
vRclq0WotalnXcz313p7UwGf3iAUdnlZN4VgSMy6dD/0cizu7i6fz11Q9UNZh3dv
ps/WNos3/0a+pkBRjZVFrPUIUhmpUj/TTzor0VsArdoxFJQm7/ICvkN9nAMvSEdx
Mu5AXmsoIB+mkegEKVvUcR/Xgr4qR7mgUiemmNhsuQI4xtb3p4hM8bgJq1azDm4V
i4g/T1B5qrihIgH5KVVJBgVuOBd4+x4jOUeI4Aa4Uyi3+XrMmZ7jpsvFyaNDEhKD
jGU22hVsodW+VE6Aqis6ihTbjsTsQKlXtA9Vq98KILUPcVJXIeNS+GlboCy4f1e+
jCBNLn2sWNX1G5GxexA74EebDDWaIwvZzRrFF+OGj7ky9Ew6uSkv9CUhhwZxwphL
6Rb4FKfjlNfnIVYMQalg34oHpwDBvrfvvF7355tse3+Sl5ZYn7Z2SRGdHLBDDmuE
blMiG5ruMkGalfmFFmiVKacFXGd9DoyqJPdooeo5saAPKQcI0CDLQeAIlQMIXTSd
MxOPWon5yYUjYPD4BxfN8TW/3Qr3OSwPXjA+epqCPrUG/1hpMxrXJNj4xonOH7WE
G/eONzdF2R4SM9EnbmwFiHhXzphR6GJuI4fIShPIeg9vMk83yiDzdRX5m1Pa0mcB
ptCupYZer/YgpG1vtvZc6mUhd69aYehD2AOBlHjMCoYL5UQm/lJ/72Jhge9msDez
Ue4HLEtxvhL0TTFAY4PyZOvEuPpu/AVaG1HpiV80o+Rgl6awtpgmYhrXoK1qCjY0
USpvdAmc9t6DXI+FDEv+SpkuGVNJPEVU/Zqr6F6Sl6i6Cccxcef3r3RKx4Xeawwq
axno/bI1mIbM42rZodmlfGLi01FGplMaaRun7YPmsPbhGtuvo1gQmvPJNV6Vn09l
ZqbeIIRAfHAuFFflQf0pbZjyVsG7tihVP3CjfcwVZPFa5EsVCmHia4m6BDHG4MNE
/61vE7XxPmj0ZjA4b0CIEttY8GkjeCu3i/WplYVEWF4sqwZ/KnM1Y2OW4+UYHZBG
K/yiFOkwMJb3FeQsKFxrTIMjlJffzUgSHKCttIh9+v9BXzx/dy7F6/hJHtxa0TjQ
pOgIq+Jszen16/Jw5bDyVYOkhdSuE26jjYavK0Y7JVfQTXwKdBjVxFKBs/Udi3ea
irQBUiGzvWUzgDxSe8fqVef0W+Gcrv8BDvhOFY9mIXVBRKcSC8H657HHlHGjuhnO
dbo6VwHeb9acdetACszTlLDZIDA0Vz79Zov2IieSNOnqEOEvc7qpyCj5I7AMIA1d
/o73nZyQQH6rm/lFB84jj3qY4jQf3s+HjiF0To5KfIUa8zGzsLQGLoyD8t9EGlc8
v44SUaY0u7AfFg6QsqmlTjRhFLYhKX/6XpfTpiA1zKrpFsBuIDSDMW8JGwkk1CMi
EFx1lU7vVwkmKJceodCjZ/CiCOFIu6nfvvGoIxE54kWkwhfy/3XxeAvYCJEEtij0
KCEfSngMAE0ZalmDOv/F5nKfPd1EEtxt0gzgUb8QhVUmE719b0RzsbT+WgyqpPXq
ceshWfecRjIB/mfySfhAuZyHZBqBHKlFBDjv20z59a8bN87Admjxjg6WiDgjyJAy
RkieGrtZCq/V5rq2oYU0GDnVXDfwdB0vRoHlWJbbCVHkHVOFaji3uLT/CWjUQ7VZ
ROpT0KB0+gDFR375NMTJzQKEICPQzQvHUv6W/NnjcF5nMmMETn6jfBB8F8oRD/Ny
XMK0H5xQLNzclTS2ZkUbtTJMCACfCdpdesC8d2wtw3Hp5fHn8AznkeqGcR9wlPyi
pihWPKWxup4wZTWoEQZUzhvGby5DpC/OlMSlmOfBfPagTXg80JVRrr2WzuuiZWWE
wQSifJRJMsEIBMWGOZv8sGa2ykRoSrj/G/7Nfz70tB/TDsH9LIwzzVc2b8ZxfOs2
pUQPFE4ig/NGILVbU5wzz1vk5qE3nF2Rjpc0t1m0r0/4DmjKiSpjzYwGDgEWkD9I
VjiKDqHRPmztxnwqHOTKNcb2DJSnm70okFwT3FJRYxH9hP9RTP5JVzzJp37GKaLr
/E5y6HI4TvStB1NLPy5HeJNgGLHCDOrP+xSYZmuZYay/uF6n17uCvtO+SwrCyTeR
5zVymI1SpbEAJuLcanzYBpSWWTq4zPI0DtGBx504RNR0uPNqbtlirZV/Pqhbu7A7
HEWpem3mpqXG5q5vcDkUfaT+r6uDQV3wYv8oh5sGTUS85Y9jaoDJppA6tjf+TE/+
HJab51/j6H+7lCJjC9jrohggkJDQNXY/+sxX0tomJ9Ebj2K4Be8QVVeogpGR/J8u
h9A+v6Xc3Sqcpc2jhCkz/drtZjlIH0lmFb+fNzSc9U8eF+GlYbN/pfwAMVbaKBtY
ko9/2zaThXAln7e0yH+l0uz83feTH3CzM91w/pxix+iZy3GuDdsbhDckW23xDAdY
b83YqDcvAqNihZMbzFdJoFRx7mIVexgf2QsYryEps0T2lRM9nyK6ca+73zcrmTeX
wH6ZmA74L3VAAcHp1lym7XII2MiMp27VubQIxku1pXNf6N3M+EUGvl4NNJFjg6Nc
0jj7mZggcipZRNLo+M3shfWrrCyZE13wVZaXNi9K6OZM+Dbj4NMV/3Q/ry5cYSSl
RaXuFtfeicITH4aLp+54lkJvi+KNGBX5xnOLzCaJq0TPDzQ19oRHgQs1tbIGn1lL
+8fEKnHTwCY2BVolnEfYWVAlF6DOMEg6CMNq3UryyGt6WeryjFD+SzqyNeMdAAi/
9b0GR4pDB5cBiS0Ans0TtFts3kfN3HjEHPNEJAdbS3frq4g8nud80LiaXr/wGTSf
fbXoUqEo7ZZqfQZHD9EnLZu2wqIhCVIgxmNL9hQCimghqMCWwIo0iopbmfdGvU+l
ScYhXpdGnsHlr4el+lqGVQilBTmC9bPmnmV7svs+YRTP1KnVveFI57kLn0yh6uS3
R1g5tPhHTWrXjI8/fhanzYqr5N3S20jqUwHT0/hL3vvZJvbXwBOl2A/SErp7GKnj
7Xs1F5k8W+sNfKydEGHPOC0YsLJTgWR/fLmxkcLKr/gXYPCb/25+bTYiTb6y+VNT
HyBKUpR3IS7M33/6fnfPciymsSq+xPKzWyabbz2is9gSxm5jxneASbIEWWK4EUjb
SLhze38oRpFJ1h79qgwjEHm9e5bY1J8ctSlJdlj0ekxli3KkePThjM4dHxoJCqD6
C7c1ItduBvOgygq5C7n5KFL7YO8QqFPQEZFBWHBVsgQnnMBS2aKRYydph2QWtzeU
PQhpQ+NyQcJKKoQ6UrQhnou52j8xTGb1tEYX5uapbwC+Cc29HqZko+9WlSI1Aeli
GX+yXDkwTikV7dY4diyI4RmQvCLBvrQSO1bTRG1f7ch3h0LKkpve/hAAJJF5AgTv
DM3WbcfrRD/cvN92id+zLl/Wzpw4oT3F1TbfWRhWqvLJybih13NFOyl3ALNhnI/X
Apf4SLOXtXo2drsKQIXlQdyZJ5dYXJmNaqlcIFuD6prWBvsRwwdfSB5Pbs4qersD
mwUEUxjx3GGjuOfPtdBEXsxnRQvT6xNemkV4T6keUaTN816No4yhSO2b8uEdvYhv
8Aof/eWfmbURU0WmcEKkzvARShSBH4uvRBV1/l00I79tWodjZBbyKxvH0CaKvw+v
s5BnTG/AMJwBGaBGkUnLfPLh3/0CQd8fp0EpMe9Ne781Yh+7aEKOQnoOm6HT8ZBe
VMJcg3ZVa3wTD78AhVN7RHHyMxZFmHHIgtouEZeDp68cx7cpoMcVgaHGgD5fN5pS
wmOQ51xivrB/M5od7pCXe6knxulUtAztOqsSF4sGMnzFizDcSLljj5o/HjJROD6d
sKewcpQKfA4TmzvOqp/2flGa4/xOcRL/LEfzGPsrToMrf79DHb8CP+Wa/OHmGHhY
Uysu41fd9pFiIWBrYallI6U+nr8ejpnIobjR0/qQMXZcKSaPbZVudge7YrNDG2ri
CHqcd5dSg2j8GHI41v4xH90NXzJDb7jhC8Yob0h14pJB+mqO2zXssvte3rK6PR4z
WcAqGyz3D1sUpkfyuGZpIXicxOMkQsyolEH7Fz70FTevhAvxPuXExORoGAvTuyXU
N1P6SLGJcMtiDE4yCZ75emO3NSeYyKmEtz2SG5Gdswhp+UlkGfy5kbeJ0s9By+/P
gkoGeBgC8BH9wD4YMt8IldeAkJP+bz0kZwny9Qk5nd0IVZypkWQcFk2/Vj9ZUH4f
4l2xpdtj/jwzs2uHhbQJmpGrj+4NjONAM6Izu3cBPbcYlwCteZvHHzfATsH/r4vT
LGRpBAXxKDUS86l9/7lD9X9DIwgbtGvWCkj4w1r7+fajEf6u6WTUZO9ftQimGrWY
iR5bm46CKRc+e/DEMoN2rOgH6NFbPsq+9j9talmNfw5U2iHxe8h8RODyUsvoF4m7
xNWwGmGa/wyD7HT05Q5ErkX+bmhNaQuR5tzL83OCG90g9V4c7FQkoG95rgBMH/Tz
N90Ov5hls8gJ945si81FQC724BjM8O1dl1LxQ0VNLsNBrMS+H3zSEpVvcCT9wCEM
MC6XXatqid51yzM8TL+DVt+bfVyY4zZqa+iETZUVoa+1pSpn9mVCLhXF8DN7gTDf
A/yLWJqrqqRXX02JoM/1ZahZgriwv5o0VibHCfGJkXhlpTdBv8pHwSzykd/j0HWK
C4EWgiFohZ1nPfKrfiE+3NGUsiP1ksNVdxLrgIX94OctSyqSIsHUQ1P7g7SzB4L+
Y+wIghyinikImjRsHGtlZJ9guETTnWLxjDuPts5Wgvu8ERYBemLWR/joxmojvnJp
gbUwqXJ6qy7GbTBFrobv7Th3PpBE4iLtrCb3yERWxulrKpoFFaYUG8jGoT2/twiC
skO2NceVvFu2m/1BqMkQZNzHGYT8CPOecgznbXGZC7x4ziV1rMOGG+WMM6A1DZvP
WEOSptKgBFm6jVhK4KrI76S2LXpzsh7ofuW3+t9ETJQH6O1ZCiJeIwpGMr+TN7im
3AbM8QKwYfXT1LY9rhLwXGC6958mtpHiiSq76gTG5VlcOAIgFPtFQTbgvVVMeiCB
QxpnmudZcE5bfo+VGTTGscRCnC87OwC7nN4y+4ab8kuqPjPYjMK8YNSpLHR8bUdv
PWGJ8LTR5oobshQ+QllXzjJXNHZLoWKKG42p21GWWUA+Gco1P9TbBU9J0zkPMB9p
mAJHwnGFcl5vNQvwYApvWTUcF5FjlafAUeRkaKM2ahrYigQEC03NwGbKBBh7IZlL
w8abh3E0/1vZHpXK/YZCLevN0ITVF+CUJ7MR8Ze/kJ8gKJmeu16egyVEPkYoWh14
gPUFjREGdsylBDKspJzGSpJbLYNJ7ne3wltmFyWrbJAaKMc0bRhSF/dT6pF/YcLm
CDPb/yoj9GO/oSsXDBr8HNSd2sejNISCscia4mdFJq1EGjqz1OI9ZfXqwJSutVP1
VSmpP9g336MNs57OzOoTscocR7ohGegIkTv4iPygsuqpMqKC1KgJl/fMbd7lH4CT
McyzElCLSet7h2ln6JO6yIDBfI6eGIuKo+u5qDW3VZjn7jKXfCdNH35H5fFOC1wY
R4bwtlFZGUxUPu90dSWtYdqbDP0jRfI/mJNB71sAMk4UGR9hM6jd46jeT8863XKx
uqHnXl5W4C1efZCfx+6atrUNitAzC3gTao3AWSaPsKGGJFfDM2Vco+3LVN8+Zjw5
ArkXurWfI+V4kq6hGwtHPVY18tk7rfegTfYWwsss9zbka/cNOCScG0SAzAhJEKQ0
mXFF8A3d5gN3ydtrCqJGKgSv3PP4VT1QMNtCgEYX9Twy+kOlure2XYGimXl3APMj
zz7Dmwu5i+GqhU77pj+LR2t4ZQgTH1iPE/bCchLh+4scRyvb6q2eyw6T5fGWeofK
aIr/ilVGO9bYz3wWIqQD8kovXa2EEp9YJvm4POLseeB2SDnH9HNL9m5M1GnvlM26
R2FXruUmbU7JlSZ1Urp29hqieU9bU8spUrl5luQHSGGicVMYBHMdB8yOVQQdLNIU
K/nMt5ofpV3FYcCt+5ijwaDWk97vDuRKJXHabxtMSmuM+JLmB3z3RXcmvf+KZcJO
xvO3qH/XzBBxaT/jMhfKtPa1SC29mNJKflN7mjZquc85QW2Rdzf/klrCZK5e/BAp
o2CiqyUdpvqrXBomCi08+15f07tUxZevoAa8bXL16+04dG0wa19nfDiydVxsIMDZ
i/RnE1+bEtgEtAW+H3lH3gLJa+s8cTjFX3fKLX3YjzbCWVNSO3tx3Y0P0HQxxxCO
34ozFqSLJUfls8OJKNgM0PHojxE24OkhcuUwl20n5AK+fqpUcCsKhwM/SNtNComs
Mme/yNGwdAQkkTFnZB/kTJrmDAzUH0vJ+D9NqV0EF1vk+S2KF9cPBI8xSFNVFXP/
tMHU0g4dGgLPobsfv9RhuBv+s5A0FjSMDV2ibatOV5UiSEKhWXpfh4r7YGDEtRkI
fnGLc+uPMnGZW4Uk3MiPF9QvCuxQoHxKux1cKCT5cEzj+vKPKX4+54JscczPsqS9
F6Q2AS2s/yRZyur7p86cKDBVjOpJa2KgsWXBe8HScvbVVx2kIuUcPYAn2VJknmiO
T+howUJG3A93IE0+NI8/HCQCIuq7Q1mwxIyhHCAxztTB08lAu6iStVldcIOoLYWk
7CXuAPDIEGD/OIip6VZu/D1PUHiQaU871cUdoxYUzwEAfGpSyqpW4FmXrQT9aq46
fduh7HqZkUqmz4vmSOi/LcedOBBHJa0Mx3ZOvqrDwwyzoSOF8rpt8m1f/nalwpTH
Ip9EPoIKrr5zCqbyrmPdqE01fQZAsue46EJ1qddbhJhZ0bX3AlWzubBveQKaF/5h
Qoy7zIMUm4ktRugAVpxgro41Xj4Gt4DOqn5UAEUwtV4Fcg42vaDFaZ6Nbjodq1W6
1WG4X1toPFaOhePf47JYrpHhzogXAG51ANRpJWXYQwKdWKs6X+i6qhKJdKmNV1aZ
IY00PR2chtH7IO7T5I9LUy4fkQEPHcn5G+NKPoFv4J2ZwqVVpfP89A/0rgDNV1G8
WExrefSzGxFxNsHewIzQaUpQwt/Nub08u7fOyDa0MVx9UMlmqcV/2H1gcSbaZVJp
yrCjhUJjIFojNHObWMZIqJd3E0qzt+I9DDe0QSZtKG/7JVZ7QnGJZW3M6xLnl3n/
BAAKNFYTFo2caVSSb/MSsv1c0476dUZyFmra01BAsMQg+/2wxa5+hX7DwKmIknVD
SbuSKgT+wFyWybl6ksqntqKWGGf7AB1b+aKr93VQgV17dT8C7xXEgAp8EtAgSTQO
FSSbyN8S+d4ZcHunCgRNG+o+ypFZNxS9QaAYOlzklsCTvEVCyzNeoGoe+LxOJpJH
zC8q+FHAZyWCzy1eId0w95Iu5WjQi740reATbM7j3ytoZgF9YFo2pl0BUcVyFG8H
UsfBrGDSf0SFeQ23jM/muXqOTQ6FJ+CGNK0VugP20RGoZf8JoIHURjNEH4GEkRyj
fbEHJGOxmR4yoJL6YF8b5+8p4W2UltUa+oYfzkG3c5gK/UNxUDylqwFktacOIOgy
9e6oNOcOhnvpseB+QW7J1dD1NyUO+6Wbn/nn9yU1hgAN7gNRrrgOgAbLTcDvp658
PsBTl8rQcuWjwH9LiA/btxFHSmRPto1Dsfbn/tYi6Ss4g/15ZSs0GjxuNlx9/5CN
SDnQspquB3wCBWDVWZCLCZ1xHDtu+UKYc3V/Y2Jol7wjJ76cGk7ChAhQmqXJLsZ2
gO01Fj+KxsgN98NDtX0cwJuFn1V0Ez86TqqyzV8iHhB/bK8tFSCDkDcqSgehv9P3
BU64D6KvkcjCno9CvEZWbXTqzvhltJuGJSwLgM/JUnftYMqhsiPTtHH8czZ82Nxr
qtlQxUN6xuB/+8clew/c2p1QYv1KtS+RS2tt4rLIqJNf+y50lQYa8l6gZifEmiKx
Un8sHTycn/UqmuqmPeY3N6T+OkxVjtzyUQcHm1TYbdSouNl4jxa6PjUVsE12exsX
9lIphA12w6n1l+4F+Uf2fu4kMzeAPdtMuvEpOnK2AZHFtsHgUOAVK50GhbR3Jvd5
URm6qtF7xIc1fOWUctLnVz0b/75HswPlXxYzH4UlpDVACwlsDmZFIAXtPJkOmNYQ
vNFDnlNAgW1JAAX0YAVQyujdR8t/KNY4WL0FMopbQWQl/pnthjqpTUBt3P5hAp0U
fZVkC3SMD53edlWmnQoVv5p8YT9gp0dzWn6eCisnJTCNgInxz5RAudsg+UL5Q5ge
jiSXOAG1+KYS1S1CRnRzqmAxXFA8Sc7DSHBabXLbGQMypLQnDpBdIA6OwuXF389a
33nJ+cG0mF/qqSGPHqsIQGJsDh7lxzK5rgBNutZsx2eKfiN9RUPB6d2E0u+6U2MS
cpgVK9z6ff3aO3t3mPzCeH0N+yZl4KphLgsaprMA8Qk9pqzNLMiPaN1MZMVVJ1mj
ZndK25m93WjJt8t5gBrYH3/w2AqkKlWfr+EUE7rw3OT8C4jTJfDTSDhw2qnA3gRV
cRN471Sc8D2CL3SOk8k+V23frsltDTXiajlyys/3xMjqE9MPfScZmi8zr1F3MDo2
/nEG10kirO8RBoWRTVcyhCuc3eN7vvunDJLmBscVt72KyMcf/Kc2uk/0BU1aeo5K
kwSnitshD2Z0h+GTLZhOqJZurj8BTNBd+D67RvrQyhaas6002UN1CKrB5KAMB9Q9
M1mEYzJX8Ved2j88AqPPuQAZ6/sZa+eojgxVw6Q2xrZRpU1ABrwiXT9FCaKF1m+5
81FvVhdq2dM/sWAJepd4JOLo4EOI4KAKbXtWZCGFE34k2tOUHD0SDVhxTSq9+uak
ig8UWnV9FTG8Eys2k9lPLQj/bucQ0i+9nvzN3KzBgKuvxG3zmL1a+DvQpBfvPhHU
NrzBBUo3cHbpDlXvB9Irq431nef4ROlG0qHamAH70mhqUldacPghcGUeRQsskGv4
8W10fgFFdr3ndVI9xZKUwpCgAT5skqhJ2XbTs8DKcaPWV199N7IuTongeNe0Y+Td
TEFXiwkS4wcjSD2GMUmrTcFAtQAP0ehS649QMBV+AyCVcVuH1KAsRMkvqAAgEBHq
tUEYSyXRbvQz4CDBjrOIogB5X9eHKZGphUIJKIVv3RnPosCHtZY4Z8eCOOojKV/v
f5BAtrL+eP7WLLEWMeHpBgJJjT+3wUGv05GD4L8Lt2dwFB7B2qXJZ9hRVp46bOhf
l50hlB2QwPxQ53IpUYfDQAqbOyD9xM9RhlLCREinshnccmpodAtfSopKfx8v1kT1
+0uKXun9PeD4b+g8+tTW5Epozp/jNK93pxUBaptco6fvg9GO2m/iaVZauxg7o/fq
rtleT6wFvzARpACcU2ebGJ5BIOBiLzoF3ZID8kfPfiRsh9oHhfwQY/vmE81Ny3Ik
6C5kGFBzP7IYwi8NV04TdA2ZPWAtR9EbBeSUV7ePHaR2qvu3GoWxAhS8ZoIh1WcD
3NI/IUpe7fxux+yRbbC9/tiIkaaWrVwr/nmj6hNy0oQsXySXhKgsVCGMwCw3VaPk
6pFfWHkRkj2uJq2TVPbj5qTjB4jgM1fRAtA6hLsLYiKtoDi4ZlZNDWublHptOoT/
RwPB/gXFQIh0LXt6LIhOvMkRLFQWWIrnkZledbTS5iuev+76veAfEWInuWjB7CLd
KWTs81UTRBVVCBZMtKmmOt2eoq8D/4LXSg2wDHVQxPcb3suOZPCkbYgJT759bm18
trlMDoDdpo5EIJVDhNDtP0KdAhhsNypWMX1gqvds0m5fNY12k2Jng0uv48KJFkXd
vEJXRkUhj+ME1GkYiB7Fj4xzKNHBBN5gGNcdXQMcf2MgQogMeaYPfP0C7z7C1jB/
mYXyHO/eisQ+OMm1FF9/ti0P6CP5VegRRtr5OnqsDMIHqQA1s4w1z4nF8UhnEx6H
qEtyGRLITMRRgyp0nHPpkYNs6mTE6Le11AT4WVYQrKP0KSUOpyOjV1T3Iy37lYeP
XkMd3XewoP61Jaeo6D0aBsQtzn6kwGZqnFDg0PwUAPEYw7zki46qoTTuldp+0UI8
4b/hP1WZLyNeo/JxqHCtHx8Nst6qS03ndWlRHEEnzvQeo+mE3TASWPNe3ldQ4Imt
41k8EPt9smzC5jX+ioUw3CRXy8R/aPy7vG+Wr5l+WsloMC7Rtmtff6HVPN9MjvGC
0fz91mqvbM9Yz72bifoNyi4+2SXcLM4jS1UCe6s0PHSZuClx+bEHZMPqRSqsERJs
J165c6rWnFx0GxqVG9ekoqCvgsLW0+d71kOYsQspjRvdo2nMJFQHQYRBsrLXnL0w
gtgD3Vs4ptKzEBH5D55ozzG3eWRARgYkaYyNADq7Va3D7MPhQXEPBIzcmEmDxC+4
mCcpZGt82SrLREqpleOJxWUBcXYNpJ91GJs/MmLR2Szwnd9jVZEzSVYraSCDPBXa
8FsrY22l3vzMA6nlapSM+rZYFLNOxtc5eowu5hA1GVj9SZa3RPxTgPVRegfjSbwV
oZHSJ8e0KfsXuOkJaSkO0fxzPMT3wEOIfHnbmvozmeMvHfDwxbxZBlVSbum9dj2Q
ICKtVIBfmTKk0n2aZJTgqhDpfxustwCJACpVrj3sbuirXtElra2GY+7wglAuygdJ
F8d6INsEwLOGifosb2D3N57xDUtXOzru9thEwHJAgeUSIUUmx1IRYn+ruqSbtGDZ
bHHprGvfquLtuLWSPrF+qAO6lgfxIOx79ESx3JtCAqJi8IQkvPHJMqGNjCjyV115
xLmFNCAT6E7FHoicWyO3Ox9zQNC+168E+JcAkZoOM05crQLlb0EhKWm6cw2PR46t
a178/i+bspxp/oIZH+IzX4yMZ0+mmPg+0GcZBGqfslrrAVxALGscItE00mvHK1SI
OS9xuri33zpRAjPxXXZtfuufOQLb9IyF+3Q3bRCaWi2m8XGoTVvQKO2SpnSoiEWD
JyNX+46LFdRfv5QtBGD/igI0LeADd7mnbtBPYJ2gP0nE5TQDPjF19Q3YOt7pzt3l
ZYoYyNioFihCQjJ1y36o3jdKIO++OCdxWcQmfF2ZmH/MUC7duqJZ4Yv0cAheZvTP
kwEDWKPV+Xc6sbSTBbjalEwQ2a9qIdVAGES3cY3axwZuPftdoorSbTD/xcZ1FJ0Z
qORIzNoCI9/2/MIl4geq/eIu6+PiIkGQlOnDhReLT30sZWVMURuAWMa2AWO9kgoF
csoTNW0w5ub7KDOR1///1YRV/iZjhlO62lwqncSCftfYTc2X5JywKty4sh+n+uXO
uFJpSydt6C/yZnl9UwrfqzyVXSfKXaUuUcsPQdQLzRxJUAfWzDKmEhd9qkQh4AMN
l1Xd3CZQtNPhd1vxk07y90A54Kb8oTqtvmLtr4MQn6Ar2WBavZeqIeUh4Nr7xdJf
UNtOGqqIijWGZlgocUBTJdlW/+V4a7en4GHQM63y22eJWK+r1DuG1lfjjk6Ovx3K
s8BUcFYxNjUCLcUKtF44cFRmn60e/3vT1XF+MDoZcYxDGOv8nQM243/JM7xOqe4z
bICCgYT08QHMOfANfG4IKVJpnErclbcAcxJzjzc7oy8z0A8yPCGw0t2dvj0KXa62
xIkM+Yy9Gh/YQm/H+J3I+z3TitWDDZCa/EoGNWV64zL5ac5ranAYeBOHhCEHWxKQ
e5dXkQwMIJa8XVHc6gR0ghr20lXrGQ4W9ihb+xvBj27BKeoKEUO13S/AmTI/f/u3
uq5DaWjLPi0gezqEqQYeck79ifYbFlH8yYT2jiTl/EiotQB1BHJVcLO7jEp0OZV9
YQDH9XTGttur+p+KFXbF3yx4yC0LicQFOXgIhQCTb293NDESLAnUC8kV4FCiWlMU
rX1Gm3XOjm0qzUjMFWuFhEAOlttWkhWfbijdLadAPX1X4wo3qNtpOZNkHfogAvAr
l3C6ZoK1UH5gLo8IyZHZtGqDjewNIP0qNzam6nhQJNw3wAlc8V8r7dML073mPFgw
irTOI0BI6fe0gp8zbgRz6sEowYaY/WC/caAv/4l3QDMgZ9MfxhRM7hBLK+NfMGDY
DbKn7/6R2zxON0XcguQYFCs8OLwIp6yV+n192JlB/zQjJsx+YkRswFaHz2E5FzZJ
Eg1tpBQCFEXRu/U3GcH87MXU4CpgtRFxLYnpp54as4TTrKUAKIZ2BYwY5C7WKyAK
t8Ih0sx3HNg+rfQcRNdL9f++BT7sGkGKMPgpDfGJItCMVAKwgYf+MJMNYvg+8mKb
HghFJ74ULcIoDrvZ2ZdjShqXjA4xUzr7pvrMmW+mq2FVPOGMwOfhlxvx4DNPVd/y
nnwEkVa7lirwSx+OY9R+0HlPHK+5i2XpmfWKox/gQGp/Phf58nVSbnaAgS3CENz1
GjAJLRL5LW27xGDRbCXmfeCoILBM7SbVZVQLs+myZDihTsJyhZaWWjNqp7I+itSE
eLbx/XBakdgObki7sSi5jESLdpMcuowXrQzKVHxuW0mZDd/LJatpc1FmTuBTOlVP
797Kr7o2faS4czysTibMyB9+/vtWNHlx2c4o2jBLKhLaF5sk8Vcm9cMu/2g1ly1z
NS60jC2mnYiwhCvFVPftYwlb3SjgTQupkkNSKNBhkWRwNMRVtRJMAR0N0sbPO9Sa
ZiKV61zai/5vkYwAEx33Q+Dm4Ijz08JgmCSBElyzEb7r3UaYVLWHKRxJ4Mc/Bk9+
z0JEdPCJaJl9m6xsKxiu1YnYlFM03VslZ+9f5P6maMhajrYRgoqUYJKLlOpTWbSX
Yzj/Eqryq5R2dfdL3wPGHi4xzyIYkXfaqWJtLh3PQnrMB0FT01n/K/yHS3e0Qgi9
78P8fOrt/jgC70oMuwKPx8gURHKRaNA+6DDU11dNqHjfelYsz1Uh9Bts+ueg4Q8k
zRI4vCGDR5y+8RhgxvduB7kQ7h6GWOaSdQd2IKTW3MtNmikZyJJh+Tin3avmJqCg
/lBNfmypkCAHPqdXQqAWsSZkNEDBA3g5j/91526AWAMY2HJL2dHDaITlgcz6/6cd
IyKJK5TygI85cdmrcN0U+Om4esKnzl7NqNsge9ccIqXlm7RNkf0W55yqtSbbuDlO
ayR14thsl6vUiZMzMyfGBVDi4pXtQl4jUhWTxufRl1ytStUxHlboE1uRmeFLuni1
1NlhnckBeEhB0r22DQPh1SrQJiLtDBUeD793cxgOI2J3ArX6YWc9txgDTGv0u6wf
bnfy7YtbDuPjQ0taTk138flusdCWu5oj8JxIEBY9eKq4P0NGi7c76TxXHzUdS+H5
d9BOtHWyEQAPVAgijyPN46GiRdUu/dgO3gB7+MuRXyy3gvBXS+UJA0NAmcCfI23D
x6iFjTGphYK1a88gytq9pu6WgvCRM7eGtajSUD/6Qj8r08zSUufTb0U6sSQBRRVi
ASGfaZVijZVch3jvUsANYsekCDr+G73+IDsHbOhnAD7uJTFXGaCvzwMiutuwuDIz
yhbaLGVpao6TF5gzP/PEPaRnFGOr3fSHERl1NSO1zOCty+vYXC4187MGkT9oeh+G
6uig0pCYt6KTuPces1wAjhOeREfn7iKQLWoYgoo0Ns9eLmlYCfkmGUpZx3yStmVw
z1FKXmQN4IXie6VYhQq+qxUBnRJKdbDvzfPuMqs7CQOKsMTkqpltl1ABnuyKf3Ge
JPVdEU09zuK5num7hkCCI5BPqRYQ9rNkNUhKuoP7QlQ1IZJm6hgM5UTkIBpNHjz2
BjBY7GrMYGE731YBzENnDMw4iXFU3on/x21NRhZxLMWASAJL4zeKY2g1VdB7RvPo
thQvQjKoaXbNqtqMPMm5RadGhINdBmx1vdHmufXIYQi/KjIQMcY4X7eoucMXPjod
GdKLOy278VbhhWWdRunO4jMLaKzH+5+DyJ8+mscgtcM/iZiIuAZji1YmOjt3lD37
QYzkjxzsNtZFdQN8SVmQX1vvd+WME6q9IuwsKSBzU+2hO+J8IQUzLmeDm+Y9qpHQ
+HEDezumMSqCy/osyAfwGVSgRZsGe257316MJ8/80Ca8gxZbOLNJgKSOrfRfQ2MK
LjnLdjhXJJPs9aBfwrSxLU9ZC8jcWBHcoJ8kHBA7Oo+FaUvEJ8SuHf56b+E46WkC
Ldj4tqSdoDZh3j6heJToGEzIApuvRi0TjsR27P2+EGaDfBYEOEkSvCVaOiCaEtrE
ZZtd1gXrpxgzcdXl5Agnf/vpxzr5nsSxNf9ceIyhuxrWVX0vFLTPntHZzc4z5VYn
hhoa/CjaKr4ykKhmmRTVLGGV8FujHV/RbYeccSc/5Qj3Ebsjp/MsqmpMMXB77M3m
elAzTP1cpJshBxcNXp4jkQO1mhTZGMf+GSIFfMQp2ColL94qyoG9e4X59k81KOGP
7dB5GNjKL0KtYcEnphpCa16g5R+OI+ufcz4T2UGj8XIg+BKCOeC3cw3kJOxHi2n5
NGYOXTewcbUhoFqgQG6EYKoLg/fvNeiR2Y+XTFFiOYmvoxtbydo1huwFWiC0WmnH
uP7D79XsHeabCEpup5BVvjEzH2eMW1lciqlGZLQIc/gX3K7v/aps2dZmaI5uOCS4
kc6LTG5+op0Dt0DF8PrH01raWF63rcQCsqrgFJN11X19HM6GPXbhyEAxYGA5IRPx
wcdZML692xPLNBuc0seyzrTHV3byjnHI7c5jk82ThHquCYIu7Z7SDoMsG/0iraZx
qfBBiyjfvhNmEh4/g8mP61bedNxn6HgKTZS98MsxuRlC0Oc9dB6r7Ifm0vbaC2Pk
KDQKbwuWTw3Hu71V5bQrP43kNb7Y4RRdE/OZMgbH9Z8ReuLPhVsZXdasObMMkb5U
0AE5vtTwnrbJr9ufcjhswbAHWAKszafbFUGH3ZKKmc7oUp+INOPymy3Ewewf0KnK
vuxDQ9/33EPskcW81UKhAD52YayGwKdyxWsEFs7p/aW3rsV7lpRTUl23/XgfMQLu
al2ai7LNJfWMORjVlXYW3SvT2kwXJNnHMXpPEnL+kVH0volEVlIrUjvZbBcOO1US
q9gKyplFnBIRFbZgGr5JsJ6X5jcDdpoGQUMt/puuF22T9RmuJsgkhMD9RH1r0dO+
1wB3t6oJnxBwdnWT4pwl/KYL7UCLkbdmDPnAsmT0CoFljb248bigZSfbtTe/b0JK
8Ioa7pfA7uCK73Z//NeTN8vhJdAaFBUq7YpzLp5cEc84uaJjian/yZoAlvG70dqm
0MaXLG0R3P8kXHqsfnjZ+WDtQST/u6IqKYLS1zmOjAVQyZDwMJRtQOeCHpl3IR4T
G/YYPloEa/J6WJapLTwds8GXfrHPlyPNWXAD5jO2ZtHo5B4sqp6YbnKcU4vpmfFz
PxVKP5s0sdZIMBdTEMmVCFycBBXBxJI/Qn7YUkkFUd8cDoKpFAVHuVqIEObkNyhR
bn+VsMXjUhuY6hjw308yuNriWIE61BJr5BQj5VANMyYZYJpIXR2K8apjT/0ojP61
16etFd9qzHAM5E6ZxNXJzBgxSoaOXxjbIIG3KlFymX13qd5z/IRFRVY6uy9y456Z
51BzAIcyge8w2WNFJh4rTDG/l3kkvjnosPBQehbG/ZI7sq0MZNKw7iy0R0vr6hNJ
JUl5XZCI+ZgXi9/FQbYLEAZG2/h2RG2h8aQNvJ8Gn8MJH+PzYKW+FKCUmjKjPVbY
dvcZfpVWWBTU68/aWgnnI3EXa1M2Va7j+6l2hGgng07sndFl8fDUQV9LD+FeRGVi
5DhSrsM2liM/+8TK+GniDJfZ6Ma2eog2mBTDeJQ1LxE0+O/MRxKhC9BhR5owov2B
HajaAzZn3JVecmmKPE1SsbniSDSEPXqI67K7R9fgRdL39z4y2YMl3WaCnfP17z4N
mV3vnDas+RLo3OJWm04LWjUlbmt7uTbjRBImXXcF1XgVhDSf9IEhmU2Wsr2skqd+
IejjK+OIE0Ao6zqfg6+7qlVEXJ8hsu83t+rGfQ9wBQ+IYc65s+f4SEqRGJlzJlnc
8G9J+UgXb/icmgSm1isp/LIfYju+GSdPJ/g9HlH+V9JSKmFQZDX0lMa4X+5uCfww
gd2teyTVCOSdnLC6nTUvw/vf4o2a0VOB9hZ4FWYNXYyyiOJfeV6Lo2Lm8eWMhyMZ
/uHLRBLMn8foN2Gl1wmjY8udH/x2Eo1XKQYLxPCloZ/WGtcQHhfMOT672P+83YZB
mkGs96+NAk1xc44jVKFEitEoE9Gedt2nkV+ZMH1CQpYg2T3Mn9hqkMZtfpE8rGsQ
N/ogmMSzaqczbS5XC47FH0P12Yk7MWd1qI8nu8eH0BLLpDMT7ci2ja+xKN2gcdUX
uW9G4WQW8WocuybD++AS+OTho2sDAVm1AyYGVqcugwF/8r5vU0LesI3gzENyup+u
XYNeRZrYfRIOborxkeTDvJTTyI75aR6G6bi48CgZaDmEECn1F/RHtIpd2FjYtzjf
TvegWigC5po6dvX9c3rGjzwRDxv2jw3kdutKvrDHSLvbQM26tuebQMNJ9w0uoK7e
yr3rXajw9CLvuO+V8tLjKT0N+Lx7mxXG6Te4rrxVQ5UkbrZzOIK7C1eNOCmNeGRN
XGJCXF/1fUiuSpDSrJ6Ok4SaC35ARnm5XHJfj+Wfv7OjQUH/6g3TaRq3uY2+WYLA
SIl7Yjyy9QWz/NJhYXzZl1V0Y4PHBI47/Q8+j6J7ZTwPuuPAucuIwdeEZctXawpr
ggk7TPiyBfcEhymK7Rh7WYz3qQ4AjLOzqZG1NcN2pToxgMALklqUGhGUrJg/Kq1a
dgPG6jNrX4B8qHgxF9N+g1N1LvVDCBKWIEOYR9EQgtvY8eHzuSZxTUKGJ/zU9ZCQ
In9nvtqYjjyf18pW9EBy8svatCcaVe1rnFl5HQpOVd0mtVGcTPQQ+A5VOiyq8JoX
EoRcqLsl/t8SaHzIpmegZ0fmwOaGIg6cYhEXf4BgM91nH44NnYH5hBLGcfRaDcd/
jGUiF8w8EgPl3cDQqRCv85Gg0tEsN8W2e8JxR3VnGu7IS1QAdSdnI4+XfeCYJ6Gp
PwJsTtB0GvVpLVSNRx5svCSLO+8VqDtkxofGjmMwcw2JTUMUMuab9nBsRbfH4/HP
ClfspaR8Apq0DCVOQSYkSjAftsg1SMjtQ7l/58xmpbRtf8M/5JPKWf76H6EVOW05
qBp71gKIxtNPkiu1G8inzymjfGMwqIe39Se+io6dU3wrxwZCFzwf4hOwoc6vSwOC
juhBUApMYiOO4a7Ra8605biFoQ3rum36CV2OPwugawHhKaU++lgQrKQk+vftz/Gi
EVa49HDs/93Ur855O4lTucBiX/mHHXmkCPPybhAhk3qFB4Pzo6Zr6fDUl7JAhrPK
9hMTV1uMvCknPc85hNolUt8MWyqkLeQ0qViCeddR1dAQkGAvQRpNgNwJmpEC+qAq
mOiLAyT8jO0x8ubQCcHMBE0ZO5Oy9PbTbxckgB1viXMsGDVBPlo5dtcUdSFHpjXv
ki6/CmHgqwRG7b++wo0paCq+gteGlZfZmgVrvwvzyvAWoI2yXru/YlUFpDe3nz/v
GzBDZ4G1i1bEmZxLkJN1vGSHC/C5e+0PdXgLbgDE7+kfyloVZ8aX+9TIidsW4DfD
Mg9hURQJwlaSD+UtUbx8sbyQEHo1zsrwdW7oIxoCg4ZVJzcgZS52eITR6A7KNLXW
pcl2Efy4vWzfoMoKIHRM8QjAhrK4DVDr5BCxY2dFsDU9bGlS2obObzfD1EuZR+kA
V6rAUsqpHO/Y3Yx+0RRrpQ6aRs4YkXeUAKmJlgmVn1DAFbfEq3AB+HVmWgQbFzE2
qiRoEGMDpfNnUvp9mNOS7Q75B0SURhjcsP2xYb7Z0gbN0vj2sdmFY94BCTgxYl3H
xSI4aSth9mZlJhRUAJwySa60dwfj5A870seVaWo7Dhex4K4MF9b2o8BG5WClS39o
Z5Nk6WjI6QIAFDg+sgGqNRRqwMDw7zOTK3wmUqs4dPXIUYd+lRMS5ParcuhRzXq4
2+zCFYmqY3r+iZP0zyekjVssMSc4d1ZTNcLFiAUPdGPvKuMUr9XzeeH7XOtfcyHD
f9oi3YcWlvG1wQuXXJh67DtwDBMZktX37+leqKcdi3Fo8z2aRirz16KVckp2GCOg
JAsH44EMRrG5JyUJWIpjyMqOxY3ysm03ZWW6C8FmQ25NvnBGTIs0uUdMBornFnJW
vK9W5+X4L2HDw5vAPRjY9d6UkrMEq2fPf68K/ZxhVQktDgcplATnA3+PCSvr7x4h
8tiDXVLN6V57B54LQsy3mUoA5WZyLqRxE8bZ9TLNPXth2V6akxhkUslgx5MfrwZy
VVfbkAJTwpRhz3J892Ye0nRsHmjjrq6BTGcaFAH+tmyGV+ar0A2LXOlonOCK3CiR
z2ohzSTKTweN7pPHW5EvtM7wK9c/k2fKfCNdf/6RwA6RZpRi/nOd4BwfU+USgqxw
e75WyY9f7m+CHUW5Ues42ubLgAp4+RZe/R6sTak3lX3eOwP1vqsClCNQSU4LmHjR
q8qXHkINv878udx9gcWntuFwx8N2/B3RTySJcOSGE5NgZWbMSRmZZSOFzNCqrBBC
bqOdpOO+WmOuZ8DMYkLX0s0Emo12tq9DR4uXz3MufpAwYo7JiN2lyxyLFL3WvM4F
aHXTRl7gNyQTpERRGvMhZFR9GmUGav1NeU5oEwiUAWEpIwAnybh+vHxJ9cmhhrVZ
nRtP4M2Ut27CokUlIf/co37TN5i7Wtn6qKsMCXSvQjsxDU54wVMqJCBOpOKn+foP
TV/F6SRytMGGD6SkvF8DhW2DC0WxBsQ0ZwQBuH5PO5X61D/VtXZa8WmgfcL99HPk
7aBilkoldwGnwIyWhFElBm5YCxiffuVpfhWcjCiVTgiuCP0WuGTBKnXxAaQ3UluN
Zhq95I1/lNlz17Lc1WlV1qgELW8aDPTVp9a6Q1ExuT194R6y62hUXBMHvcW3YhDc
Qe+sgT9XbCzeJOqQzfs0ofyUPzRo5bYyNsLtlxacxm1CVhcgDMq66ZnnGGct2DON
EySZtqRg27ObGS9lRbkh97/tYNu27q04tkmWBegUHF9Z+w5fULpznYNWSxtU1km/
Kuz8JYT0pFhx2ONIn0ZkZQZo5fop0W+asnIYiwhHpLPQ1ZfkOkESLrp3oh3kjZjY
69/F+VGci47aU58YEdfMVjwXSdmdWwC34iaqij6jDMNKPFowxs87j1nkcdadZ/pI
WeWVAssWjP+UARIfwGZw3XQ/0W53tu9y5FhAW/cLlDTRXuiPN9VQxkBvLucckVcc
ZV1kWz4dr3slne0hTTaiXThsxysXSZXshtfGpFz3F8pXw8zSbhMnLfEACVSni649
hnztjKG8V/nD2uNMJ63ajCSywRqWMeh2vDTOorHY5Z6lHT8XNHO/+Tq8qUcondcJ
+9LB/+G1HcqJxcpgLpDcIXteolW1fvvSc8TAhTA5gcnnKq0IR2BuR2Aj8QBwxdzg
zq6s6lPzewoXwytFBaCGUjZ/nUlkJsbFonQcUnWOLcPW5PYUqHnhOs9SS6XORXIs
UJSIeaAWQcse2sfKMRbGa9kuwCgzclqvDNz1uLMAVd+8Zu9C1i5Z2+kypAAOtZIw
V8jf/mvT3A3B3aPEEupVoE4jM7F3dLFkgsubog3ttHlg3/qNbh28WBqiSgXwhuSe
wpWVPEs1a+QTa+pxw8FoLYMiQue6Tlv/wmmSFg0kmhU0Dn/FbxUiYjefKP3LCy2z
ZDKV0fRWupU+W74gHKsM1CJFzcB/kFnIisJY6C5KWTgykiB1Sq2y7eNyVbtUVNy+
vaQ3xCAhAhkltrjRManS87sU/eLGEiWr9+E6C9bw62bH4LMahWuHvWr11zxEx3GT
j+ePTQz0XQcP1923IwpRj93kfb1lqcsVPx7z0SjMUZf3/MN0B7CSizd80trfy7xC
rYclK09OLurkyHydHkHP0/0U0pk4P5eQ+nygBixDaKqEG0fttadU4XmtXyYQLDmW
qsi7sHUsnaXiMUnOtPRllOeAkui1c0SKRr9qcm2f+dnV5hn201cZz2+tIJ+20uED
MgR+I6P/Z0dNcpa5izd/s2UooE85QcQj/uKiUTv+ar20eKUIzZVDaZp2aYdyL2Po
jY9dodlg7GhtVxTVBOGKTfpuf8dXQXZDUMaeuHKxJFL9h4bMxRQ9Q7Sv4ACxjbkg
cQlHxKYknpMT/UMAaTARrpIIsxerV59HR7F7p8CxM/jZ3IwGEEsssO9x8LBsV6m9
BDdKeSz5moR7c67GeF6X4QDBQXBy2W/BmmkzCeH0LtDD9wuwtniKQXywLABVxwz3
SeGhY11QNphwrCU4nf4LOCvGOugc0efbk+VWjY+9zsd2qkqT2akWEKW0rxVoJZuI
XjV+FmuSQiBMUssIroiT8WdjV0MDmAocarFtf2wpCi/C+WvuV5W0dOVEhsticg+q
Aw3nvOKFAB0V0bgloi2gwaDfvdbtxJufqmPhCy+OVOUDQ71OjV+nOzNREGtI34uY
LaWeyCVIn3LdnYxCuoY3ICnA5FxHvBTPJ61Agd3bGT/3BxHAynN33oq6ZimaaiMw
yiLy+dJXewi6NIHNFlyXpctmFJtaqY62cEZJxRDrGUzkoW+3NbfV1LmrYng/6o2m
FTBpPpl3tfa7vDELgaPUoiYBhaOsOXwGeAwXs616m81kigKiqLOwj8zQZNUTbt+v
hRCFU+c99UzHgsad3JxFY+QzxpfCJTEDjatoRhEq4ms47FI88FGPbDnCEyaUSNeE
zxnqBvGIygWVFiSxcJwFBWJFjmUcRbzysNTDfEsgAgmHpVL8SVTH0Zb7U+bn3mLw
9L1bakdSlAZ5h3C30WRByyh5KOUEj+qYoLfC/w7f+VTsV1rw199Vqn9WC5Su6l+h
vDFXLJDJkY2vMK3boxwlu7CKI6PqPeKWOAqOh/GRAcHalcaoWcJg0FAY0MYlb6LU
bbgmYz5CBRLCCe+CNHsOyGLHxAPeuTi6bpQNGuUT9Cx1oZbY1o1d7zTORSLtcNSb
DvBidnd+jE0J2CJxRMcKcX6L4ykImljYh9W+yg6gQQaz0jgtC3IgpdKrz0RLOrnt
48rWFPvihOgalDU5FgeDu4vJvAlk5CVggDCEl/t3E47T3REPbJ4vguxbd53ZEImN
4AzaJkBlUlPtJonpaNhjqKIhav6aKJVRlXhgVeVfxBW9EYnlxMGXtE7qqIfNg23B
oaQD5Z25KChzwvT4z9JW08ySfvA8tVeN8PnfqhD+gKH9inGcitNgllRwbzXPyO2m
EPOd5Ro/0A7AIGnCDe1F4PRHYjUQpNe0L9Y6rACIWBX+8LWD8jQ4x+hVcSpzp3rw
+hw+6HJ4p/pRjG/t7KFarFZaqZbH0U6w2NwoMv6K5NYHx65yKQnXHAWaOL+qYI/J
6Oz6OL4fTVDyvVJ7Pf7KsivmaVvLZEW3R1LIfa0CYoa0vXLMziirxM83YLMCKJOt
7lLOhz1WM/5ildxdodreYGjkh7u4onQB6SFeAIN4j3g63ISIzTCN/d6MuZeiGaxH
E+YP5AMetyFqtAw/N6x4c0WyH8Nj1mUf2s3mpibw4J9HTUIqGrVU5mWoHWJov0OC
6bwMrlitwgWvUZUd/t38/VRW8wJ1Z+9KmmG8gaAGY2YylHefLLMGBJxJbB9Zwfi5
tEGFfc+sh46I6yzs9vre08wbyQ7IhnzDUYl00nqaufunOCxcEtI0igUXTSmW/vb8
21Opu5oy/Pt7hsCwEPY3/VTsPGCEYH1D7KXqeSUY+p721B4zs/QDCNILQXSDSCHj
+sJlcvtT1m1BEXOjnSl5tTytw/6fnAV+sq0z8wmCL5gUipFd3zUKZZConOwjGkkp
Ke5CGL4SlYeUvrV+53/ULuyqvp6llg3by33jR2Os0j6xHqWQ5ecfi9FO8ZhuNpRA
+KUTxTw+6gJzhprr2BpfD6oCnPvvnV1ACFc8+1orMkVkcGCeFq5DTtpnJGigJN0e
2SHtOLOJJt06HQ/VhSiJGmLNO7oODiDI/fl+nYRqKkO88MumVdKDTFpPn4TFPefF
uRwcJYSFIe74ULJSaDHx629q6vIgOnGD7kfjVONSz0w4T0cyU4QbGwotNrGgGfzU
2S873RfukqEbzC+rBsyk8Lx+5+1ZPtHJTyhMQerQoPkR96EaM4ymEGWsrjMHvsi0
YGmRfmR5JeMdGTWB5EIAeQhOGI4dtC/nDJQwObOSdMwITiQqe1J1amd9wv6qNtMY
qOCCT+BrWFzdWAa/kNolt0EAoH5c+125idGrVgLE5fr147D6s5fS2sY1ilYNAIWV
H7WtFyT2tvK4n48OZqany7YaVljI405NxHY57hDXEqZQ/8HeTZ1ItC8o4XSONasO
QzdaS6m7GosDFp2beAhdxIAsrn0fNmAZvWFkO7b7j3ngct8RbcMG8tGRycqqAASX
E1WcUhmr9uCOdE26zVbh+KB5j81rxbAjwE/FFkL8QRxP93M5cX+YE5H4eJ6lryv4
7IAfhyXj40TH2Uj0TbfZlUyRW9f0a7DvriDZnR+pWJFRc523s+7fOJRA1ndwDYOy
kEV+WVdxnVC+PvelVxxVGXlVH7xhx5XuVsLA5RB94H7kyOQk6JRS1Qvb8w95p21C
tdlhOD2G6dzfeD34PCazzhjzT0r3iVD5jCdgCMcRARuj6e3ei4W0LmjgYxf3rodp
E7YrmHRJBV4IvKt+RJ0az6WwqQKg7QEX7xv9O8hLscGsLr7slgj2OA2ea3dQChyK
0RIeOASAwagQvesHDh4UeH4T9z0S0BEN+Ai0Tif9vrmg5xlRLPef5mA+KP8UNZYv
NlC9pfEmLmHiEedr+AwVnHaDXaPCMJK2P/F7MhItd0Viv0PNurVBh/ILshTB8lH7
FxCv5lUFqIDHlq6xfRqa8DcvD5lqL5mYKhpcTndT1ZbzJn7id47US8FOZFseGivv
OMPu3SRIsRETyWj7a5LxDQJ+T1hktBbpl/AulEXu1OW7+tvOwNvfZavicqXPxA25
qJA0qi5lc7Li1XyWG3xNEYcirhiPq3dMFyAmIUr9i0ygJ3OGBxy+7TWkX4nogA/v
vjQ9O7pYKPrPH0v6LBi9DZAMLu436SOcllb0viIgrGjmUuqQHBkLl2JEgWZa7NzX
KHXEG2x0Wuqc7VNBB7YdBunlnG9j6OVCmkc8cD3mkX5H57B53mRSq7jfyUd9EHAv
oY0klxniJVIiJr1lbKsiX6ctSYRLxJeKmIjPiZ+OnYZSCN0U73zi8KpQPTJAtnV8
QNR2PXRimh0W6h/n+95jgU/2C4DpYXi2PH2SxEpi7d8BP2QxdiF4DECR/+eoNura
/DfGp6bm1/bC36OgyinXUvXvO8W9Od3u6lg3q6rgGxOFbv87gaAfHbPU4FQw5Tf5
PUD/Zhv9aLKtEN/W9k5+d9GSXqrsXQrravYPZynAtyyJ+HADjJqfckoWJhJvtbyK
Dj2WfAJi9TMFsvCTahJLgYe4TcSpMX3iHumFJDVju75oyR0lM5QMEInIrOwZeKrx
W5g6/hmOZvO1nQLQmFWKRMOQjyA1oQ0oc8lQCKP4pvUk+Vb6kLhX3dPAaKNFuOBr
xBgCblhv9SMLsLVhtTLH8hWNfcGXjnsmaomGNTbqJp2EACDgTvbYGYVNfKSLaT9m
8hs7L5d6NwmYHkbpEwpKfnl/G4F+Mn1m2sNhO3VJsO/lFvkoQ704e1IJw/MQ7EM9
U4zXNK0rHRUi3g1BDJURRO5KMNt0Rh0Upesgj2RfBMSyXlERA0Kr5jrVuVFlDJHs
kaSx+/LAV7inlFx+1oqdosIl9yVpjrXtQrg60dnlJY8LFJg+b4C3+gFnJ8FfQaAI
V86vtwUDMgmWq1wfijb3YP8U/JhSYDQYu3QLSbb1sTyRaUn2gRxLnFYP/PZqX/fL
ghR2rDcEHx13az425oMbIBa4ITAcmrvHSLicRJjn9oFsTsHqTN0/gKD4HA+rC075
4zXYBX+pb1TvlHSflttrqA8Z5z9x16JGtVU81PoBos5syy83uiaQdQQcRLrPF312
rXJVn/6n11IXPJkSWdCLUj2Pqks9MTaj8DgfAdiLk85Q+i8J5NlrXTYjGYPNZlP8
5cmKwLPI83DJvFAjYVmaxQIc1nx5aOyWXPlQjV9ur6ziMxaw7Ukgb4ihMpmln6Zb
UtgA1E65hSVEicoj4OkbMA4HxE/fU5xGfpfHlx9Dr9qi8rSPkp7f+13J3mPdFr9w
8X2pFO8ijHqKkKdWHOFVeXj3SJMT/7Sb5WpjmRecM3uDXzmxEZZCwbIx7dDtpHUK
HhLgn2qhtF1oC6gkMcjDSMBXkvP+PzXKCeQl6cA0CJ6kqtTH4LLcst1k4It7IFpD
f3tWKCkJSIGIr0hhyKayxtCAEH4uh3FTPm3BEW6ipOrE4IKHbZJHZ3A3CLXbtpDn
3AM0E9is+P4vI6FLnlvvHRoFTZxlAAPhLhHVEVMcQhtVQFP4Bgv6eVdWriz5q39c
ZNc7CnraZeG/BijIhzOxgQYMajOQkeN1ydyoCaVoeNi9vtBXiQZWXN0vVMMwKWx5
wA+x2foLBZ9kl3Sj3Gu2m7e2cWMFbt4aPku6FGIw/Ikj9J4XAykQ3s9QoipeFMpR
DCO/F/SoKimbhNos7/hR9dl+AlqFSDWPs65bmqQT2SnV9/Q6cG4SmFpIzVBqX8s5
ck4TIRLPTwR87zfQxeJB9igJ1x/8qd0aMkz/Ku0fmVO+ypG0DnlRIY1CPTWweJcw
Ez7H6YcmCmSQD8hrJM1ZOY7aNWn+RI7Prp/QqTLe1w0phwUvqxgPiGC09dZkxMg1
MOilmJ7sH4YnMamMmOUkdzYXozfhk+i798ie4aogyp75Pmpzr7JiL1FjEsgckSLG
ZOm1zGunyOmNhK79ronbpmqua5pMLnW7qFr9vtfDLmM7cdch90XTgAmQlbB4PlwB
v7nN9WhySxRfe0sfS5WIhue5u8Dz3efsCGNQXJbQ4G90qyTASKHbBjURrJEmJSmc
aGFfYy2YdsyohTSkp/O51Wqs7avttLLX3Utt5IADjYz8gr9qRplW9q8+RaB3J/0V
hlVmkEEyDVr7tdJzkrUbPyLya/xIM9RQz0r4xbWLLTjtGOm6jJtPOUYF5IFDGmMW
/7szvmlR9P8Ic334GBtmmAuxm/r9y0Ydbf4cvAuOvM7F92huodyIVPlM7WkyO4W3
EjGNGkLIaRl2JAOPQMwPRMF04FIUN5SLaW8QPOdKdIIltfnvDtieIZh2/NDAtoMe
+iaPK+UmR9x66h0GKsuG0vhAZPq4dK0N0H1WFUTOWjM8/pBwX36oDxUHC1mgwr0L
bEjjumfllQoejeU1ju4dZuPMoTLX8qgS8NW+IemGCJRnKbGnhjq2O9H/Wmz6Tp7Y
etdF/rz0PrW0PiK4JS/SggJXUIKacgZpIeVjGWeS5CDQ9exFE2gjZXi9K5fvZvOG
Lfsa4qrBsqJ/Be3RbYBhjHe/ZOss/pb+P1n+Pa7IyEMM+i49SAn3oRueDfO1L6Pp
tAp48wzfJ0QDDH1IIIVAp5NCXcUYyPQsWsfPmNkf77O74Z/oaFTjqXFodRrnBSQ6
Y4IKz3of9iQ6GmVWSsBuSSgwn9aPgoFcFwCZPTMqxu7gju+jPBRVlC8OdffnH7Gk
p0vzE+h2lBxzXeB7WdvyVotkC4ae4PKVlOc1yvd4dC2C2WXOb3U4xCSTTJJ/vCmk
gLiSYNolAn4Xymc7iwzCKoDG2vJdruT2T4gRbLZn4EjSze4jCtTHUhhIKJ4FJA2Q
zMhPVSe6yPna1ZyN6FdEAOSxHgqe/jRM/ffU9t3qFttELGM0x8k7vJJBs3oaEJdQ
0THvRb79PVw/5ql4g+cVQEmu/OUngAIGdSUmKlcCVxT9uTyzq0AAjWV0wkjcFwEf
2b/m3BEta9wtv8+Tme8QpqAyjdm4KVBLaBe3whPDPCEJ5DqVwAcWi+ewWZ8P36E7
IN873sqGZXvoQhPMafkB7lH2YgjSCRwefdj5w16smp5SQRcU4Y7J/dIluNMW3OLg
6iC9JwNpotrkP6lJJx04vzC7d5TxycTJiiNduFW4/b9+Lu+RoQn2170jxY578xag
7DsMbkUgbtr6Ofb24SkBvpCLKI4OSlsJaNSvIhK8ObyrdgJPuAZ1Qt4ve/5JUni+
I7Z+6E3Lq0Lr9aKOrotpQpsIXMKP3PrCK+/iZyCbcm90awgV4noUOEYwmQUZFNAA
Q57KOL5VBJaJ2x1gx6qNGiYaX7owOI3Es+xrFJ7BF1IrCf5pPlKPlYaY3ug7E0Bq
3nIagdEqUDyaN/CNK8mhB8xqnvcBtIcU8fUs0+7eJPp5KtquRI2AhIwJovRiP+uo
HwYmQvVWU5Ocpq5JHKeMGO3ZqjEqPINhg9Opkfp24Wo1xcYFlEI9qUkmWYJsDg85
c4AYr/tG0DUAYc+B+zXPEouE5ANV8IT3HNIJVTkwMQGLqVvAlWbAurzSl9/U0u4q
Pr+uidka2ZkqK3kB4gJWvZnef1qYNq68RCUM03sngd0uhnEgq/XWQjWB7xuDsql8
OVOYF37ftKA/xhyJIcy0c0tCxX+9tU/mRyIZFczPHrygi4+kuo8atR6m/aXuHeOd
iB7fHQo6erZqRAxLuTZNMYHycqC26TjKpRHqlS865S4/rZRGTz7mGWG6XkED3SDa
fsIRGP5+yCicJjSuv+McBNzxv+esMxkJwD6tWTlyEjyfd8YfCnbZoB3LMOij1IfT
Ia26qzW565iDhPMQvfIzasH4ucSyJGhzC0YK2N3p/C+e/i/eEVaxGTbb3XCboauS
qILwUp6cBj5LzfbTYPaUxVDHTmbjvkobLxJwICa3ROmiSjuAUTurALgl2Pzarl0o
1Wc2CQR6Gnl+x/yMrXkHEKjaxU90kA+ECvgKkKSfIJOGLefbYPKYkBDxk/ycWgK5
3bETOo919uGe3WAJcNFtzxhBYEK3WDAME+OpMDKEhUoZFIU70Y3IY7z2Fx8rAmgR
ZrgFVon4GQRRlHTrYe6sTfjLjnS7ryM+9rT4n/pRmRk2lSg/HhzKid9Kd6pROYyO
6DR2h4RlDpp44/x4BEZAtAJPuTfNEYeEZsrzUG/i2L87ZVD/q5Bq8+ObMX63bLYX
Cv5rGX9xIbGEUYhp5XNl7XySoCWS0ktkIwhddccf8NnZdvkF9z6wGQPGfYJ+JDDT
DltlX4CTFa4iqXhJdBRU2OYkx+IoCUyvFRBwe41qtF/JZfe8Upt55zdHEq88vDhs
mgvWu7gjv0nIWsqT9kKAeyDPFL7amIEeSeOD6Okdhm5oI9nLh1M05tCYeQgnQlza
gk4V110M01TeGTT6Vn4/QTyUhhZPL/gDi95HCIau2vQSV1cg8KGfgH+uquVl7y/c
IeAc4UojOacHSRF/VJDBE7cSXAC2KHxsVujfPkh3O13FL2LSzIqYgcqawWl9Xqm8
1o1x0BL6gH0xcUWfIKkvUO/8m8znkNpf2sZabKjYj19x9df1pG+TTj1BKpQEti05
XFqWMoeHJI8Hyj98J9feogpbEvy3IBHoHMEdl2wznJJJFjuvLQus3fx/YcC7Fn8V
rrxrixySndVKWk1Kv11htECY3GGHJyoW+dKXzHKTqtvTZ4U5wAyxejcitBKIG5dG
51nJM3weQU9DTUnKaoxHxeqZOU8WPttqNNERatvgMN6IquWwoGN8ohPiDmCU0tdY
WKZGW8B2EJPBm6l5oJga2gPca+CkPSrVolGAQlmf3Juxz077YEhqjXpwcmMDIXrf
EqTI9r+wLIfIwVXkdOGxx3/SdT3GkfqGXHTUjG1ij39GASR8jGf1g3z4zh93TeHT
YS9wBqK1mnAf4Y4teAru4k0usbx0d6Eo4P1LxB/uzNfpou+nCxtUiJrCB50mt6Er
5lNFykQVsh0tU9NEV2CY4Z9PXbw8SM0U2f37aU6F2jz7/Bt8xtixQNkPz3HkqzU7
vduZS4xKFByrXgoS2TL9X8mC2mQcDXNjs2UJZA2JsJNen5fJwnydxTcdjOwZNesd
5Qjr93nwhWVssOZd8Ri1dFLyzViPWEzeV2D0HjP/wXwoEan2qfi5ncgrzcfgHjRl
/YSupUlgmFG1Yw4vzseX9jIzPROqE3p9xsxq5G7IrUQbRdDKq+gdWZCY+LBZW2MF
T9S+MZrtMROXhrWdgkvwh9JhIlYLiMVpnpgceoFGfATnviR5sjWTvjkpkvctCaNE
1WwHnmjwfWp9YrhfiVngDjHgUF+b0AHS901bTFLZm+kX23EbKkfNCn7c4TxkDZl5
qfQP+4/QtzXPAQyT6/ZDp+jou7Yl7OOxDJDi5aalx3/iCJ+/HpPk8DGgICXaZOAe
ZHkvObtX+jfXAVrukHJ0rHRr9p9F2Ej9wOhvTQ8xbXLKjrvX9TF+6W44qsxU2a7H
O3UFihIUMZZRYN3MUCHfFpxNkgGFP/9dN8rR9kUzZvmahrh+5VVJ5vuQoOS1RweA
zmv/L96CRxfYmER4atjLIM/sR2547YlvjvHov7mnQqcqijGvxhsjTnDwcqinpoev
IGXj1PLCBJEHUSAGJ3hHGJn1Fbv/ngPukPMvHP4xUvHPLIMt9ZV2D7L6OoVvy5Nq
pPDAEibi368SnTzxS3WsjYV3MpAMkVgsoyGNdhLbhTA0bChsGXdjc8GyzTjAVXgJ
1aDdEpQbnPGgOjeKgkaXjszyXLId5r04HE2XNnEMUgv+4pacNVeRFg9Spe6KrJcZ
e/Um6zOpAEtK5yDexGyeQmbCFoMCgXWFJJBJJXiOmlWVY+1qe7+v0otdSM3h7Y0T
zZdTr/sPj82ZYOh+mckN2YhUnUbj2/kgqLUeQrp/vMc3dcc3RNpBV7Rkwrw1/y+7
Bd+kQtNY8U+pgrfDQ/qD/0ioXqNdFKS9hXGJ4AcPwyBel8a8HMp5B4jrWd3hXDFd
FpRxdAkTL1F/2QWlP9/sqvZeMIMHUrYXQwgrpFkGd8p/74oYTe/rdRKbP5qMSwrq
ys1KUJSkhKF1jNqQNMOHLOaMM04WV6MxBdeqO1CKUGrTREbgEds+xZaX6GAqlhyB
I2YpFkyBocZhdLZ20ZrjzQRY6FUN+GSxGLuL90SAnYMZvOk18fen6idwhhUKMnV8
WgzxmWamRXs9K1oPGwYCJ5oYx6nqHnI6UgQ/8J1aayf5CvM7FzRXTkBV/+qbTYC6
A0qrv+uOZY/OyDQQS5UkRZziXn0psdrUhp8cwyYLK+kVaC8icmhhRSQkMOjPEqBq
3w26HSolzLckmxGydZDNLs6AsYLv5ozaMfqEbksuHThVgG8IreP/G7jItqSHfUhq
c0AVw5eUcgdxiPyzV05BQTMtP/zSdgQi1mND8klDum8Zv76JSo7NNfLF3eiAZMLv
X7B/aC7fk3p2hLpDE9WU5cGpk873ZyayNYX956ioWLzly7XUeEaoBhyYdMWPJg78
iEW0BgRpUm+k0/0H2YXPei6716jsey3wsaLVvC9r2ZznB8ODUBC/Cs2R77WL+ZIv
XZpZQ8Y0+B4PmXy93q/EOEISma8YcaG2mqt92Msw1rbPlP6+Dep4QklIHgJGT1yl
Vr+sr+CMlnC0naO3OZyEpppe/m1kHrTG5ZsT+e3CMBIsNTT03H13dvUQj3tU1/cI
907v6b2tA5eyKYxfP+f9BPT7USHmFBps6gDFjsgIh03XxiqZ7KMI820CcF0HzS65
44a7xbi0T6QTFxutvuIp7dQq41DFnslQ9ULaRuo3auEnqbecc70KAM6zcFqq3upW
n0Ud/mHW6Hk1cKfDtj5sk3Tb9UTuYGzqXmP3O0upxcXEwviJ9ak3c4rK/AkpwG41
YHAXKbx+cKI0e/p+M2h5Go1a6onibUqK205nVYEFgd7DAfnu2XG9CFXEZgFUocXt
SwVHE+jn3MOpiYGDmaintA2QkyBaorlFcABFmwmX4J6ZrYCBehX0jDIzVvFeOZbo
2OJTmeguHlrCnTbGOhMyGd1M/W5jw13jHOhWR/upafXzcagaM/kKW1/Exu1G7HVD
CyqTeCX/jLIA1kDUJ+hsNFe2YrZD5PGW4EbkwpgXct8ezIGuYBEDskrLkrUsnkXx
r41NDrP8C64IOKB57xRPCBQAv8uSJyVm7mn52EweeDNBJya7H3aWEssqc3XKlhjL
Pxhy1twZzFDjAexuzZafnHEFItNC3/ZvVPWPauHhTJ5HbUJ/imRCIpm3XUvOXXaY
70cbvPAEQv1MB6Uqz8Jwb8Oenhj+Nsza7LO334oFyiA2ForSbfo7LbGW8NrVRQaJ
4S4SdkAdw/7Fxs9yRC1q6PiLa8vNtb6Pp28D8wKYuyf3yITPil4WDoLKmPuPRLY+
i2vmD5RtTCj8Nn2Ztg76Wwwwzsfzv2kO6xuGtyC9G9FcY7yfhxUPokv7ljXkuNjR
AazB525ke9hW5ohWoR7WGdIzA8ZP7KDG48vKCKODVi7Qidmwbzn6JPDyjQMNB+RN
RuPtfzGXobGKcMzTNmKHKBgKifWxD+2brUOkseUFDJcTX4gLqGD4A5d7//KP5cAq
dv7uaRwhCa7IlB6LHKijFlSAFi9tCJkDaXvPXvXjjVF2ZL0h2OKBWNfdyzCOOP1G
uYTA7zZO4PRjvcBfqZv4akESAuzn9VuFDJWWxBW5bs3OK8leydYA3XVoAD9j+zYE
wXiBBRhi4ENi1KUmi78Q/+Q4Xj8AZulcXYYCr897jAsfLNo4CPhm76WLSd/YZ5Du
v64einBrSBX/Mga9CS3lI8ROd5aoSepJ3mMEe2zV75F19Np+Zy3+OXKrFtmSkUyD
0BgYPy/VbGW6usp7dRhEdYEMUk8gUyczRwNLcr+lyp23jvYTJpX+npE4O88t/pK2
h8j6pVMM64Ksj/yC1hNCOHNER1Yg8tP60H47vluIYK4fZJ+7ILUjtc/yFb72IXI7
2CiIRO5AyUtokNSF5wfc8OIGYJcYKQ3ne+QiLxWmGfc7vc5YC7mJZLpOuTe9SlPx
ggEW5NaQYVSf0CY6329uuWP4hKAal+wWrma+P7b5Qu0cYFeGFZZo6GSu8sJ/gvC3
0tQWuQaIJ7IBwjaCnAMM5DTqLOZfzrxOg0YtT8A9gVJEjRUAYLhy3ccjNJvGadZz
+DBzPizgc2HXpEw4Z9kJcUdAwxbFoxLskF/unGiGlAMddoEYgP9eaxHVuGpi7ESN
97sehsg1lDE803pIwExoe5vrzLqcccHbHdrIVBA+1eEyk+Cn2lQdG0PJwPcJPsc/
CcELUGMVn5YDM76kBVa0XWHP+F7hw8D4tJBC0TPmYdGa/fdU+0qM59hormPSAsjo
lsjG5yspRVGR5T4PRxxSB1ei6K7rKjOwd7hcifWGKSmIgXSgdC3cRjnl10vtFmrG
6Ekv7FVVQt7Elp9lB/6CmirBXQK3oPNjiN5O4Zw2zPdQrsetKo72N/qa9Png2/BT
QpTswLMEgoFPWAhotrNmA6qTNtQhEmokr5WhNrGexIdlrRmQg9L9f4jOV3KM/Yuz
U3ie42aByB22R81WV4n+46IMdIDXSg7FOubIE0WYvWJMUOYjS9wdRrlUlsq1iQZd
8qHIl5bP5cR1xcAwqt/AQfQ2QYQ13l2UU/pSfQxw2SURUO/OzEUy9xl9sPlFAw/U
M6jaq98BBBsF+yrzOcod08kg09aeDjaCAryd342d3z1FfAkVJam7XunD1wZTlLNP
ahq0SzhwLijCtvy4XShYPLbP8T0omHNR5E65FloaivQRfcXIdIpvV1j6wzTR/P1M
UdhMlFQqs8tvQedKPeKK3gWYKQ5I3LGwuctcFgWnq+PaFBe/9xXPtPyDYcoXrn9/
pPv2xOsGqJiApKomtlpJMuo+WSSO/4Cg/HL5oLwulpK7c5D28gLy3YizRZDApuTM
sLwzaO93hukYE/8I8cpplyHCb2wQzb2ka3fNkRIq18sNmDuMB8wom94QNyayKvR8
6pTNahs2+v40GElp7QMm6PgybeUc/9QrJ9evjWkDrXLbcBVWkCIdAvsxjY7gHPh5
M8PVfXdG6wdPAAsUnR0XGteCTMDwp4dVn6ktPJCcAeeXsmTZOfTW+sEDJRS7yCFh
PSFOKDqSvx/tFY33sY3x/IJNQCdEaIaOnWRhiQLBoqaQ/2FY234iL5UzYOXh/4gi
gkmCxYPtKncOuMQV4hq+uKn8Z2wPDTk/QnI6wPo8ALlyZ+ZiLXKM6ms/2QUZZnUr
dubWI2bwqMRYTuwRuomj+XczERw4H8eSIR1T+knKpSFx3EJ5IfhtbjDI1pgTPHM8
4Ox24HB3McG8n/Qk/huMFPuMdFkr+fjRbBVH3/BNyBcERYRFdwwfM844vlwNd9a+
xvnzjt+y0pRdd/S/QbaQxqN56UK6hrSr4C002pRZ+PtmnNHQSC9qKuJJyq+4rlla
M39V4UVyiLk+wtEb3GAFIhs1nEoXsp4c5NoijAhJ7tcJZtCbPzQ178f7ikVAIR37
dXbrVQQdIhVD/g/yvJs1bSwvEk3fkjRtOtIzDrvb20opwaNpkI6XxBaf6YFSzWNg
6uM/+ZsL7QaMfcct1OcgdoANazKYkxYkCYCEeEypPzsQaeOu9yeh+IB8K1xQXg62
xiNN+2CXatZSSfw+tmb6+W1rqRPcFwBGWqLNZmMXdO+akW8JHeff56K/hm5LgtD1
vnJCpjX2/kCmf2t7BJxItRoItBKamlWUN7xka+73UuMNDnD57NTql8pzzNxQxBZ4
1vUTznjBDoZaHHWNCR3TtKmGj9XO0dAXYN8YpcPMq4Tap7TcmZt/i0ODWPrSpdjR
V3JCFEPmqNRbEKagmw3YHbe60qqy+GH5jON/FLw9gk0njGllQyvV4XWNU+fxm/CI
EwNj0p91o01cO9UJE8jVT7ya2fEco6FGQRBygIZxwCf6DHW2t5JU5Je7GVLv5GrJ
03dmI+gxXnYas7UCIVneauv2KD3WiUJ9LN1tCLIi0DCVFZZ0j0U08LEYkMcci4ul
yfd71dedVnpZ9KrFZ/FN7oXjvh52J5q3HgRUZMB7hx2SMavZETLqNCe/fBQY9oR4
/NTiUztj9lzxRn4Y1fWU7zZ5/x8cE1HeUDtZc++dm3UNsJGIwZrH5bWGkSq1dnoz
l8wIhGvrsjJdMJXRTp7dtAcCErCVstNU+vGibLwatdDNUNKi628fz8oH+hAXQf8W
/rpeaI7R7HH2+o6Oa0bhdTquQNlCSJ4UBU9iB0aQJld/CiaMEmvXIPeC0xgZclWW
1E5D3cATIMzQ/4LKQtbUMFb0Hfs7TRKsSWanAG6JuTRqfhTVe3tPypGzU3TTtikB
5Mo6nJQZlxYRYKeWFSdCsn0n+o1N1/XoMl7r7MwJnEZQ3e9Lhs6OGtRtReygAw74
ZRiQ8PEYrkSW2wJkRpq19EPG+rtklkWvcWOejHHcvNGUryLAZ3FAE/iGA8bQysOX
GrEsyHQhiycL5pnLzyZPp5N+l05J8bGuK/CpdC7wm/PnyTXmYudaO3KDur70vo9e
Fz9wd+52furLB0D2peNGvv4jkS3mYxZJcSbxOxToAnVSwp2sWSQpfk0YfJWDDyZX
c3fVNr/coTg6rLCElKpoBI4V5zeUuxfBevpjezm1dU7lEXzvmJPhghA6qR2D8met
0bohOcdn/UIN4LBbp3Y/+NI3tHM9CldmXjjB4+NE5BhgjRQtItw597IcNTcxXCcd
XElyaEHWMoO48TCkxxIMjdnquzBw/VNz4Jljb9Alq8s6E2QLHhEXDtRc8vLPWHWN
8PGANNsDO7Lr3O7TB9I6/iIGhhj7tIjAEIZgNKOAJave0xlSMRibv7rMmpViH/AW
7BnwpawXnwK5RLsjELdlj61OolVG1eMJDjFwB0oK7MDyz/gHLv0L6GQyQBY6cOSK
NAKRyiZlVdWqc3ulgjtlSJQPN7EY2f3l3TTNWO7+BEPDOwkQpkRR973PZ5AZkJXc
ZRnuytuSuavU6L6hduaFCG3wpLZWNytxXp0YIm2Pikp5HGcik9jnBjAr3crptN/s
bjnP1iN8eL6PXdZ2iOzlyA0auFgA2qHn80adISwW5IfO250g9L6eFW3NusIb9uom
YU55K5wSNYbr0tMw1jw3KMrFzBa/yPG8HnOt1iSKGerznZ7ykrHV6hbdO3nevxkC
0lqJAxiXSm0gOQE2zMguRsKh2TbQtENSCCmN6s9s4NX7ID/S0EkZXe49GWfSPxkF
tedsuRd92Z+WSclcICZ/Mi9YWnnd9cqu9KxKoGLBeDi3kwJKN5DdpALkK6BpXbjb
t9mT6lzZJEZoDLeEB3973Uo8oiiY9IfVtPHaWzxhbhkmo5Z3ACwq+eZojBDf2Vb/
OyTxHSyNZeVkfbboHd7zPsZqY4WHfCloLnXWNjT3q8OYV8JcN+yuqN0prIhFboYc
uIC8UICwqDkjTcVvD2tScF4OSxtwyZ6A36lDIVHw/ab7X4DEYviG9TMVHdvp5+Bl
IE17gPqA3huJdSDA1+Ul/cCt0S0EAfrS7N/hCFrJUL/CF40pi62Powxw+FdrUFtV
xeKjelTO3Z6pZkPfl2oY2yuVvqrZpEsKK9JIn9d6+FKfj0Vnov3gyQ5CH+Ocbb68
egWN6uchheK3sF6Rgfb+7D8JDRO31P3UqCIxxobqsGs0SJtnbabHlmT1LNStS6Oo
PxYd/NgcggFcVkg2p91R6JkTsdqhlqlDw2aJzMiVoCRd3Tpdg8lzO59nenwLs8Ps
ouy/Q6p2O/LDxkbnmuMEwJfvMYZDEWoLW+aZhLboZ3OLJYVyak09slN+wWGKxVSb
IL8q4MC+tTt+eWoztiZ55sOGJsQ3YB8x8z9npyjYucK3rIybORX+l6Kukmojta4H
lSKTljEVZP8dP94qMQTyhcpgvBJ0bPHFsbxgOUabG3WRFtBQ9sVA1dF225nlwCgo
9Q2OBr/ovFaR09ZYwAmcTMZmBcaD3DhA0N0lf+y+Tm/xY0S6ewe6V8o/y0gjg3n9
IhlQgnhPeTo8vqojk7v/V2BvNRNBpkercmOUkwmvxKoUT/mvvqaM+bPgCgdAdF6n
mF7JGJKdTwpUMM03ZZwLtMOnpXoZjOuxsAzWCdTBevOvvzq3m/AJYhMvx3bFUTZ6
eH5hUE+wVJnyT8LGLGNQXPB20o137JAkBzBywlw8ebYBBbmZyozyVGHFqOErGmTk
EYidZwmy6o1nPg/do9k3cFkY3yS1ExTLaCa2aD8V8q/4amHk7iKHsnH2F1QZajza
NrGBvIcvt/xvkhy51sbX6WUa+Yu3m5XPViv3kdjs69qd6Pt0vF3u1oc02ES7wLjw
4bZKLX1XNvrLvNHJ6iZa1MkqhEsENji2dBujf1kr+6ilTHMXBi1KS2rlXUW/E2Um
PZofEFyW/sNZVFVLpBiHX5wT6JJd8g07S9iswhqOF399xIVw+O/adXjBOSwv4XvU
0xeyRSqFfXrRUHJJ22kyh98j+2twJPjAKln82s5/zCs/SoG2Hn80vm/gWs0fkLe/
xMctLOUCz3EMZ8OkuQuY4wJ7Am7MqrkRlPftnwOnqYkpmt5RZAJdsECHRCCoZ5Qt
/zdULThfwvCuZakaZcbjqLVHb7jGh7WYPRioOBeZt/Qusl0kVu0tP45u7Kjv6cJT
guMCFLU00s+AvZ2iO5YO9EH8X6I5J2kHP3X4B8tZnUbRIuU7x5asnYtAEJtmBudx
ZcIA/OYKYlqxPID4PDUFI4Ci1oA1BqaYd5g5LdNfaNxpOEItYAQF2GSYlDG9urKi
HtvBBBZr3NtTQTk1/iPfDu7ISzrGs8DggRSrLRtNV7RN5N7Z/9lZ3QDPoGd0xgbZ
W/QWPgKbMvaz31mLv9EPHRsTiAKTrYDghubjRbUF3mrwJm3cxszvKpJrOABqHxoD
znpiimq7oIR5Ubvv8uymet+7CdUZZIbtiZfAFIcUjtb39uv08HkLdpLsyg31bXyp
S+taraKCMQkNWsvq+tGx+QE3qCy62TFq/K7tbpvBuClZaDhP3OuCMGRefu1Px/3P
Npw8bT8RmDBymo6TUEvBQXHSdenh/RV9hr8aNsTlAOTZoaEHeQO4vvQ9q3p84M0h
9wwBV/BvmC3v70Ko4bEbyHdllaT/TnA5jQyEf7D3VGf4vFTSRFVFQo0c+m2W+X2s
uW3u7AX9tj/No1mnP0Zvd8MuHaad2O2PikZz1uMtBywSdV01iFgvfMSUiPDIGiBg
eXXg+H12M+RUCe7I+4Y26BuzwIE6Sm/OgC0ZSSaKHOrYaoYjyn7WKv2T4ohCYJmL
ao6nrRJB52vYojPes+tRlgYuNDIpI8MjUgPw8pB6vWJ6GsS2m9a9N8TpVrUaYQd6
hrUVr5Me2Zs31ElO2Oewa+5L6GxEdeULSIG5Y3QyNjlbm+UOcv+ECED1xp2ZWbE3
yazYGkKtSPhRnurEepiHTJ0II4WRg+itaU2r2Dxh6qxW4BpzxL0nbujdfsES86t0
kbOcPUfv3SK2Dr8VlkiVU2L/QQdrRQVRn1+TLOQyUm3nfcru9NwT+FZcS13aUfTS
brg7aChmsdr67idGzIytOst0WUJbm7eAqt2O9/XOsB5VIFKSaDn3Hp4bt5znsNl1
tzrvezwX5YS2LMIb6KUizBbjVjiGlTXHMP6dP56FEzhENB2PwFdBoO1c+6wpIG8+
FjMqx2IBOBVPISvq2swaXC6fZEDK3Waoo9TO+vIsjbsFC3Et44eD4RIDB06x5T2r
PvZrebjvPGE1NcI0vQ4I8303TXdXdJmNa0gP2qRrq148Tgjb9TdAWi7UIeITee75
S587fUrJW4K9PHAza7mMgL5RaRnzfxAjJDYBwgOnC67kCqiWjIzNzrHEoG1Gyvlq
dDmCehL1PKMwER+LPRVodpQOntl24crmY3cT0C1w67ZJ+8U/y0mT1QUDewp+oNOw
uH6eTx262NUYRGgmq92PFqJd9hXv3YmhUwdd+8COJqy4JuDcWFpwOSpLAkxazN+G
XlUxmpSeetVXhJpB7Mj8oZf89t7gcjOE+QoVUqCpchPW5gB7McOOGOHGHIk4ZWbL
EIw10aXUAlUuZZgaiC7J3OVQw7DdqBUPjF69vlC7p4vdcTf2AXHLqYKUZfFuTpSD
c75GWexQOh6M78z4vgynWjaEDDCzpBjNibd9iSpbWMdPcL/QZ2bJiEvuiExMd1+o
Qd+Q65F0iG7iRahICMGAa1Xbha+mQzRBGheVk9u/WlPJtEOF5U40J2LYavR5RDTA
RuVBSuMGLAsyosaRN6bG5oIGts16sPowwfIzNeXaY7f8MaP6oxAR4GCbLwIW2/zf
fA3NbN3kMLzHIyInwWzLVsupvAIOKRjy1xeCtnOY0HfGi62KbFufMxvFkj4IWprP
9+ki4gu6EHVVf+k2WKCxUgGXm2j6KAZB4K9I8B6KQ9hgNfE9mqUn8UNT3LaGaRVs
wl5vgEoJhcZFCwZe3XpuNQVkMnYT05OJxSOLE1sUxSYeZwafssy73rqaN1h0tGys
5OT6qoQWk9uW1VY39tlQrXs90HSdgVFODtyFoJM/awaSKclt5PdRkQEUbH9FEKn/
ZNWtNPhinq3uecNeG+j31jEtwINLlt6z6+qEZJVqofNt7Al54jTh8PwVtDiv6z34
Xf/cGKbmLIcRNZ+ZHBAIUWujrnht0WKxpK0YTIvqEDJP8V21V9SbsFTFaVt7SKd0
ACdRQjeclMO5Mr/OtEQIojzYZp35z+TRB42XxkSfC7eh2sPaKYvdUYXGkIRYITya
AzP+fkn/nM67qEtj8RpdwDxsPkliVaxB1PJ3TPVMqWVnav0xBwc3V55k07Poa3Jg
G9bek0R/RsROgYjaCx/ZcR6CZCG+emhoSmg2qGSTyC4TTEl7q+s7sjscBy6Kzba9
PdKTA1oYH8wOF18dHhS5hoQ0QadTJxQ6NXGQE5PvWvoEh2ovMMbOYmaMPAE8qdNM
W203oCAvHFv2YYkau/w6R1i0pMKh2qIOgioyZuMVQQB5ZyAVFV/elDEGPlFiUvnq
1jFjbmJPe/NQZptg+DISCNDZzbqdiGEhdE2jT6trjHVW0ROYsAX4R1FjpJUguOgM
3HLoes5BF+rW0YfvqoLAqHS4brmdSehcOiMgAY3DEnHDEab5iwG3TcWc6GeA6LQ0
imH8hFgrMYxM2PBHi86657vHjcVoY4OF8JkLa0ed8phJ2moWrCW6gUkQZka8eMVp
R382cI2hS+dCeXAeq/nqBHW8aCpUEJHpU+TxfoVj37vd+4elT0poGxgD9BYG5Cbr
Pnfn3YBjeU9iW51uoVailzcOvtGLNELxC1kbkBheCwskNO7qTaVAqgp4J9J4xien
2nRKeDujh0HzGeUmC08szTMOOVy2TMj3YUDCXv7eBwVRgRNv0yJVpE7FN3WIsgIz
zOLK16soncJI7QWb4MIQyKQ776Ab4EnlNwmnVUa7C5OFWYZDYJiZr65tegURDz1x
qJ9fe3++XmZTaLq+25Qasjut40AH58aeiwPypHw7Oqaf0g8NwVMon994B5dhOYyK
7OQEa1twSEe9ATfCgqUFPFDvgTWpYiz1u6zryZZJARL+05laCAJppUK2mJMZ6o14
D1/ugMpRnPURoMF3HqS1G/Kr2Dogjx/1OxcTIdUE2bhmbtrwwa47phtSTZiMlSu3
lmgaQe4DGPtgEuCfXduBH0s93NU2Fd8tV3jKpA5SBlaF02z501sOlVrDwRcBFjiw
JMELLjWz+HFn70MGICnXdG7iAaWk+NiWYgqYImC44siiJdkPMkclDPDLmH1cP8DN
LYWBGJbOkQMUHGekV34XeRAhQBO3pRGbVb+7K63NCJtGSNTeuDtq2ytfGNbXauZX
UENKmHYOSEnFKuEW/7XkjHLg2L560omqav//P1XOQ4vNuXj713m6HWKxHH/rIS+M
hwFBt36DrYQK/nuNErFDpOcwxalaFXHxjeG0GE2k/+5jwkHiwcQgx87J6DDRPH3/
JiCW042Tb7X+VjDYDnTio9Kk+pb39+mlUMKU9m0UPnhKFy6sUtAfhwqbct4g36lP
jlRBlM/1qbfIPOqRYAq+dY86UXxagA0tqhvlZLDZSuBKyei7XQXOszu/veouN7yC
tFBRaxkcJmt7OD3OeRvGEWWNBnUv4fwu2ukxzGjiF+jnF8hdazRNC3VaKn8pnKVL
DBqDFZLMoC6gyBsVPoAhXp+NjCTauVrHNyd6tJPHStDNwjr6gv32Lbeg27nCsfIV
vA4IOugsSjaF6shgIfoPPju7zWPMj7KDDqQyz0yFfUMx5UE6ZrX5PrKX87AIpRFF
ANeJDPiQNE/Mn9EDYoF7ZSxI88/FwcC+DppvE4WCE+TDrLdcE1wC4FyGgyBh73+5
5LzYMiK2Serwz+V+UKm2l8ZnNSInALh+KTihzFEmfI/O/eGpU0HKUQlr0r3MXFTE
Br7ch8pYvNurhz6LKrA1o3YEc4P9SIL1+gcOiWEi6XLoWInwiZscNN78oji31VMW
IRs65InvsocOD8lRill8jSSEno6skesOKtCYTSyebZRIe2spygGyV34vWqsaiTZx
QupDVPhpwIORQ878ClTjkoyMgkKsiXuS0u1WiTspuwgaszpwievCB2Wfly2Q1VIB
WuKO5HY+TZk2GqKJPkxzne9DmGMJZ2/mpuWJrCAl0PyTOdQu0b1/ch/NybNAyPXc
IX4YLVtrZtgaFQru1jVisEocuP54rLFKwzZezZst/Uytm7nRN57+ocBW17lCxnXA
99bCzaKx9MvqvKSz+I6gzwm14mTnop9zaz1ATbPtaTDgpI11Ymgwxd7FKCTdRUzP
PLt49LylDE8vsX16yBY5PD5bMRN2eltcWI0PMjZeU4bGrGDAGCFnEt8FGoeh7s2E
OTARE7b1qwSH64O0SjbHrt1wX0nCMI/kWutsgJtMNyejkd2oKWEzHXYBNV6a+hx4
kor40d3RbSMQGIvOYhJbItDe0F4oemnLxUciHmFqvHy1fTRgHrOma7NBBYKav1dq
7To3osO2c2gH2c8OqyQON3xubEG54frQRqad4Net6QR0eGeGTEUourgSrK6Ta/7q
+4aF7aAxVuybQsRPciw4VW/DBp40w9Og/GkPzhfrZKbZ5iDw6VobXtJvst7+6NUI
tppV2bl8Ovj9xLZO30WuOtYiUZ342pi0VOL+fC0gbfhtjVFop4PnrsuDQAE45IIG
VbT0rAq7JBg+20N2iP0yEoQmzSKT4jzKaBVhSbQvM9UQdmyeKo4yY0q/Ejo99Wi0
MZ9FdBE6yqB+vjlyjLcrO4AVQDsvPu3ql1hjud/MUiQHSEyytNT4h+Pdf5gHQ7B4
AqEwmnpBG2bDv3CaaZfrDLICoXak/yByglpH0mfmmyhLC+6xc9eUVF0DvFSvUn/k
K39J7bu6Za5FxTsHzKjvfW5OCvs4WGLjBJQmgxsEQfQj3fjv0LLlsp4wi9XUNrVv
osNBrvKSiUE2VfgTnUYqhy5xJgj8T/ky2rznYecchONQg1DY6n8ggd2gYjVPGghi
CFFJTtZk7Jjf8N6b0y8mS1bS/H9CIu7uS6LMO8F9VVvI0BjwVL+NylyBJIcuMnNp
l20LTWCEK1Qs+l7HIKn37EdufFPbmChcgGIL58NaL5pUnEA4qaRjCwYJpgt/fXSO
QifVSTpJSMLqAaeMt8weyFjg2fiDRJ9AAFiuAlBJ0KsuWgrKiP3DEt5yfN9iUGu3
7rlNDb6uUEj6kFkragZg/tEjwcn2L3OVf+zWtsquRVH6ZxVCRacRTZfUk9YXD3g0
8DwKAw0Y8Lk0ckUll3WYYTMP84mFYvFW3mpfMMD6AxgHz8yMQYGmGv4/iD7qzT1L
jIOZs9NFSvM+y08+9Zx5HG4UIGQ3Li0COJ4yrIyX6yy5hXXku7Ll4NJHNfNrV6mF
RUKj8zXHFz/GssWSTxEAsR75bx5A6X1pGtbwnR8NsnFx/xJc/G0BOKZl7xuSX4mj
t1hf/1xjaa0e436egI1UzpwDZXyWzkSvl2k1FFDJ+Ojd3w5qiLvkVrgz7fLK1vMB
NRzxfxzGlRLLARC5HHDfc5xKDw8jCPQWu6qo2pr7ZHEFKDNHpxprzqLxFuevmoHh
IeYwnW5Xqq2aqelHPxG/bQBDYaZOPT/xLPK1K7ml7FXp46vTDrTyz57G4Xr9pWBp
SU05qw6I5jqKYkGfnIR/pKzfnNCxie2c8qkOXN/vjW5u2QDPrYmHL7Y0LqQEuiCu
2W4mA7jgaR+gXJmNkMf5vlSzVITDHig/yeZsVPnl01RIP97vGYaKwf+oXNkJUZpV
dxueLz648TgA6osCBSbN7E5lpNoaPByaxm/JSzm17nqiiU1/ljY1m6+IVbGKY4Ik
L1yJkEeeozFne0gWedwWo1GFEVoK2+mCpozHOw3m5S/O0XcLxn5bSBHTvplNgsUs
D44Am54Jj94WMRiQnV7o+NuYZhZWdzFF6XUNItVaKCvTJvxCAlPTTfu9PW/iiqjK
uILBevxI2a5R5bvdHUwQcxVwsEhAmFjp0p+1PCdcRqxxZhV6NzYtjFfmNZ7/4Jm4
bXQpDXAomTOfcL5PuLk00rpV6t3HcicF8I7DwCB5EuIAdeH3WUTpWvlmy47n6ZPv
iWlQeRhxIGzcBnWqLbXhCrKoeChpgyjjURM3FMPNMPuT+BEbg8LpWJ536wat5RqO
tESA3eggktTtnYZc3ntuY/LsLa9DadzLBOq4Go+2XwedcJ63XRLqXMaFeDI2zgOd
tyd+pB6SmwMJQcrOjrpgtoGKA9B/asHod0lPGMIFLc1XRELdvdixnofRsJdwK9RZ
z9O8GqYoOE3zsyeIaN+rckTbv5hFlG1AvkkYDyNsb+Y7gVf424Nrbhbcfl39HeL4
07dzccDhm80XB05+tgio1tCfo9/kEMWVE/zK484ndWKAvknThn7/OQyQkIYGtwhz
rmUgmDaMAOpSjjgzEZLstZAMylXxln6pwRbl1+vc/eI0OuAsiyBQ5VXbaq87zIfZ
p8ib5I9O/C+dXkIihgaeRQ/yPwMy9PGddJSI/w5h4D40i49jlFhYnBhFCTmSdX6b
5eteG4UgTJ+TWQ1xmWhYK1EFH5qjDT14eHTdh1ToGRoc0bIaYNJ1eLxIxaVAyJHq
E2ADTcJ1r0+2ooSlbySxPGWw1PCwRrLMloZJvQrGfXUF2IlIQgdP7ZLhSa1bjYAb
JrFUjabmQYKHWP4Bya3CgjThgq8v6JMInu3fX0Xd63UIaxyNfFVKliSvTPBcDyy1
hxbAPOdJwtlA0qrVbNAFWkLUlVarR1lveHmo0PzLKu7IF33p6VfTm75eClU8LBgX
7atGri/QNmRxjWyiV3+dC1+0xcQdQSjCo76yZBiZ8sNeh+GHaa+LZKH43eWsNR4Z
Tzotpd4aK0wtct6gEwmQKhv2M5yEWyL2OYcDQDNdR6VNOoC2vBDI1KPPKPDFuJcK
6h2ukfM8CVdgfi2uzO19er8QFeRMPjStGvyc+PK+UDizv3iUGIqQNlf5A0ikfQqH
pYRi2WCan1mU4TZHWuL8jIfJdlgx4WiZb+EZxt8ZErqgqHxa5rgi6Z0Wj3clElOS
qhI69doKLP4izMrK4uiMo4I34eiUNy+lx2OZmdm/NLnbkWAIJ1W1ct69zOLRLO10
KmfVQWr6/nLv8E/TVydiFRKD8CnPr+LYk3+aE987f5jZIaGn6O5mHXnnUjhVPull
pGARlw/h4r+xYhYeNfzv4tEDBU9zt99n9oA1+4HE//GNonMBXUeyerevjgPki1TL
Ldc6mK8/O/IbHxdVHHmt4brox2Mx6EdDPgMgbP27zWfXgu0/kjK0YGY+sze4BjA9
azpyNW0p8+vR8cf15FLoUOQR2lFpoBdXXsrYMyGHhsvhGyHi3RTqJeJ0LGX5r6S1
PrmoEqcgZKB3W2+kwrtQa95/Kr6D7HMfIX0fqoBol7ar4BljkLVzPLb4DuOrz0Ey
sQEV1OSAI9Nzn0u0y9Me5b1e4nEJyL8/bkOzdRSSEN17aHVXNAbZVeu2YFZo2SHP
+4Rj/0XWwaKcm58LsHaKMe4zh+UzbbvB9tEyVtxAtZuRJZr1PL1NFf8dOqtBroaR
i8G/+s1Kiz6CBsKuBvhcsliqBOFf4MgqCoDeeT8FTIBh8G5EvSRElbT7ltyI7Nrv
RH0DQl+5+FMiz/91EVNUs9GnwOWnIQPkWZ32ZbZA5SJBviqrlT3jkfoFcV0t219P
Ao2V8lJx6uigCnFFfUIvbG54uFjfNodODY6tMhM7bGkE2fQLaQyQbqDyrPaC/3Oh
t9koBJ1QGJyho1MhHY3mMd+/7FZx2/V/4Q35L2yU4dViY6uR7jTaJIZ2oJr6plNE
wSSxr2Y1vmo+kXMmUSX9aBfuHhHgcbrqg5ip4KNCJXwSUS+C3mhrOQQCj2sNgBZV
SXquAIZKeCp+UOfc6zjHMhH1zaYq+zVSMayIwqYWH1hrSyasd1pqVIDVBpYUS9+R
vjw2j65kh9Gk3IB1fq1GNp1iqlFfBw20t52oBnD7VR8ERrA7Senm1WAKepo+Ut1x
KObCKZnVGEpJqiRZ0NzAZFAMwvhf8kdRY7WMuFLrB+a0UTzQAaTHAe78nDlsTPEr
p/cUPVPR42D+nvsI3XcNd2R2NB6ApGk2q5m6RmKbnolFgbLEoI0uB0lz2JladQwp
D7My4OzzLLe3COvcJSe/GTjXK1Tut8ynHU7Q/gkEtNSUXgrTs6gd99LDvX/RtCz8
nIPn4N3fGbqe7xDriJ0or3jzRGM6r1tD0Vc1XaSEjSfQHF/8MNzVO8AngVzRsDlO
hkcrKYrr5anG4W2M0CjobKwlBB9pi+wu4csO4AjyNuCazXn5ywEh8g4Se+7AZjYc
rD24bAzGw4G2IhnhHSZZz7uR52O06NRNhp8qDVrqhdKgAM0LQlsK9YxGnfECJNf0
/TzwmFNLbEfzFpAfjThVRSuQFvnhpsqMebnHel281osCz7KEHq2IG2Zlbaa75gU9
vW6PUeE/DVjphSr8ApPGSa2sBlSYlGZ0+p7gkaOmQ8hh1M5n6nh5loTVzfFhNzvb
X07Yhq9HQmNJTZF1wYjkF1UIgdaK0rn1bbH6ZyMkk+qKg0bZWgNKj7P8qmw44fen
jQwTV24P4kF6Rg6uvUd69K0vckjCfEHNWeF8GRugKoXuT51eigOT6oU2pusL6t3m
svyHVP7JfcA/4neCN3sFfWeiqoEtwENGsTGhYfRAwj7mVmP42IYc17YF8Rp7MnbA
TZ/fMc6wJIUJ8hb0zy9utZ2iZNwwlp20/Qfhw8KUK0Ioet8FzXUUIPUKtArKq8/9
p6AsHrhi5Q+zgLJs81UY2aXb4jkLjv5KJtDByurRru9V3TjPkL1iKUAN0qo8h7EO
9NlL5TpOmV/khFAlWeHSPLxR7tNi2E7/8H2JgRiM9Em5CLA+RTfSFa3hmgm16/xe
ofs7tC2YmrfaaVYRP53U/M+ScJVZGuh9qqElzgxcRdnKN5NEY5rij0AC91o1NIt1
eAE6T+d/2p2Pa3I+Jn2YDdfVGPnQ3WxA53NeaYgfG8kFfKmjlwLTLYEYzTb8s770
BObAVYkctWqDO+F5wuEn17t1x5MhieihlU4x3qbJDubkjzKsRNxmJyLYAVuyGFct
8+bkJRU3cgJPg/A0PuJUDyInCNrWLdQu7Ntmxwo5zxHiYjSqG30I8IA8Nb5f6Vbr
iihn1vrRIZkdl6HMBnXZBZUPD4QjqsMemTWx63MxNr0ogoN45Bswt47/304xgtGT
FHarXeu/QrHPjroFHQ33hPdbYkxWEvYTvnqu6eoPpr7DCshl6ddvXTFifZbXQHWC
nNUwdW63tYuFSw3+7Y8xJBzmQY//9p8wJtEJmpx0p0SLbMXr+5N7aoIH0v1Rvbb1
3bNeTdD4mlOVOc9NI2wmlYRCfT1y26Q2g/03wYgpDdPywoRhQxR0TenXtK5qc3SR
MPuHNsTy6OZW6QMw9/Ve/DIYSYdom/LeU0jKRdpjnuThVokU9FoanWCMbUJuDoDf
RXOMYN5ozhXIuyM+66PhPS1jfKjpYI7GPeDcF0iggeRfFlk5uBv2ksHONYnM/iiG
IqMIAq+B+JekkTaVl0ZdypAkL4pmQjoFoEnU2FH0iskBehVQRAicCnT1YbqBXdIO
gVCYlxrhpNjn4VaGVGvUo3ceD5HWI0YMGu7Ewa3sMwTVmLD+oJglPodgOLrroJRX
B4NKPtJG51iiv1U/a896M8Gm2GvdGsdR0iquN3UVPuGLXKFYgKsB4nVCQpK1Xrj1
QQVZfYCAklOhtKCHBXUOxVv+4yzPWGnB+uvfgmjvRJsnHlXuZ8kPxtgcrLhJAivz
KI6Y4dkdMLsC6Kxgevz706X8YKe6d/jD8lUcoiq262Oe7ouJkA7iZtdxONCp4ynr
ovpsmKQ2HzPg3byM2SAIdE7OWYX+fmiW8aQzbpbFXcMwA9PE6MV8Nk0himOgdhXJ
zjmhvkWsTK3fsmsyodxur+twFaP7vFOQ0nYRvzRPanbef355q35EkvhEhl4HOhNg
W49WAR8d+6WNXRQpB6aWkvpSiDmzl4oJtmPwkL+dWzffkqU6UDH44WuGeSqOMKJw
7yDPVYViobCggb1MAhQu8L0Df/yXIlVSmmfk3WiEA+HPO9YKzBC/GC+cC+kwpDkC
tlvGxIxogZzfzkXp3EugZxkEdmnvZqnlHPDe83KiBq/usGVfiKqcK7ehpZDUWZG+
xtADXI/m8iDVrA54Fn3Ni26vXv9fUh8ZNYbWaGwaZdLUelWEGcpeRoSgegBp8D4/
ezrT58RgDCpnBfVs+MLASmJGw7NnnkEPZU6HkbXqFHh8pJdV24m/mQXHPJnj9kPq
SzFC8sh2pnz6yfoae09i+rSqT5MJuZZnkxy1dQAD8WdZrRP0g7IEVEb2dcWAIdwX
YbDSdqowGly+S3ldIuP/rFz9czPWR634HNkWVwpVjgO1lNt3qJ+MIVRge5gvd03W
cDPlfmypYXQOqmKfAGayMgghq9SwQOkxbLx4Ie/MexxHhlTipJxlj5/tnp3aFCgx
1Pt7B46QIXML/CAYxmcNls+2t49FEjAKeANZIO7o8YGNBSjP9CjX2kjNtImGmj11
y5YZELN9CWw+js8xot5UE72aIkTtV8phvbeyUZQHDtx2ab8+ApQAwFTWomu8Z9hr
r7nEntmHI6tWuE1e5eXp3lY2eTooUUHQXHJmdJxDYiOfOdka3/IEcQIrX78IDt3r
Yyp64Rf2B3P4pw3qKoWQWPdeKrWOwj4R0q01ZQHdTujex9hkoxjvTNnm2MMCB7ri
iLPNdItau4mofi3FCzVg4zmbiypxxz9vq9H1gAaY6+f4lvG6pQejYPzzYaG9FLpN
F2j74tKvAyyXYciPPkUdkaN8GIlXCsVufwBdP8SBl4g2/myrmNRPbMLsiPXF5IxJ
ShIW3YA9CA3ruIxStPyAp8K9OKkp3I36qajbpEAQ2px43fh1HEbg2woDW5/dksjU
37DLsBFlgZW7XtCV4/aJtLycqp4xlLchIVnEji2hQRATWcYNn4yT66JoH5xQX9o0
7p9MjduRfBSP8GnFVINMskiwYHyYw26vDqo2s2H+cmh2UhrwfnLN8IAkHu9c9vHV
u9/r2Eh1vi2BU4CiIFLXDZx6jrGRia/ebqZCVABF6LTm/AFpBE5aS2+Ff7Q9xjge
4kKN5x40lgQx/MIomm4vrahUdqvZYK3lxH8+bOMsOvEYWe5S1BY9Ed0BTa8cLsW+
Z91r5M8SxhLoJD2Fg9/MJPAdzxVQbfMR+JX4exErcDMM0+dpxhI/61HIKM37FwIn
txxs+X0hyteYShRu2+Qcj8OV2DokcExg293ggr28+zgAq77JH+cS45rv+dqO3TyD
pyvHzoEZhubN12N+s0Lbd0cSjhGkzgLpkPCNuI6oMHF2P8KEP7fJNotZyy8FZulS
fHGpZD59pWLXLQPr7ORsXLPtU95WD+YrLOzq1Ku6ENAy2+sxN7TD1YMC/DRMhbuV
y9uiwHXPSVEtd81dtT9aQJPYG0QH6hcmEkVEocfg8kZghwHIOR3dt3VRbl2+/Le6
Jv+v6zV7GxrAt0ESi6Drw4HZ2EbE2A8V2PUOYk0fBfqAT3iDdCivmRZi9D5QeMmG
6714BBeufOKHvprSVZlVa0Ueo9X+HJfb+2B9kv+mzCcZ/L9HiLKIpvS6KYimFkmf
D48QfcEAvVLjVh1nDK058UB64O/8rxTfGBDduHywsCS+p5HY3dCCLn3zKUIbGqIA
X5+5YwCZlkXT/37ZB0V24mblE3n4WZJarXdWhhM8fT94t78ldOW2P8vH6JIfM7yc
ILY++Wi8wMOy4zYvFD1y7hp3KJdkFEYD7l5ras3S3X1RuFfSvpafJ94LZrhHNHtN
UQw5TWreteMWKpewtWFM2HqKC7O8ihASzIU0KrBI46IdA8u97f3QJrplHcCmjofQ
IAy5z59wpIrcwn87GCQlJjX5YJljVV5O8DlMZTBwvlyUYdWuhxgkGqVVAhaLnxUj
RuaKfKv2ezQsvP49rj9p/UV2mkiayJfzcjEAUphDOKdJWLkdmz4b9xips2fAcGYH
yR5k/f68C/sjFnmPmmVhDxr6F0VnjxEEzoKQCCc4F0J8SVV3mWzyI93yL514P19V
Y7g3woCAuITl9mjm1GNKKVwi9RW7GZi3bOF3VVMggFEliRE0GzMDlOQuLbG9mZ4F
cWNEVz5JFZk7hM73FowHgjsLPkzi4nRySaFkDNCqriyOj1N8HdPjEJBNXltjYJGD
3R/RCHUYgoM8EEI8Ss5BDClWHk8ZQNX8hcjx2qSaGwBLWSQqlTTBzpA/XLHY/fxu
GHFdmlm0WsvotUjGmu/XwlhKYyE5u4s0AgN58fx35ZXBlGn8/WERtT9MjwsrU7/V
uO1Gy7+pVs0LNhF+cQVycLto3E6SCTcJLVSDhz0YwjeXY7jcEjzyycKneCkXNJLe
57qOx7FJCtJGUFm9Pd3lWavUPN7BjqMmgNufLQHqtud0TxTXBOiKjf6YImwWRm7W
TmJfb7I/lHDoBe/78u7ixIktsBfMgMEAMP2+FgD0XBlKdY3hLUgzyUrFU2ObON2+
xzSvDgIdzFT7jnmgSCtxLsUUUlXr5jgrTkSvceoN/Zs9OMzWrIhqfOTzZnIwISux
biOKdFYm/lurN9400CfPtCbDlfd61DKLhaJ578t5Mb8EyLao3pniGYerhWVRXfWa
YObtU+iKyEh5Wv8GcIFkHW4+E+qYc6V9UThTywp836pTJNUjCpya6F4LqjtHm+eA
N3N3SH1YHaxCzf83qRyjqSSU7BSSmHExlo3ZxRhQ3Q6mp+SLNIO0HljUYzgYIx6G
lxvYdQFV2Awv/LhjNX3L6r0YT6F8iV5ujXJm6fXe8hA2LZstEquK2m+LFliEkXRa
QtDGdy0FcbGRQ8p5vx5UiwuFG0CerRo8MEFSPStUMIgMsF3b21XdQHapujAvWZlc
LAdqNV0gBnrm06oq6uLx9uq/JCV0KtCoK9WOFkkvP5F6/9mkcMEbOcjnA/96l3EC
XYILjTmUqPZIldYn6+XPPD7w6MrDb5XrQ6nL8SmsqKKQATequsQZw1J0h1ZBG1d9
+FFe2zu8gShLJWfzkpKMgYhGczzWN/JZL2TCSPUslEt0sbYuUIWasWMJ4WxwBiSI
FoKVyy55/NboNjAQ4yfjmS+kxtsFqeSyXZafy5LyUE74SUFpuJY3GL+fa5zy8N4C
Yk7jDJmbIkyAinxPbkemigVLaIvwaL7HssetmCLB5X2W6T/+aQPZi0imCE8y6jco
hGi1F38Q0Qkyi+B7Q9e7nl/WcS3utfXfr529rGv7FhzGvpIN3zX74LG8GgiVxpuy
tmhvWw2l3zPTjHgPLsnSNSxGbqIoL0Ir66AMOj16/LXyG8UVsYhZ3+t5wXeEBSAk
rJ0nSxkHjat7bbA/LGAeyJUOu1qVCP1BfQcjvNMVKHe5Q592b1bPLC/yBH8aY5Ce
iImSAtkiUzImXiwAmp1CEwwYlGtoWxyt6XLrhalAMYnqNkFLb1wLuYL9QOZsQcvJ
MxRG85JKuFjU1khm1+SnpjptrVhnMUOehX5AO4o6kpDJr7ubF0QRzoWVIqQ/ofd3
+NneijlWk+V3Fg40u6/GmBlnjDjC7Jq0QJe2c1+nHMsT3OL4ZsX7y68tJZU1LrI5
sytw0Y9WVTw0t9acejwp1j1BtnZssYZEBVvYdIxZ0FPOsq3lMhchXP5Xk15lnJlx
rR3ABJhuYuw7ANjxq6M9EeT0HvkUwGKVbuvAxMGWq/zdzSLWHzz/CMquFfhCC5Wz
VQQt7uF9WBo99bfdxu6A8rnNkhPZppl69EVnRQXCbvenoDqn9AH9ZiDEBQ3hq/Ce
T9DLodcmnCOPA87MaBB5zUE0+n7C91fK/fehSo1HsX4RqTyQNrn90F0hVTLQP/IV
2oL5zJd27AqwH7eWMjWEfPL5Mx3sRdai4FXm/7wZ9JTL1dExU2JOpPdsmj4Q40xV
Mf/xQmzeH7r0EnVLmlfZPnrOBrJtX5ynobu8qcYKm5GX1Dbm0tumXzpbFJaPHr+4
jGHjrik+vKSMtMUO4c4Q+XYEEol1Mp2f3mcWO/htkg3s/EdrJsCD6gwByrIarGzQ
+hPNoC3C/h4FPszqDZNUiS/K0mLoDePqOm2boFPE2AjZyI0DOvsv8JC6Dk2MxZ3N
vQzoavblSlgzMFl6t6Sj3EEg1O7F5LiJUmkhh5ri4HwKIa0xZti5jNi/dQBpi09P
k++iRqipp/3dPOSUzc9V9KZOLQfa08feazTxRKSg/EX+Qt9sHg2sLY1V+GnZtxbW
WgAXx+2vtfRonaN4ML/VnvHKf/MCJvIyKICPSoLLs8LXDVqSc1HIGKcdKOa8oWzv
K2fH3Ymi2OM3zEdkriAKOOgSgp40sZxeIGeTORbBPgTAPOAjY4xQv3RIDTz4ZIgf
ikkuUn5rDpp19mzW+5aKkvDl8+o686CkxCEV7GG4pGCotqJmB4VTdIx2yuTCH43n
ZZIFlUx4GvZwm3cO2AYV14VwOlpD4u6TT+gPwwbNKRte2NUZylUFU2gCLD2oJshw
nzNmuEvAr7dLH4fki/YGMlqLrpS8o0l7ckEonoSH8JyLNbPaGuvRiTzUAdnzrrul
3AvmPI4LYU+qaeXz1gwPB2ci9W9nfkrens8TTYhx6opZF+6ebOzyKU++e3I9E25j
x5rROpSpba1SHlKo7wtVp8mArcVxUhdtZNEbj5nmQFzBmW6/ZUL9Mech4YEWgGfo
VbLoWvZPMGeuyAY/b1ks+z3OXNpGHsyZ5o294r/PhG+SdjRyxvSOg0TcG0iO1zT4
KWXDqfJFdhXNdrObQKNTj+lwXpqi/IzOzK0PIqpm9cCSKTxhUswuYLfaQBu7WwJS
bzUpZKki32L/BZgH3//UgSSCz0iql5GrOT7i8xTIrp6pIg0p1HihpD5qBbg60tDX
rD/0JTqZIReG2mlrNeOMZ6ZMZjByXYgLbqgI2rfAoBGoLkNKJI8+D8mIlcjWkedV
3aKqdWzPrFRnRtVE3zfrW+pegeClYODDvjDVOHznwGqiNZjDi/S6mzM5l9Ui9PAs
LfyLioseHG1zjVFqLLaeTqkProCZWc1/Nf38TSB+R8D/aJ9DGnUtCcuvsB9PUif1
9TDBTnc/3v3Lhkz1v3/wj3iboWRKnsz/SWdqQrSD+4lMOvMyreY6uOjRxyt9ZRvE
atRdoysPYIKqQUrGN1pUrnRW2GzlMnWvIlnB+uNsLBiWDOQ1eA79edAXZG4FU/hD
NxeULxm7o8hUmvdnLlzIy9S03Swqf2iv1MbzSUZw58P5nP73kgGAL3jG4+zvzagn
d4TBI7E4EEofsstH35L0BJzS4zKhPM0fXjb8VrlDQUUhT5367bA2YlnrHMurOSxv
DOywNKrDwhZz2WsnTu8MsCmOeg7eXM+yAo0XN1pbF/DVP3CJvV2AhekaVD6/AMIE
DAzoXPybVannSCD+pE8TfTHT7wBaDdPzlkWAG/0PIrrlXOH3spy7ALqStUGVc4ur
/0/xsDjTxO43ceTjJBHF68R/Wo4WP7MUjr2LeY13Qo8kJvinKNl8eMVgyMYWG768
EW+z/PyGfZKdMV5YCrbPdqX6lfjM6LbTRF6c7BaQG+pv6I7gv2rKiLfeTR+XhxiK
qrlArnCvVUdDgfkVq5sXOBBD2qxMJc0D8EeSLZ0iaPXXX+86ZQ3qqo8rjW9lewad
5QoeK6PDgTfST9qL48n+OVA7Clpf4anxsCj7EcJl9J/El9hkz7RLDU5U/nlgahTG
HyYlwcXWyQ+dH6fhJ60mGawHFTUmwHNEaKbGsOpv+7yg8zzH7s2QPZFiILy4jZZO
LLX56iyl6fnUIqPhSrd/O5pGda5vwT3GTUvr4JTff8zsSxMMDpBWQei2VzA84j5i
S7CCxUAk6hG443DamyLo/zk9PRYuZAoDogzsEPM9fahswRpm6e9vm+YzQIUKnmsz
xe1VHXZfc+FdkBMshcGZoMvGYskmZcgV6ozmQV7xQXftLDB0gOjsNvIWTitDZdzV
Iq01sgw7lbra9zsX2YLOO1aS0OZ9JwgCVAqAdxjkALhS7z3JwuBB9ZZcCPBTnt4d
lNrf/TH1Kl+UyjRLv/9+jtDgGMoKjM7FPYnNVwo6EoHI6PeeBFcq1w53r7CXqSgF
tauOqV/cmED/kNctqwOUW1nIeYpOQgkhXGT0bbySJM84jTB4C6KWe6w6piUmsCSW
52eJ18VVwjcLZ4Ohv3U6EqPLNrSf+LMiT0hI8sLOSc9OOi6NHnsc6dKgRTrm4/c6
1yyccYMFuK5O5mxRGus8sq2U6J53cr2qBYsxyddxGjr6q8Vo4DXdYPooREEQ0mQE
rLBzFWuhc9A+OcWklLJoE5GGimD5i5/l/nfMVgbDqkjwbyvcjrRgh8ml9gHZA+mO
uE2DXEsQqny7kGAhMxWe2t8hei1U5G+EQU65q7ECIBwbLC/2XoDK7NpntMfkIywG
vo65rGZuM2mf/nlHIWgVKyO0u5qEwjmhb1K2/PSGWBB7k4EcPeUxE+oVyMx4p4wN
Gkct3D2psUzlLvXHhChkYmpZgeCCXzPiVPFhsjGw7ZbxN6mWJ93yIXhwzb0FQgDb
Vk/zUiHup4QPSF71f56laqxtMxJ8P7qFJuCxXOZCJ9+2DKwrJJA+Pv99WzNKdfQp
W5akRxrdrpIqdltVL01Xk/CpxsQmos+psXeCpIy/VCrBmPsssJsorSDqRjVS6rZf
u03myJCQFmFB80LbI6Gc1703yf8CSVxyH2Uwc7eakqki30Zk3I7cAe7+pkW4LUWU
w2uxeDYVX70LZEYlgqulKCmNnVlLak5O0UnKRnU0chAUDrDoETqV3qGtnr7jFgTc
fxudgtZO73csahJwZmZUL1pkw5R3A1U1EXIkI0I1AxnIYTW7JYuUKKcwd/TXA9E5
xnblltiVpDYpcfGu9AQT3/DjJJKPb5ilqywqnu83zC3p0dJSfNS5EOSMG8FC2Kg5
jgXXkkXD0bVbCcj9lQ//GYUiIX/+BeDVgg9AvPJs9DCOaANk4ONVvzFK5SigogSV
KUofqxvC6edv4CT6jbGLn7AogzLqP9QJsqfbzLGcU2R1PHYUxD880lMPLoKuUniS
qMY0rFkGj6BNC8zOcfZuXmx3P806taoEWWpJ6jfsyveCp2iPeYiHVHS0SQOWG2/p
cLd+oTpjvPczPph2SakKQxZHePYp8HhnUHaVO6RJhd9gvRe+DyIO6k/E7rgwR4d1
pxZFrUFhNGNodqJYDg62zj5zfkZc7btV4KvmNoiujPYWchrkbwokE4FPF/Lw6UfW
kZIS0bL3T0xLF/3N2N+xJsyWvg+cG20UkezApwz2A2TYrvDASyTBE3L2gcx5czt4
IbBW7y7ctVXRbGYaSptPGh/amw0wo8VNAZ//dhGJZBZXc63OPT9mEmikHkjCfF1u
P3L7RwN6C2wunZHx2j1H7LGQ4mVrOKnBaF6fuaN2x/dfU4OQJThs9pL1etr/sIHJ
i2SpCG1PW6pVCN3ePHvNaCDDX0CSeTnR82h8rbYOnBQiVNbgSdiHDCTOQqGshvfK
UgWnuQuyNcyWh7wILTQ2/QmomMUSRy4e1ieP48Hp4LIf1D37a0pWpIdEm8YSk0IE
VAeEpO7JiUhyoA8yfli0PBTtsu+comZisIwSFtgpeRFc7yuxWMDot2PvxsdBOrri
SZRqigAEUb0WLgmj69ZdbuAv3kkfdIlztfZrGujqcd3i0GFc1bCaudHnrBQdQA6y
b6BShFroHebxFUO9PE06MBxZAeg16patw2K0BPG7MR4kH0T2fXp3t9Ukt2yw3hdv
VkTIUrSm39clp/AsZ8nTRm0AqP353EfTMRHr4M82xLFqP3+jcJfH1lXfjvX0PxbG
3UKg1Gj2DAPWEtrenj8HZ6f/WXYxE92JpwbQ2c0HikZdk9yJC1wlXEbpKslHV5zQ
jTf/eFx0iR3DNXkBhdk0smtiUwnQhe8vwxBD21n7Kow6D+s4rO8EXeRJhV5uiBzx
6S+GCvySwdLQDA6RmiktSSW9G1Ou85kKGUPngxxT/IOjZbWnWDZhdwDkAu9ItsCw
8f5LqRFSR4T3goWSMLnpatcCGRRm8NKDIn20iXz1YcoEMAr6LWsNBT2MHGNIiSVk
R2YOfB66zqE84/7NjjLgGTkJ+CllaoBJ49S5gqxy07077Q2mgez/vJH3jlCXW0TU
DMHJcAXHWyT5s3pb1qCgKIHAWnGMpo8m6NYgrSzi0B5MFJPM4Leo/O383LI9qdyf
QtQBe/88kIfh4OviDzCGGjaI9clbdSiiRPraZS51Wa/BJPFA2ctsik6yC0rq1sn0
K1eyZt0KrtLrggJ4mwJQIq9HcSVo4BwkOksOUKJpqUIMhZq7OzCM8rvfggyeoRcx
F6otTG7hL42HVRqunf+yH9eFBhk5OHMVgowCLqD2e4oT+wNvxH5CTwZy9ezpw7et
aJqPKaRjOSDsc4WQJx8T+89bklXX/JJ1xTAJKEfw10OTMz7MMr7vD+Pjc+W/3/7b
fWeaMSogkZ4NJBeezC3E4hYBhVtyNw0RFY84KEPFYQ2DQ+q140maW/1iI5Mzcoe5
cQqP+bjEjGeqTqenM+wKLfIItA3gHMZZz5f9TmFWM3JkJo+Na3xGqsrvJPzksxwf
V+3oUn5ZIS3EWJNFPqg4lh9JG8MjJxg8fSXaQO1QePzBmPPxibZC8ctgSk+czdjk
kVF9A/rVHh+5hwl4m/c3NB3fLNNWAryKaUPGGBmEBLgcG2Rh7BXsEoLGrBJCCGTH
9DWcoSme9subeWNlkTgOY+sxaKcJhO9zPIsKHFtTylSR/OVNHqnL8C+rfBF5E7VT
jeQ0QLq/ci682muN6mEKk2Sc0iLGXPrl6foBwewG/6yn6flcsZh+NWvtMVhcpukw
oRipR2fHl8bwXEsjMHWYAI/VPhF0GG4pSqzJBP3AGOBX8xJk7OviY3p10oIIjH2K
hhvfp2oYDurLivwcQ878OTCPtFcLa7hsktweP3Y3kv9iK+WCFDHmR/YRmLzn0WPZ
ijGT1jX2KeeHShEgVLSG6nksZlXBOZu+6Pbp0u6D6gx42YoIGba0qOIp31qZaMLb
L6JVgtPP0PFsZgKnsFc5aUn4PKFrZtzB5WzPLMSHZuYUKlLzvcD51ANiRaazyNim
K1uLKzWOIPFRayYJvDnPR/8qDq8APQ5pmQBLnIpyaPwPWKM0kdBWyzVJPWNnFC1m
eEfEuykVhpbhdTQTK4IxUSayRBKQxjAcp+vcr0vFUGPKRClfbs/AfFyJFXaJEJaz
d8tAyBbNC976jFxF/Dy34h8FNSx+Vw7CTzqVt86VP4FOuYLNlp3hJ1lT++CpdV5+
5rBqlmSZ9E9NZpA8PsKFlc4FssGALwe3kiTQSBAwNREQgxtnCwEWJoc6StoTkLec
kDY9oqkALBpF+F+F5Ht/bNGGD8UIattdiluSDWhOFwdD/4XhSQqjLo+zdCpFxyiD
M3mgLRjFX1nui3TGDBJn/c58wWO+qKy8Jke0j6Yb2buSDgl2H1TpMjRHcD+UZyDW
kEm9HUX7wny4izkA7hNltDYI+Lv0lhWs6YVbmMzEynrRlQAA35XeFYX3wgaLdtDv
B3ga1TsOUOp1MKFBOQbJ8Vz++f6eqfWQAOkIlsfrhVjsb4Y+3FYXcQFsA7lmtTTn
Ro9o2r59Utl+ekRb+hCKjMDctZu7DV66cJf9obOzyIcXRZ2btRHm4an3Blx0edih
BXnZFEgyqCeecsBV9wze94L7YRWnkQSz6WT+nB8wPM4eQ84bos2htm9Dvth75jV5
0ctNQUkqLx1EpFkZVaw6h62Y0ARnm0BgZ40NIvJv/1sUqVoCR8O0QcDdJe5ieSLi
/Cp7ZvF0RABHha3XWHks5aFBlIfYf8Ertwk1EaucxF92yJoAc4P1sctP96ml05JK
qeW08z1PrRQr1+c4N/AL73N/2sPL5bzR5rLwHqaE4wabpLvrKz+sz8T2fwH4Me4x
n5nNDki+yRdX/5Whlh5NtI9JP8GVWGlhkbf83LrA3ip1rtZqejMeMJ/o4AEo+Neo
Po8v+9hQE/pMAnNFG08hvAYPdAFdmMXDflPSr3j07Qxpt8SEo6lZoJIemgHtf8lR
BGHyjvw2NAf7mgQSBpzqu5a6KldF2YGeF/2tn4wURcVxU+qFdGeScUk7d5i4KfND
5Yw+Npjz1h+H7iHE4jiwRQBJmFAg/a6nKveeOlx8+rm7dN4Q0obbVUE1ihXG2ieb
Ds+jLLABM+D+J4koukjUJo0wppeGuSsUViVqPlIcpTrC2co3VvWSDK3kmVP98QQg
g+JLBZRQhRw+KGQ5pbUtOqnJ8navf3MfIL8sSgS0bcbhyhJ3EIQALOFtMqkKpYYp
wVN3TkZ02VLVc9d4hpHA/+PIMf9UDuIseS48PirKsAWBAvtAFTqT+FzKZnCbRQr4
y/YTYX9mEgdhlrMr5zREuV9XR2kQtlcVCOSUI0XLb8PhYK9fLmaxDlio33DYuNKA
L8/sZNu2O7MD8bgYsu5KOx2QjI0tS0rzI6R/AMaOPSlxRp8br2m861d9G9S4T3M6
tahzp5a5AqkfKhbzFLR92YKu6w20l1ccrtgzD68JIhABBKlTra8C5aZOLVri7hop
c2FFI/TqUVB+E9IL6BePtHKoJteyIoCZMEDdEPsjI7CkTuH5/lo4jfD19tbWnVBF
EzFJGzkRL9VyW1XFX+7x9dNLLZJdwu6Akn9ItaOVL3WAAce221SJeDJZaFv6HxVC
H79umTKSGeJjs9R23iphTquamDrDu21OUAo5qxNkec2Bd+lsEFvNFCZccBhNIsga
SPTek4lFxzOc1nFZG8heI+SqAEtb8z1Tq+rQcK1oyWcnCTPV/WKGCP0MExjjW0n6
m8c2XBw2POKMkgxmfn4SEsyjopYbX9fEnoSpOHds3I08+GeuimxiofZj4/Kv/57J
2a0pT+mmq0zFtiES/c7MdGjunUVktWYdBciZNgWDiGFlzyXkOBHTgj6+S+urTDp+
FbOAt7d6gXi+HmC0owqRO2hlnftO9njk4BalMKeiGsWanR/uLNYP//RF+d7LdENF
cvzEmU5N0xhlTBSW7aHuW0nq6G2JDKCGjrBNb9NqT1N9bhuubjhkMZeFMg9Zxuam
nmLC41h2tINhBImiYs0cqT6wc7KmvWlYpWRUCfpLWkQ8pPzJzrkAsB9cK4xSfAIi
4+bFMFFT0kkGZ7Apt48r5ygb7O30oXVCq0OS0RGfth77ja92EhA7eDCFpSSmC1PF
IhkPJOvpdqoe7Rg12KKoy0HA4uDCwqV++9mLJJpCFlry3/vQJT+xSarJuqEvsqON
baI6ASnIVnqw6MSHc9AilMlYJ0E+LMo00/iSQ8RE572z2hh/6dZlRzhJ5ATQbLv3
aNxLY6om6jEu9IrOpb7CV0g6mDy3ggn6AOYuq3SlsAbXzZe2P9Znagon9fLvbLNL
HEKaH60C5qfkNGvChAzYTM4vXRokkO1DJZZ5k2WfbGfVdZ6MSiWy0N/HpLKkprJc
FYZZQHw69YT8q7100kZ/PNfLQJP6VBWeThgXVfgRLbPvE9r2smuRLzYDpF4p/g5g
riwOEewSjdAYZHJjki8hYSwQf8BwzS7B+rBWdN0jCkc1TfT1kkMg+cy5sHIfCVgw
YIHvlFmexYL4WcbcaQFEolnqZaKoqqgrufVhnfQ0bHFW1A1a40jyjwxacy81/AHZ
NG67MM9uDMBb30mgz+BahiBweV3KdVCUmERQzpEoj56SgJVeKq993//bcYs3wVg7
nns+v7v0YC/QsqxRp2BUn8LscnYA/ce4QR3nnPpI2oRtG70G4M/4llsgJszlm3Yw
0uwi2GJCABAD4Y7RbDAP/VurEZDshDCE44+Z6crHB2tJmuWcxLuE0pJZu8wLDnGZ
Cb0DcxqxaTFjq/rweaSe9KaowmytUttSmrpDyww/pfDghRc0C6swtePwI0PpmVI/
1LUliCP3PLW7E/EjLGZXT9GmCBjGL47tSMNrQxqYCK1Amh1NkqQA6Ae2kOPefn7i
NXhre3k9NjiqIcEXySEqS4ObVAKFR3J606wZyXxUYvDInp0MhRVQUZTHiFvbALG5
o0R93I277aMKbkh0Sv3EXOplexBg07ruUQGErzH8E95KPYDPpJ0E8WeORuGpQUNt
ztMYEO9uzE/nKcBsz3mEbBgr4J7HOvGqWwNN/J3JdOYLFyAScrvmI+q9GkjL4dtX
1EDroiYlvRvsIPul1INfFUUISNc31xLw5nLs3V8idtCq8TZ173OsQ2tnhpByZsA+
wXhR8YngjrkNq98VgMHOOeTxEadUz4gejilcoCv+9cAeFHmcZlE4+WHo/+nHmeq3
oLsbg+12ZFsB6HVLbdL4W3nZsbpr/bce9g44TLk/LlPwqXKiW75Dj4qK6phAXmgz
Vh/GZNQMpC4uiY3/NkUwINm01Z+MGwZycLBBB8vUUgN966fEk5ysJNMBePVRTq0t
x0N/7HhKk/D04sPX0Ks+IsM+fSyqc54dX6YCAfVyVQDoGCD34KWNixLLd5ExX9wL
e+KH1ETUAUEq6u9gA4qiKQs0qwsUoO9ADzPkYszg7KJbpHlFD2wTuUkomH2FEDox
FU2eD4o4tqG/7ACmuz8dF1fbukybI+bElTzSOFjJCi7VIxU2nl6l2OWXb74AQbZR
ymPlm7Y5VqxgawUt2zzEF+0UuW8xtB7mAOzeKGC5zK+M0mg4EOAai9oZHKOfQRGO
+lYjZ9AucYomjGvkjPzbkGFnLKzwPThyw47n1sGmIXK/aupg6hJH7aT6NjFYt2/+
AZ1oGtzKTgsU0Hbv3CXy56hI9RJPvzH+M9BVwOIIgQqkHUs8HFgvKiiuke+LUj1r
/yPh4SvwzJ2+v9TlxVk7R/3R/Fdc50uPx3G5WXrHToWlUUZmTPT/rVvSHkSZYyrZ
R9yNIv1O8k1McjqMMEBevTFn2jd+xOREID38HJkHc51cHVR7Ho/bxHPKP3V3bCJ0
U6zIpFHlWBvLcUSwblqolld1Ib8veyoLb3DqSTsidv1qitQR1l5R4pV437d8EYTL
BxtZFU27BQ6JyJ/GbyYvMmJ3sujBUHEzY87pstM9o5JG6HoOFSmdR6sWFgLsTW8J
DMiBfgyd5KOi9q6Y7PtikUtmm0Plc5rYSPpnVYrI2bCqFMo/OT0NWnXIf+KUOdy7
UePeDw87USCRq8XHHbTBBPtWRLWZc23vd+l9HO3HNDVmw2BsAeGaWOpGwuoN04dj
0UAxP6XNVztCr8R6GXRWBO4H98HgB4DmPBp74qCqiS8kL/p6yt1sR9yjhzvL+e3v
bYeajy0VnMkAegna9xuiMn2Fis0DMhRPEDycfJQ/m+KOCpwXhRBbY/Y00IwvIs+F
K4Z6sBppqz1e8pkEMZmo1sp7CpCWWY1/ELN0YzcBVhaq+llT8OXky3vyV8VMmeSU
wNROuDMeKUpsjuLyCu6esivyj7b5P0zURrPyBuCB/pUnt3zEVE8y1G3LGcKxximW
TTYS2OCwSyZHBWT1qVrBFpVB/RC2ypfX0WlA4wP4RlK7OSfBBy2MSPEkDWsFVXc1
ioPgAeqld7nbLDcfvyRb/6YkUdwF67tk1A+S1SGfhSmqs4woOzhDNowmjbQgZlzf
Ge4tFcOQyOUFOLiHrQ/llb8hg5YQ2ApfSw7oaj/Rm6HXN9ToP9Llq0Qs3pjIgGDu
X5vYtzqN7jhlTanbM6xFatY8X1hd6v87yhq//HPfMRJ1Whpw70+5iH18fFBMRBmU
8zzhbwIn1Za+fWZubGTR21O/Nl+A6pqEPbPhk4cVLy4EzSG5Pba+u8+ORfwjeRc2
K42p7vr9wS+RNmMiUWEvCQSIg+P7dsW7aEGNccs4KhRLgjOIIXz5nBYyN4oEvhaz
3HygWkSWkP/Rd9CluePgN3pkdOYC+uq+Yw1sOoPF1OZjfPgt81af08axgnSc97+S
YrGwfMoAHb+YUbWMOTW8JGNUTf3t61Laf6LF0H9+kxnAunPMvxOglidaFyF88YCz
rqAUudPIO3hgvn3Czz8/cRgQ5Jwj7lROnr2tNZcrFQa158Di/SKb6WbEGV3C7xoG
ikpXJYQvEaxX6sxQOMyZK2IZS1Ak9OrPloNLYaRKm1S1uFvP/I6ZCizX+fysw8JC
YhKOYWj+4pW6vWlKxPYjrrboB3xk/3YNTGRNUiAJwQRk4Tbsd4KVUtEdkvYDgkxp
k0LBhMepRqcEcrYrGjmdd0BhUQjUiqJ0ICxG2Ka+sZ4Xg1MLfKi16IpAm1vr79Pf
lUXBsIvFV/mTcKYMeI1LRjBP2hWwQYm20u9DNKojECZNt5/Ewj6nkw/ZNYs1l20D
NFFa/j+hSzQaVveYI4nciLVECgp/TWBP4lOkkA//Rsya//UNYVjbTBgzpyM8JjLq
h6MxwsKvF5eSUpiubkKlbGJbOILm2fd0sJGcCiQHqu0m+USx8sZ3ECQxuSU/x/HJ
OmJtbK8FbqjCcqL2ow7IdPG4AsMSELBXidRoCan04JwWsCl70LhV+ouRkJwP2LzV
v05XQCDhy58wX9SAN3/uyq9OmeA9JU16v8DQ7VY040g4KZEhIlS3z6YEuEJcYpMI
9Ofpy5xpqu2yrEbS/c5qJcA9kJdayfrRvYu1dHIgDyHU+cobhdbFIKvxN2XpEITQ
yNHV8aWfM/LqLTpC8qRMllENgy2k+Nx5ShGkTFmHBR3iXw9FnaiHqhC1Hy2U5TiP
hJflESmlY1u5OJDcyeQWxK9hMEMX9r3ZsRGiScKoG6AINVUAzUes7trnoz9WpvA3
HsgQ+TBjGOWeGUJpfCBjhj1ED3O0Qk1zuHiiU4Z2cCVXy9OHIIV4t2P/eAcGGVxM
rjZRWLBC8+ZbYwtlUTbLe0nRcEkmihJxZwQiMAEihg5o0TZdp/4VoazUbtnG2/in
JFQoQ+Dpgv88ipFofn1kSdsB0PKKtL5v/1MW3SyUcYASqNoFaq65WF/xql+NrQ4y
68QcPaT7dAtaqyzcn0bC3Ft/4A3/57Mv677XfspGrFRkbriOSig77eEFerZQuAtG
F/sQLleV3AfuMZcEGcHbiXzaqkRX1ftb33LG7z//0HxoHnC4Gu7efxXdwTQK1ZKl
8oSt1ujcVNgPA+ZKH5SKD4tnWIPOinb5SFzx1rz30EOXt6Q0clMrDY6l+y8IV3Lz
gnvmL6lsvxPfkf/olG7rkiiF6BurKIHtcg4nRmUMbibpVdssF+1vlkHzkDZwp4xi
Lv56RJ/V9Ust4dorb29CH3kw8iTpzehasj6nuWM3kWtrTOxt2jJQE10Ao1DtwTvS
dOX/Cbl1pzTLq5fmYiquP8kjmxeK5zCrRRlWrHyeBKh0xhH+Dp1MXrpaCLEEliTI
QXBb25EbPNB9DGC4NBlTcD4d+B4I6AAibxGG5Oir4SKDwEGLGHlru0yb1JrHv4De
6ACVA/pXz40ySXwf28B4NT8eCHeiQyKHkHbs2wQrEnISEYNdK0T6xUWvCDU2nwPL
VIaELKL6k1fb/CnhDRS88HkdWNSDDDJdGFQI/9zJVXOmoKD5dfzq7/yYi/g32fWW
OePI0TP7rb6FUuNPb/9HKPice3bK7tPpwb1Jr5x+q86RA04jZL1bg0/qHdyjwA4/
6p0EqTVZrlXYxuoh6EA/hEkgaZyGY9KmYNGmuRXT0wH2aFxkqyYJWQ+2z/pRVXHb
ktN7mCwiNIneh0/sEMb5dIYtPwfIkyrZ8OuWw74K0zhaj/4CORvw2IS85KRRe0lS
xEU78v8bP1wFqUaONXOQ926thl8U+gvZlpwL+L41AdqPpI2VxHseQRO/dOKJqpS0
Oda4vWKe1pqjMcuLsVtTVcfRUFtInHNYdqQiRUNHm2eiKIXRRWqhV5BHy5DpTyUL
Sbw9S583eVRK5rJcIhFAvlmZZU3a40C1IO0RwS9J6WRiJWzkuMc5da3hbZGTdEit
U2CoM6WP6yWQlBXUEF/wzRhgNonUc10OiNJj+KajVbO2Sc5FCR6ofd3Cn6nVlkkK
bT7Gh+Mn6ydsP6+gMXpTqjY+AbziuZ9BIkiiOX0KD47LE2dYJmxEz2nT6DgDIpA7
nHznvW+5z2dTwlDVqHUrSgFl16reC3CiAmLDMrL8NSpZ98upBXvSdl/6idHbrC3O
ZwI/VdatvYpuu4XtGsGUpYP82K9STdORwgvmJdJyDjmuqERAFQwrc3KB34roYpyg
dgC8Uda3OcYMj+SqoIj2kFUpYZxM7m8AO9W37bvkqQgfwUs6U45INFuIxp8gMwtg
jPAe9Xpw3+ceI1wQgs75C70AY2bjycUNAhWPtfuSh3cqihA3pAYXA2JniLZXlArc
BTdABz8uAniMtmJpYJuKRzGv3vW3toBXLe/29gvFrYeVyLI10G3jVs6U6G0o0qBA
1Kbxl/Iv1npicL3jULh9qb1wmC3xEitzUQnOb9BPr12TPsomKjumEHK5bA1BavBW
fYIuv9ndKR0j8q/eH0LwOvA3nzh0hGbD08P1Pxs8vQx+Vo0mS4GNGmdpCex9zAfs
6odjZByQq2cxsl6U1lUxZLJEYSDJZDvwXFVMufYeRJOpYoBzd2J0Xit+kON7Ocu0
zj0LQlB9Hw0s8VrjHJ/aR7EET30hfqhGmJehT6+bl6JWupxk6dmgWgFN1W9oJQ+W
y7rZgqIDpFeGZuN0PqAgvo0MoIAuMOXeJs/XPLvhCUGFasf7Gy4sjFxnZQLYoeDx
oyhsAnqzI5FuyE3LadAlNwZPnES1ZDn9VWiLpMfv97lUh/gO1QxWnExoZ80t9IjW
Xk/s40kpt+Op97Fa3/DNodOf7JeQuFsVsc4VXjnzBRxgFspZE3efWngMxlGJ91Yv
viqlLITmH9TCCnDkvhGs/ixPRDqpg3XJDW3haNdnYL08ANWXXyEkg/ZsORo3/Sg1
EPsw8rV6kA5nuFu4ITyKJ15CnUvzTTwH+IdiBPZehSreySA94ONA4NisbiiNrUaD
X06Bc6EFHQUwAfk6jzyNvQv9nez6zvOM+4f/yGS+UkBmIIbf0qfxP/Av8kcGrK2v
cJgJe2Ra0/7VtO0cnFRisQc0EomQOaIXz/PApm4Uy414Gj0PQvtzBPkbh1f5Sriy
34kqOx6znnkcBeClmi7/kHcR/iJTRU2VTvOMmDG3kOdpvDGAVI3u/u8mWta/545A
w/cD8XjxcY5D1PE6h4uqXQGBrV1diAMCz26FGQGC9L7tCCeUDsDjQLO+Lau8xBWE
io/5ChpXHciycrQbwXX4dX5R3RaMMH6aiXamV3b2CZ9bNcQeFPbySBv2razpGspc
UlK0jbJlkgvgL3r24aL07WEOsWYqEnscX2wHaPuu0TuZr1NsayJHuqjjEXN0RFMR
s7U1CT6qXDFixJN8pUFfckIRwsTDnm+pLeQJlvcSon1jPkmG7E8AM/ktPplXB35z
5nz8s5bstdgjdLLompyV0GbApJGQBO/n2dRhJsZSq+AXG+iHO3VwVb1YPP+1VhsN
OftfUaHyi7k8E3aDZFZdh1YAQoSMiQyN0RkjBsvYDXK9y4LAF0DwmNeHtNNCkL9/
LFbCxEyv8FzNTK4yrlmB3Mg4Nzyk1OyH9kx4tlaOaQbD25xVjEdd9qGE+nD4CNlm
y+9B2NtbpE/vaNLWhglVPhSRLw0eVn8ZOTEIM1xHsFuuG2xctSRhPIJralz2RET8
lPc3qJ4bxP7kSjOFhbv7ZFouli/f5Vb86+6C/dIQB7amx6CaaOPVq0DmILeLXX1k
/OqciY4bg/D5s2e3qIcwzLtiYNknJBHv1E0M5KeLmac7dC9HmB9jzU1EpeuT45Hj
n461MIBsOSFPfcy5QojtY877B3p4UPoci9ctAR6QL6zs55+En5O6MuHahNVqq4dt
hIE3o7FNayfkvP5XwYxYFRKm0ZS86oBy9QBPgQcI4pk6u8fTjGZ5oTsY1P/Mpkok
r8c47st+U9WfcHj1a1R9vQ82ZDInK55wk6SUPWQ6boE57xwtS9ncl0sOMF5wnvZR
BVJWCCrfjIXsVV6xROJjldr3Lm6VCUnVrhfMMDgOszpcYnrl5UG3IDHiAuojmUvD
bQAGsk4Jo5p265oU+Fd2tuGiVsvfjgfAUBkrTUO3k5U1TopkVsidNkUvpJ/oniOP
QE2V3snosWBONOg5wVzJCS7UeY2ewlqEus6ei37Bo7EWU2m1qKTa8WLf28DijpXe
Xl6Qr6fUDh175gp6OGIQnv4QSgK9NCzbDO1fwxpMnORPmQtZy5l7gNMbdSadD+nC
xkvQOg85nXxs8SVMZmtkcqNIQJydDE+X/DZ18pN98gXxOwRRAbcU4iSK+BIwN4Dq
QOzaIG1sZ5VZAL1ocE5mOcbuQpQfbbO76yE+iXRVwPhwqGdSWklvLpqztyUDAwM/
aUAODxRROIxVgx6mmMM1Ywj7E4fWCgyXHjb/1FlkepOFWhmwD2iZKFX4EqVA3P3F
kiS86G7iKP6izkIoWRTJMElpwJ2ofrcODQ3pX/uMF+YphxJBfwF75rAFX3fdubZk
xyw2fJZNNNOhRab16uISlUct+C5Xqr8aOc6oymUN+46EPdG5r3OUyflKrA51WX55
AJ6R6ivmbBhdERQbQF6qTzvvT0LYN+I8rrlZx3J0rSV+0ysjXDYc5IcDs1RhKDVM
EgP+vqAEdsSBRWLeyIF46NDnNrhaz8UuWi1V7AmH3TOSzai2OlYyIJzByBZiWjwF
xeFl1NSYp+0AqEamHTGn011z5Du8+oHJNo17FPk7KZdv8pECSrXWw10NSkYa8H3+
TtSbyW21dzw2FaQJpSmHqTeIzg66Xe8Q8DC6gczxs7N5ra3Q9DoVbe5KovrBXMVf
byuiPWywzDnAlkTIHbCatHp4xpI1x1/1VYvvp3gomPtJWYPDt1+26Nk1iQCj6LlI
fi6ZkeX4G+SRBcHhj0WOOthJhlszcwphODD0neBn3jvP+PPld2KXr9CEJJJ3t2Da
RiX+eD0Im7gvQ5ySII4X1tQWTAVqlqS9cT8GCj33TypkFkIJA5z/neK9ylSGWbo3
PuUrXAFtbTcMrfXMRTOSsNf8cd8z/KpUQ5x/oqAeaC9Zpn5c9H5s3hkKoV3mU7W0
nEA+EsORn2GeZbBRkFwdy8LXkZqWbI9ruiV7QSzcBrFNTNAHq+Tcm5W5DBqI/il3
UmDmHFMqSQNHe76jjDL3O2bu4zUv6xx8jmmCyYE+c81WWU5gvsRv4Mei50s77zB2
lzuMJZxZ2cV1BeMMAagJRe7GwONwvYjkcfXVZkyE2NFcEine3p3l925dzwcSfaZE
R2Ygn0i+7Wtr/jnIQC9x2vj5z0+dHxezNq5qwuixhMoypYeUg9WfLOYhWij7fQCn
qnkjnpOiXDZZCeo4aIi0zS7ccLEz+Lxlr/D0AAqltuIcQX8sD/c2N+jM/9v/Ujao
3bNOPetCjxB5Gdj3txHrlMEJfxzCpNY3ggEe3sOuT+mwLdI5DFOY0GTpbRz5Z+09
Y0ITWs7JYtGNIZ4NORPXZxlKVKrP0DJH2Yio7wwTGoF6hV5Rf1clxg8zXOCAcuU7
9IgFOPdTpVqHei634mpjZ4H5aBtgOsz+WiNeJUkj/9lXQPjgfiin3u/1dbM6cNcj
txHldwI9/9+umYia0JWy3q3gZqWVlb1bommnyRltVOV+vUgbCo9U4cfksdJbvLGs
/yt80EqoftuT9a3E9fcAgvyfRcjNAqSzGqNAhj2Vmt8kZXWEjAbgy1Cq7BynC8EG
m4QM+1shslW+VKEGSRszt/Spns8Uz8EQz5Xps61D2yVfXFGOxokg+umh0+mIFyJx
pxzVFQeRgjglgiEqPj17BmEMxMAc9BFxUS10SC1FJVgIPC19czzasyo1fJI3+ooa
er71WLUnuYgUrizGOaDMr4u5OwNePJRQuIh6iMMK9YkH16BaSEy9nPxNSO/0y5T/
OZswYrZa66AWgM7qDAnTCeZz/Ts3LBuiLNM5//eYwhWJ2sD1JOVb0zN84/tsHgLd
7lt9ULz27an9DaXgEKlajHqyyapnAb3gVUAuvKElq4TBzHyodLwE2nHKQw30J2cm
IRCnAqd+pDHeBCYoZ4+tykR8SaiL2h9GxShmOefkJEmgjkI3juUgIe84MewRFQ9F
XbNM/sd60Yb1bZB9zdLzZkV5qIIJ1hzLIl1cMh6O53VNMaB6kXGQ/JIax1JmsqU2
1hss0HH99r3yNvhbJTYqsMndFqjXYPVoVL/X5/OJDV/gxZ47VsGrdQv4J+cFibDp
uAEX8ONQ40DbqI9div6lTS7NUqv4zfumlM5z5lr95uKYK31rwopc6LNUkRNObPVF
GU7KlxA3ggPG2kEAzx79qRGjGW8COzcDIaVnFa0ZAteXL+DT1wxqEQk0pyYJ4RXk
gPHNOGVgrCgoKzL28AYHwCJo2HzVk/Fdwfvi6zB6UMCdzoYRFUmRIFrJ2dblkzAw
Z5jyl0I8e5MG3M1IRrcJ0xJar2t1Dd7AqRLhUq7Ltj+GEHKeO0T8yesAWIWbjMp6
fxMjkMwr5r6tAyVZM9K7eH8EMOxMylHPWYos1PXyVX15elHCwW+OwkzERNLCUFvC
/Zjslt0Qd2gNWnkQ4EHhixaEewF3CrUfgiqvYtkDj93EKB4aHoRAJJuuPQzE3nQO
VgLjgoidOIKMDxn3auA5AA==
`protect END_PROTECTED
