`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBd3VF7gjgKZ7+d+1uTXEA5y/53LZvDgJSc7pi9/i8KpXh31I9hDVBZnZqhaI5kr
cUI4l126YhWLWe7mjlO3j8uGenK6IkD57u14p6Cz2MRLud2pCM8fhSRyg1/LrJJe
KfMoq8k9uXVJAh6clfVI4LaLJRC66Iaidym4sBdzz0tGrQBBwVwfjzVyIAtBJC46
AdffdhC7dgrlwnhvMfb0I3EGopefCWWFWWiRI2gKiWXm8weYzHAV4pOAcRTCpqCe
y7e7weC8mQ+6+qQNrZ3yhb3JT5UmXLD68p2g2cXUBtn4KHJHOHtJkBCt8jlkdxik
vZrpvaw799SY0j1p2sKjxF229zks7hNfjzPwjUNHjd3gbWnM3zJtxsIL8/YnOUZj
tW+CF7VuTrY7cEiqK/tdUTO0o2hrXD8qbh1R42hXz1QvHX9xaHvUcQT+3yOCU5kX
n1QhxN4hQIDhUpkT2S1qw1zh61qj1VOjdpUR0vbTPX29V6sCzwqEGoGC17drb3T3
RK3VR68qQZtFGFaAM5o1nc5V1xVUZYRYeBD7RhsU3qQCezukg4VxdqGA2oormD4O
KRQSUESSzbFBTV71m3JJ2nv3q70sIq9+sNN9/oxzI3JlBvjuC7HlllTbPpziHGAU
pPuN26kN+Kl1TNRe5K1lj/9M/lrU6eCj37dsmEpkDMXpDLvsZ89opEp+wJ4ZZ7Vb
s9xUoiw36/dgPdWg1Bvlmis4Jvbij//iMDy1BgbvWhINo7p+bvogqAhicNdEwpI3
sF0T2Un2BxIAB5Gb34ldCJjiX5FEkmagHxEJRkf5N5kzIXaFNtbldFMvivFW8+Oo
OACrgptKLVvxIEUEZTVbcWz/b+ifo1VCIByweY343AqixxZFyWr5bRzJ3Mn4lA7z
KD43OBoppWGPiBIuQ7H+q7ITF4Lp0Z0/Z6yO3qa8sj3QEaMzkqRtEHnqmB9E5D10
pyi/hZu5+cIFdpsTtr2+3Ayhc3ee0nvph2EI2mkuMR8wpqA6H3Z00DqU5Q4rs7bn
sRvHYg5BDZ/YZzwGwya5QViIv5LV+YxbrJEroIHjlSWBHKEEPoiznp0FC5iQ7oMT
3m8SG4q5OJ7WFwmNI+ZaOfWGuw0rGaRS7QShEJgRAy7oWH2gluO8Whbs5ActItVI
AN49yfcVJQdKeCWhENVm8gikYAmafMOiHDoqZMDB37+DIp//rwEWshYPg4lWhtCX
HPEFb732/WL5iSVuyUdS33SKmVmA/92S211VhMCbcpFoLaD6aTGVoCchWA4mzmD9
NVIK8s82bfDrLvJIW/xJRJfVNkHtts4F412O5sJsU9KuWj32mOzrb588cN9aW8cj
1F/p5py9Y0mhbHjzXV+4BqaYwZO2HLGgLXP32lbM23YppunCyof9GFfCSTQ8SWpY
u4sPDK5gAsoi2FYtQxClQviLvLbKFkp1c9PKSSMwO1YHhT/lp1Ja6CB/lxbFIcWD
oHKolfdELfkY4CHeelSyT8iUDOXY+mRDMt9MAjSmMCVAkU605g4avfIGUFTPV2FA
sAlwXlgzGrk6Pl5JJP6SuEmKHZb43PiOCJroEux3cF+PLVpsIG13XNtpxSxrjcYs
VFmiM/S4p1yvluGzsMp+UDlH8XG2tEtwLkJcd0QxshYwfiTXVUDRmynDvwm0Ecng
012DJO+zp+J0erYxsgEwOQcyDV3+ot5KmTeEZrA/vwlfh+ob0t7lGqZ61hwmoohD
QR0pv0Te1wdoS/mcwyWs7sq/BwSfG9nU8bTQbMaZwCzBwMw5YKSEMz6k18iAF0gs
5+HmDZy9sMoEDEGN/oGtKH3DW9VgQFxYwqdpf882IfmA/TaoE+Rm/3muKjeNmpYH
NEkNJcsn/IwX9fYp+c9t+BG85CzPTKySeUT6Yh0i/TaXNaObWlqT6S6MPWQLG/+r
hcF4g8q7r9QN4eGg7VUy92xUofClUUnfZ29qeuq1uBZ5SfEqxq5NW0HhTz+HY3DJ
`protect END_PROTECTED
