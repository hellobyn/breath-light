`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGnt6/UT98HWfx1Y430crdrO3WG/72KVd+aCEyeLY0UE5y5ivUL5492/RcqhShOm
dBvxhAJUvyeiXv0ibX/yQIvM81iuA5IAH2eGXptm7mfJGZ25Kw47cwQkJHEftKiZ
Vqp11uiwrz86h87qGgSoQHZJ9HuuEwUpRr2UtXG6cE7bWUpX5AzDj9qFA4I4Eu+u
M7nrsnzM69batoLV74EdJtusz2tV3CFjcFv9vhfN7ArpGYIU0RbTxulf1A6ZyY7b
Qu5TxRPFIXfz3IxLyvzrsAQ7gYN8k1a3+xJ9mRiDYDHoSzjuUUqHmFaH4e/QO1oJ
x4aHqh6cZ6NgUAA9nX3dfWCT7OUJ135bTrmPsHvZuFVjTTm9COoTlJYnbF+ZEaZt
DCD0ZnIJ6gymSIv43VYcW1zfEGdQWTbD6UdfMR3xiIVKg4R/daYUzXpqHoFHTI6N
KbIpm+7pMqR6+bjjoGSV/LGRYSko3+yiM/lK0Pctx/YRvCaL2JRRTASiDRhk+gws
8S77YbLmVCEB2lTvoMR3I5cdYlLu6JzytN8kWSZWmUqH57Bp29aEtqxfZlf4MyHa
cUMSg3N7wDXffvqN5YvnclBLBTOdh7+GiXWpsSAuov2b6tE7jO4AL9ZoXlTimU31
3kwVw5hfzqXpmx4J0x+AjB2Y3I1JNjCYxhHPYjy37n39qvhNTZagO2kW+4VVKM5D
t7NrbP79GXsr+9ggiRqKfCK0MPfEJCdX2bnoZ3qrWEupLaeiIdviBLoObUz4SE5/
dagw9fYpcbzT248Cby3OuQ6j7FiDoDXBpXCtwVyyi+sGtSzyMHnFcoyabG036WC8
0GjTSH21Iqnssso0s4kDVeR8MUP5TzblvkXX4w7nk6hA20rLyKQflBayUkSzphaE
84tUPCN7NTPRX/LXcCbyfzt4D98MEqkHQI1jVv4Ow52uEXYECHfbBfa+GI281ews
fOPdiTHtzKro5l7uli004CuYrxwNvCC5ZxeJxxK/5O3i76ezM8yw5EuBFb9Zvxt+
UaxPfw/iCWmRufl0pGht3teIn9lxNGmhewMylqQJ8hQOW7ZSTMkaB8fAwXO1jZXH
uAnms7dLOdthmtF7T65hsTRc+KrKtqQYJsfxQ4ldaQdfS/zu6Imm3AEG82Tq5J17
LS7YmH/AE1BnkUofYFWtx+TYv9DdNUZx0ThLKV95zuuRfIg/s54Ws0ErDKwoUyzz
Y8Jdro2e89+64AoVhGxZ768qn+I/+P4HZq/+ZCboAMK+c8Lrfwj6sj0JH8z/GetS
NL4f+AhPMq9Gz0q1kvTtc9q8/rNwktyCNu9Ui4d9Gqo/5Bu4Gd6V1mduop+PV5ep
NPSBPjUIJfjSpyP2TLGh90meehlnrVteLuoWmgTdCElAIQvHO+by/ZhFs0Esgm4n
1AQyUm3ijcN6Z9Bn6V8oKdXV6n7ipdrHafh/XFJch7SpzotMnqzEClq9N+g1KXtU
s+PgC6Szm6UQCCmN+69GV+14fyZ9E+l7IbRY/AW9JuyY6jbifdaVloedsUWJLgzK
i+cY2MoGtlNCJm/wsX6FNeEsa4rvnVp0dexh3naEgdJBL4CYMr7TtjOn1ldfrqTL
vE62TZQT6Fl8+KThRWaa8r8KpaHWb514aR7YKwuqG39yVgU9IpoHGrS1f/XM1v0s
BEedWWGq2wRwgtBz05XlCa1sItqWg6CKWgsQJdmLQvzZcavFBwYx/ob9RmHN44XL
JStUxBLZWd9GPyzQvmr31U5WuN37rfVh7D1B7S7V1jEdgUadtrPutSW2L343yu+s
2W2SXU6NnXJNiqlD7E8JAQ7tQ/Qi7LIWjygd928dDtzh2XW2UHYZvTElCzZbLoBU
wZ4gmTxyMhuT8pTQ3XNC00J+mCT8rLHEUqiIjTopf7jqwcFc8l/GLmj6XmX4JEIT
FuyFFVKt925xPG5nyaJaChDOJkvNmvDG4QW1p6gUIu2MQPtqo06yUnahjZAfMOla
ptLC3ceVbIBX9BSFj7LSuwEDz6zGPVve7mzdq3+TD3jTjGxhCyh+DVgfcFNszFsY
7CKWW0hKN4QSkdagN7Wz6rUi8AMEsywDOFaw9SyrpZkz3H7YCyDxNZc2GB5Zb0ji
/MC6VwSECs3A0KJ4rJwtJBmvDuSy2ZIQLqUzEQ7vjMwxYa6+1FkRv6IXirFNQePZ
CGMYGi/YPQhOCVmpByoDeUHukMQcewe1i8kPgCpjOeA2clwC/7EdbWYotfwAW0j0
5/tGoaBCkX49pw8n4I7ptKnscQoNxQ2AqR7/Mgm5ZLtTH8/0h/J/oMHumaHXQ5ru
Ria3VbztIEwdNo/7H2BkthJe6Wvfqy9dQG1IvCLY1LoRonyR7IHdULzK5SU93iXm
HoDGJl1gGXGlj7yuKf0ttAExKPYD1Jj1gk/atnYsZzS5KNkMkbUore4+4bSgh9YA
`protect END_PROTECTED
