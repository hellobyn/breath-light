`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+U3+Gz5rF2hKdCU1EUyhqhM4TtWPMTyCN44Hz2y9FzEK5rBgBrKlNli7ChMZM+2
sRI3HYrDMId6RPJphsCi3+Hdlvf6QhDUe2KFx7P+v8cX8IbhjruNzxCmLuA83QNI
n35qkabIXWENjGsvIbvcAY9zK35ZgmKnNgQIMZ5EVik9lLWlCjGW6EHoEHNuzhvA
k79VfPreTZbF2huHF42XdJlucSAoWCEISPDHq2tQ9CXvMuMfB9GRHrP5fxW4jiWU
1W40Ic2qH55CONVQjKCSKJ14AV3gD3uF3CSNl3f0jJya79L2GzVK8e09rvzLyIlP
yC+sE6p9zirBFmye4TcQTFd57Fl6U+toBmWI5mszT/1yLeREgWsUdI6SV834J98P
YP8mGrw0wyEB29vTReHuyC+YvDQsf8mFkpSpoVPmr35+9H8VLdXyYQNnowa9MGnm
bAjuKV0aquJqREv6BELKvTSzhWqd8A4jJmAA8FYFvslScEky1lc7YAou8ymm9GOo
MX2saA/EQ5NdtU9fxrWMfIB0sVAqNgR5DVwyXAPxp4Z/YVdAeI9KMWv4jj6/76P+
BrO+lDX0ztG0GIQcsU8ggryc2j0Aomundufxvsa7KR/i5hg1qfzPzt1CrhnVDbNn
kY4TATY15cCfQ+89VaUnbs4txTALGkWwQfa/mjE/7NvaDabujSQzNuAUjPvxGH3p
TCo4xCeSSizwulICa6q/Wrd+gkuvZK5dVr2bHU/Bpc3IefgR1LYd4bFTxQkPu726
i9++ptAeMsTWnbcIrl7ASFes6fmK6LmDI+jbDa5GNv/evasBQgJTDwacJyXs+PbX
SoQTB/C0NXNjqsxbNDl/DLE4sIUsLuT3aPK9Pdw/fG67eynAPZHuxd7YEqn8/O7F
4gi+kirsZ2sPW9wnvXOmXbKUNlW88bsdK5mP0yG93A98n5SXViLyGHeQ1om/qUKA
d+YdxyMT5yRgGfi8cZXYCf1IEnrbhOvJtV78wGsyyTQHzivuxHJ175DKlLGSGiQX
2A1ppHJ6TkLrm06K9hESYI2XFEQ8uxJQzQiTjLm06lNd7iG5sH3mTZc4Ih23f06V
fU32wIgZxWN+utuHbbSuinOxMbK6jnmFWH1mik4FzTFODRlaQ0tRxEmwIu1YIqIo
30cXVJO34dDFwSUjhWWiRvWSth8Qy2M1nHWNQTh20vHVzjvFjELhqqb24qKJJm/x
7a0DtudyKnkGLE/RpvsUSOb0TBwnBdoZgHtPLMFPzKmIPOrukjpNhdyjEf6sC7ny
durM0GNduanPXyugcjf8wtrI9XFPklfIGgFVM+BfSnIIQ4ghTH7LMdTa4uzdcnci
sdZFEjs1vOfDRMFF4/LIckxxFkPIIfRP1w/9vsWlX4wlubFPyX+HalrSGmjDnooW
Z/qOzOC1DnbC8X6GW7/Iiif7t7yRcENe5Y3iYjNs4GwQBRJ2Khw/RnH2f8J+H2F7
Xkb1j4L2VX9cpyQGObkMYOQpLA2jpjdkxm3j7CAA9TryfoZL3uYXOiLKeMp9kvGJ
+RUbjn5pBAGXmTTjkJKXzceIQFzzKbtK7d1rzrxwIkcOWBSxS6azeOST3ZUN2HdO
qzXAMOT+tQvcRCVvak+rjp0vlcAhAjyPFIurSSGP/omDq0/ZSy6bKVnhqTG5Qu7L
EasfZYXgwC2bKfn84kN1/R6hWlvEaSp6gHcInw60QR8=
`protect END_PROTECTED
