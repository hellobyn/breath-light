`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jG+33SCZBdlv4aE9t7GyzMJEReUT9001yKJKQdqRzPU+JXP218Wn6uEENIaL1aU9
3Q330bQsVMZxOsg9MI5iqkpl0o9ode0NBBThQ7+d+bV1u8laQ81JLof9OxgsXHIa
N4dZGf9OeFZ4f6GyU+kNtLmdNz9RaXFGAyTouatecVB6ExlDA4LbJEjkwJ4JKuER
hAK4MMDMcQr9hWIevTFIkYwkH91RUIqMAMBgdKo/EQDSUoGBgDfqjaJcCZdufOhR
/NNnqzHGGisppnahzplFOeYi5IXKEbKHL1PsgjfVARwRWk5NE9TIA162I8EXH4QB
0gF91yyLC99z+3hU7pk/mSzrKRCZmbA4TnKxzdhTfG3n07vgEMm/9nG0ySoExpci
PfBNH6z3JGqd91YJcBP+txy+Sc2blbRaRsiuVN+EY5zNPcxS3VYyRGGTq303iS07
9Fgjgvztytb2Dvj2uL6rvoUSteovbrqDibZDthQptkPlZ0O3GKejbEdXySHCepeT
gRS2Pf5kmMcArMwGip6EoR7klFVCc9LIBNfdRB17xo4reWbrhVrciuJVHEFCARKK
/xvCAkTvB53V82KWOSzdaGCUxQUHLvf93cth88S1P2NChmhF69BzxV+CBDZZJKee
esLIQOTqkILUrnoGACCwu6cMzPrCU4+vzr4xfUvfN8rT1H0eD26OhoQtyzIIIxI4
K71CfD51oBvHE8Arv6Zj7rzhwHalO2Ch2YZRKlf9HFi/AvAP9OD2zTtbBrXQWIeO
T5pwPjNgKxqW2ynieIfpgcdlOejs6LxE+F8mD6hBFytg5f6jAGsckVHlRlt4szeJ
F7u7IiCdlOlNyoRjfgZH3sVKL6EM82wqZ2yMwzrenacO+nA5+GXBeTN6MJ+n8pci
8NSCeHZb2YOZ11emMbt1xmbFuRGygy6BeFvFHQ2/fw5jzPePEC3OkXIeV+QKGVM6
zlXAKeLNFoJT8MlQlywvi2xMLP8P5jlWEu20AbqkrdCT/lhSA5XU+V9wFoI9BYFk
BReN/kon4PkWWSVe3E9mF7bJyWgM7Him4zrni45QE35qKM9mbsXR5w2WbxI6ecDZ
Y/v/wt09LQdITKdaIEPaPleb28ydsiOY6env1drNXfeBjOXE/uEaYKFGSyMUiGLo
w4QRS2HkZ+w+G5O5zNmRrpF+/Evt1w5b/7LTeEa+VlqVJOzH68ewUndHs3GHKvSZ
vnaiV7Ll4xp/ySONOD8oO+F33SEX7MV2/FYPso8ns8NnIFArfqVXbu+V/qJtevSt
nPoj+1JK4qN25s6sYXWr8ftQ96gbGMbhDgn+UD0J3/+W3rKREG7tzVUZEf4arhdI
aapVCQDS8t6NJW/gJDtMRXnS59ZEzLuPwbUfHevM0FBRzX2J6LY+jkcqMr0uU4ru
`protect END_PROTECTED
