`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fwrix6Gm5/VaEJZ0y6OFuqjq1iJ3tZ+2w3siKDOFwxnzQqAtMDcuV7l/0ZqipyMV
cDQ9O1r469aZrOWnYO1GKNULYtjc0FPxmKfxq/QY2f2HTIF/3l4BR6stGK0wDc/b
YmxqJeBNw/w2KlCesw9IUOfqDhpnXaPgEsudaD3i8Ch6BAmAu7qe560h8VCygyS0
i/aUnUzHSjh7PohYngq/nZ3EON6znLYS/RXZkVv87jCkZzoa+8hIRjsBtnFfpxso
6KAgBPd21Fp40yzftvUVa3Y3C0VAVJlsm4Mj9TeDFZCewLC4tx9FvgDEUfM5Pucc
P4ofCZ9+8SZk45oKGiBFtlTCVB6954K5X9H6MXVeaISl83EstFqanC+AFvsYoNkl
gFrpuqa8g2jJksPrSkxHQFu4S31espZmuZx3fQ5GzyiYwdV1QOlJyPCJhmkEVK82
Cm9fFZ54qWDgQGGnAvNsPYDnc77QL/eyUFHt8mSA/IfROArun/xQkA3+qOJM8bG0
QR73bYfeTIbArzMxWaChMv8SGhX558t2laj0s/MqJgUaq3lTrivHwMu//5plodnY
cF5ljZZMyogngVaZXrP7VkVVEMT3vOlBdSWPMOGtutWmud4Pmld0eze/rE+xOAZ7
wD643A2DeA+zZUpsU6D5bDslaeYkyIUoSWs6bpM8n7cQvoUXHU6RXi6TB0/fMcYv
Gn6NAFTMXhpT+AHjWoi93FShR9Bvro1KEdfP+4zeh6ojCnPg4DGtRjPAmqbTNlQ4
qZy3vIG+yVP5a+1v+Xvy5SkcJglyTGjIUbYvYo8JqC+hZAsTk43H1Vd5JAImUK0p
CAsRhklhbqnZ86wQ+KfitC2zU0i/2RpfsaY7P6WVxhuS7IdJwwpXqXk8XfSxBRHf
ArIUQDbUfsi4A+oMHhW4U786xVkI8rEeyK6QwbhMCoLrBvsnMjbErtnH3MPE7aYc
YTln177GzbfnPTWn2kJ1QhDB73mRGT0z+NdUjwTqOUXBIC3HSdq7wztnlien983y
2UsFBaB6HxOA/Nw5wTEHd6pTZQSL23H9ZTHwrl0ehN23dOZueBtoRkc1K93Nnprr
b8JtIHI9GxtdabTxzpkg1CAmM+/IozQtGYUqPs5ZGv+YTha25kawdJek8hznI4FL
8ydyYk8+9469EZxOh8J7T23YDOERk9Fa1TGz6T8gTlLVY5xeMlpN+Qk/okI2hnVS
G6YJxrv44KXaDWZ7PMDFiEGKnvUoA9ZcZS8zHQ0OSyIyjaZb+HPk2pEMYkxRUwkx
+wc28eBlx7h/1ZrH7wp0ElNtIq8eXRKQNxwYuNgTmQY=
`protect END_PROTECTED
