`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jovdfJidIsKnKqCOXSTMpjWPzXhqahqUF4yBRdT3ki9TiFC+Xh945zmTMKZuQG0v
4/6/afijoDZWULr7NklcGbucAYV+1ZHi1Dj4ciqu8kv4/AhmSk3DbTJUpPlCSRsh
UXuGK/Mg0xaJdwx74nlR5zb1/64wxeQxKImMg3VEoZxDb/uEhbH2FGz7aBhaPDCT
kL1PGrGCHby8ZNz1cCfncdHAOzrG/TI/hXop4527a673LGq38bhOBmOyfxxZmxVD
nWOt7rFRqZB2R7fXilwlpIrzZ6WuEJcM8rJ+NbqRHuwiCVnH7qJgdfeIOQWS5Dwb
7D/6Y19qgmDjuJPydX6pebt90UoF+lt9fKXUg65EvxzEINk+jk5wL0C36Abw/JGk
03n1eLfiJOvq1oHGu0/EumCKZgCC6kdnlaF8LwBPIDpMLb7vrUJcqKu0Zgno1sCS
tD14/DR0UC5AFWEWEKdX/RSkaY3+BGTJxyPpABiWr3Df/oaJtbKhb4zKMm7bdqtD
pF5M6846iZEXmvVJI6fQxc/I1+XhqsFDrj/riufhzePJnnOQ1qlOQ0GFqi4zduyQ
P1jgfuLHv2ZoJ3HcXCIXvINX3jSuBKYxaf1UtpRyPpVRMibi2mziQiKkOPMxic01
iwAd1rlMGP+LzGq1/tWUmzkPnw0MmF/YuFPIN6C2p7VIeMMiZ+Wsnpf+NC6FEqUs
8/tMz0NJSJn1qmNo5HmmU5OLeIvoYh0L2FMJSTKckM236u8CsVyyrP9TL4vWzEPT
EZD4nuZAeI76xZm9kyIQQ6WGVIB+UDhR6CauCojxDlVAawcSBhWbeAxZryGkHQmi
SLnadgZbbTRroRoQshHcyffMB6CLLUyHE+SdwdsnCsxwUXm3xQ+K6vVBgIO+s7PV
laGDChdWasAY78AskfA4/OWU9Hh8IxFEUh1bSOLxBsR+EySr/11VrTxZ1GKHyMKM
si3sVQvYionXxU/y+JpRbh/qnDzEyT9PVwkzNwRdDWSiYqE/zQdqKnKFZwebbdfN
lbXtdoS2PFrreSlNePcddm2+Nu/fa2qlkuDOl2FOie9sw/qkjgINnbq2ulfZ+g3D
flFBeXDgnx+7ueLsgTNwgTtg+RKLC/at1YpRecbRcO2jvYfGgaZ2RJY19lm+6uzp
V/iCopkI8/YlfGPPB1amb+Zw5PCT279SxtwEYdDkBlOuAPohDmq6un4Hz2o+zhmF
9iKLDZBTwzNLYz/9aADVIBwCQ84wX/VodbJQGEN4Vnhfua+fuNbTjRjLcFiEQe1C
ihA4vZGO8olajIw4xQ3sA1hixTBjshYyNmJpaCKkSM3oSG9sf239x4GzhnGX8aWa
CRbRM0mjnk0ghIMRbqOYNExKg3vtQIvjxqEZ38gwgTbEM1K5rtGeAHL21wgUBeAp
yoysaxEIrPxoCc/g3O7M5DqyGQ5m7FBW1MTgJ7mmB87hvGVVs25VAGq56IdzCBmJ
`protect END_PROTECTED
