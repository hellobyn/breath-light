`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dTQjadyQccRQ0mwJM+7FO26De4YbkAmNiPXmVw+WrT49W1tU8NwyQPbxZRpE3DAU
f2PR9MvOTp//5cJIGI8yKCVLTJPEi3oRZX3vqtQPck4qbb0YjE/An16ND38ryhcH
rnGwj2YS7ezzsOEaGtsyscgJUoL9w97Ka8dl35tkPKy1ClZu2gkPStJ7F5FeK8ce
PDJ3Sed6thY7ua/Py77Dy/9KPs6V7YgGUbZ43fyk7qjqKwIJnYDdc4wEXwtjeZXs
yyrwth/ASx8YLv85ECd+AJVoHWDDtE0BdtXA6tuqIJRXPlL70Q5S1MyZzR6SEuV7
L6Vmtdc3KodFTqdAUXco0KvUZTXyaptG8BYR9vRF8n1IQizQ+QgagJPJPBhlfcH9
v8k1Yip6hPcEUYqdVTnK1o4q0bi4Zi3j07O1Aw4oOglkwop0y7X+Y/+5uXlgzQtW
U9uNidhacmegALwQmxUcPpVWgue8xJqwr3cxOeSLayxRP6rNNlu6VnpR0A7fWnyb
VKmN8mNja8rsBoEejrgXIK77dpAOW5Dy3kNyJXefwCUTTpefMbJsrocUgpYOYUcw
vHtDFQ9pjyZU2Qn+SZrdCg==
`protect END_PROTECTED
