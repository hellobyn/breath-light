`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
McxeYOZDSJN4usf0OhfHcuPLtxTjXfvkIsiCY21KFecBxIpAn+yUZOmBPg9rxtkv
1CoH+sDT39rKD9Y2aEz09T01tIYA0tUTE8wdQMmVEjDH+OvI1ajStNvWhpcQtktm
NmbKPQS4OnKqDrmhDiwaweU4pOCtPk/gGRwuXAOsFMwSNlWI8UULHzW0po17+03O
AXlK3HJ9RP52rnTIvHX5le0mDKDyLoaQtVIcRHxn5FEwIiB4aRIgWZITtnQq4dZw
DxOZ8rJPQMyOMbfC6Z0a9ZUXrLsprvsXar4JBxFxadCSEcn4ljZmmWUsjQDP0XLs
sQHeLDxTrUN/yliH1/XFMMPziSmCwivvItWMJtvtTrdJDIszP4Yka9Ovh8NKxmpE
wDGevmRWfdioQaOeVX5hzOf0nFAic8+BISqHY5YfJXhoxZ8udP+ZAf9qw3/QeJ0Z
q31okjrPFIYoCASrPk3qETfPqNPtesf5o3wa3kZC/9sWNB8q3CGBRdTOTOtwoJgc
FbNlK3FXmhveQuXg429AYAs2VjD3EN3JiXEp8JULjBa24xDF5jvh4i5hEjPlG9+Q
Pvby55BsHQp6PUlULnFljfl0n6W8cZrVF7QDYEYk2+KhCJSn++gvQmNbBDViNQHv
AaadAmmZbgsmm68LEtLm2q4kDNyLOiHNOcbLf7W/B29vP39odnX3zkJu4TMePf9J
7YgdNZQd6d45kdSGn4EmfqMbeiOqSbpbr3QvLi4fUYQix+9cf6doGuU1DJijZLT/
EXWqwN3FVXZDljsjbLRj7kTrtNsqgOQNHP4StfJ/LT0xsJY9sQrJrtnYYS/HSRt8
9crRuphRH0/A9FKdBT4aLrZ9+rzYMzufakSJDjgGQqmCdPpThvqveAK9W6iewONI
n2+geq8uC25a0NcXlqOjONn8EAOyVfgj1A8R4AhKRCJgoCaQEQ1nPhzBsHrpp+QG
ikAtyvnpUsvvBSp99E2xFhatFJdoqcKhAcdMzX2RG7UIvAnvz1Ch3sDNcBPkjgtW
yX91ZgO9gc3I+qtARbJERpR3Ht0r7Yz64wDGUqzE45H7dfAB7Hvn6Ukxw6oRODYV
SEF8eQ612JPJ4MHuplefQ49i7D7Vy5JZF7duobSgXHuYT9eKDparF3x7XgNOvEn2
wqjHZVSRNXRItqcbuZvAePDePW515JYDym8DtXO06LrhTkUipPpUr9dhTkrbMUtp
GADlPKr84FPzzvDoDRF8N49CDlMPkeFqqf2HPhxIC4laQrP0AQNthIx55dLBEMqe
UrapDSN86vn1gaYIM0nOd+nPfFoRErRwyCxh3xQjKsho2g4EfchroTZ7HlAgLz4P
Ay1y+pwoLMWegSjGMKXPSK2o0tYjzXqoODaFuPIEP3FyTII4kms+xSIJ23ckYw6Z
AlJZpb9Wz+NqPVj6Fs+riJtBq4BLgGIWHnLX1PBlqY/KtDTxqtxYST9EOrJx+zMn
HQnvcXQrh1IicarQ+wUa2I0W+OT+a6j08W+v+OkstVZy43EI8BLLztHZ/m5v5bHW
42Wl3SqMy4z1R9/m043dprFWBN9WdTFpprKnPjnyC9RbiJ4t4Xh37PU3OdThKVgS
IYWLaCHnLT9LAfQRYLA/217vxIA3//2iC+Nh8riFRJik9RM9fqSP02Z6/l2rpNSj
opsrTKOg8Q5irILbWvouzjSni3RTraCzBh1nm9cYj/qTzbFxjG7bo1jQ12Iu/ZR1
k29dEk9kunag8cCyv4bM59jAkCyuvAY2dnzmVMsCq1Rf55B6CURIB/tmwfvT+4g2
l3N/Jn3D8JUs6yq0QfFkkb9u/1G7fB4T70Q5ZTrLgB6WxgaMQGO/eDNjOmlU+xV3
O6WOGMgFcKecaNSaNaH84OcqCIhKfG0JNKbF6JwhrW1iwQnn465fjGLkNl5F2Coq
ufZSZAsarKOWUbYwWppO109nUgHuKXFRiVSBl+TU7iyth5/HEsd1xxEP3hnT3wmj
UPXzssuQgT5XLY5oeKiRukimCIG45tk8g5k1bWJBKuaJlcB3BQwJ9/fbFX+xCD9b
L9UV3TNqMsqXPg3SrC1XJqhSVrYesm2l/2koSEPwXhug7JEIFY1cjgfy2yev42ee
UH47rPrhu++aBfQkN6TU9lvhrvw3REcf5ktict2XIs647lUFuuK1Nrwn0aRVu0sm
43Ea4zgGnq4wN3s10TUAFORn4vBqqqvBDB9wbS14RH7mycNpgHAYGxkWEXJKHXqs
wJYoUyHhsAMnqmX4JyOGwdwNaLp+patjKLm0v3NwM8u7DIrmykIwO7EROIgQEoT9
AeJzzNqJaaeUKh5atPKCbQS3N10PfnAbIYqUwr0Pu7ydM4hkIKQcsLShho9Ojsvr
/3GeUA9Bco8FozoRBH1Aijk5MIk7lf5BHeaNIvAzWkOQGzSBuViSsCObLd8g6GYF
6YeprUJfbuugKq/8lz4kDJG2JQ/E4WZyIUn6XQ+b+Wcmj3Nly41HJV+HdMMaAc2g
6NeBP0OZGeo8vRnO1u0nb1J6j2sEBFvV/KU2phcX+4UAAt22a2EaesKRn7NU8ZFz
F94EybvR5t/ZxsHMIM7YrR2jhhYa0StFrsf4vQ0f3V367jQTEG+AIfEPMGyW/IH6
7uzh51iefEn4qHK8IGrjv731u6mWLWJcf7EE64XDCHqBt5M+tqWC4fQLz5S3VldH
Y4aa0c2PAy6o24yETK6kvABKJLL6LbkntBqp+PwOBYmlgogdtrCqJ2kYicbfm4SI
GpLRTePYn72Z1K6ZGC8Y88y6Kvl0+DmDIx96ysruAFxx/qqcMgSugW2KZq38bC9m
Fd8lijuCRMxZyZ8vtbG2lmyNmgad5yqdCWMizpT+gczmGUglrxOgINUgyrKcwZbh
7hy+lX4franxf6X9M22GQijkw3MH8SAmb2Akgk9fNu+pyk91kPHSgSJEhVYlwPVt
ehIQ8bGuhpwBEiHQ9lzST/CLoIQwscbynymUwKofNVUatiRQy9Sy2huoLZOV49al
NG/KlED9LAp84tpqCaVTg5aFvyMjQFeQ0lOAy3nqfyPUvFl/XfGOIp0Akq2C3bow
KeuAhplSyqGE9nLxYnvLU3fpyAlYwpNY2K+5sJQ6G2Gs4AszhlAvT0Rq4J0fafBg
MtCh+KcW/Q5jomyT/vuCliQHz3BSkpRL24+/EivEH+qSxg/rNUXTR79eCzX3jiBk
PRE8xCGyEhQbsR12B6npkp1RcVuhBxJOS9RyQuum9Ih3iw7M43mWCfUKXLvFAKX9
cLKw4NJj5gkjJZl0qAd4+4tBFmmhkMj8CykvOeT4jtikTiuVNTMn3gYwfqLDa9rt
teSGI60plvLZR46teCqaiFGNZ/q4Yo0rvE0+bKmoC67MnGrbnzenjUNzeyJ9pSZN
2egVpzzuY200tcOutvdWZuDkxEKSEkzvEN27htsvS7aUrlSSAqAshGNFOEQPHL+r
hCJj1mHy1iOao+B3Un70cyko5yfDRrGp+4ty+//tWNujgUb6GWtHxPBm8/7iFuIv
y21QqSbtm1s5ieyB7L4RXDUn+zzAbMefaX4cydnAQi09zOdBGYKdozOAtbuUv9a4
dWAzaWyJlywjfcEmSs6csdndNZOt3Lp53g1muiKYdqQVV/xVNZqEeBohwvCU9JhL
i4kfIKrHz9uQm9zsaFwTbumhqUvbn/HsG2xqC9HQZKDBBlUGw7BBv35O7IIoxho7
a6FdC6oABSyyAnxuvp6Z+1k3jZRBJmD5tnG1BuE94cqp8TDqAYMLFphqed+k+lK8
U/MRngN3lzNJbbQi3Tq8oDl4auYlE+t6qfQFWUuraORV2vJeCK55l3aCzBbAUTgb
xgRehRyGIhdqPEbCpvTxmoNk0DSCZaQ5FhfdXj770CMIMlypaPym+OCCoQSA0VI2
i+dbKdH88rHJ/s2SmFfeTLQ6RL2YCO2eLvWgKdjpUk1lXZHRXMu/bk5bjfV5fQnW
bN6LP9H/XvtdzTt7N2Cla9KeyV5JsZa15enJ598kt1SsNTQBXSY55LNPklPDyouB
e3Ki8nPxoQODM/nqVFB8ZmZeYqbYogcwpnhrZab/C5VU3MF9MjDZfI/XV/KDR2cX
Mz4hxr7aVVnzDgkfW87meaIitNpWWEDKLbyBMY0xcgLM4RK7BUlL0enEUDx2ICAW
NYWr9lT2bB5OIn2S9yFkkMs5kGkQT2XosadFKDHgd1ksSIBJaRTInM7W10NCUv8i
JNxCOlx+pjhe6GiUf8evUf/c46TdqwL8KjD9bnf4wQB/LBVvY3BDWUB6uxEZypPL
qNGvfqgpXYoFRdAfkfCX9M6jtFfpSlkg+w/Mr0WLDCpLOw0DmsuwugQpqWT3t8vv
yu0czFA0k1a24QaHocP/16uebEGDEMB6eIkCydKhMHTcIxKe1yto/Gpcjc6VCWbz
RCninXbxpDRqNrHQYY2xyZ/yH2dA0VV0YWHvhmrQdjlBMZBFMAjiIdHerYOiLzMC
WNqbzslcEB0YJZTGPBzCgVZhqBj/aAT0RH+7JWZ+LtaY7bJCta78ZpTwahqvpwrZ
eQW4tdu7Zn1LW2Es+s+PrEIxHl5w+mSrq1jwfx+B9e5WPI1caQO9HsAnY6CGCgR+
xitbSacr3Y+Rs26Lg8PkAUiQ2tqUGXzoE5YeNTx2RGwlmT0coaxQFrmg1hRaDOEA
eXYHAp5UL4HgYRFbbpoB3IdWh8Z4fcirYUfdjgnn5bsjY+ZkXZh39Wjd2rHw4BY+
1OACFSg4DaKtdiueMV2s5G/3NNHD7bRqlCaVxdHcH4HcQoATtiz9BxesxnxA9b+a
0eGbdbE7w7PraevJ+gMTrNLsQqaILdsfjltGsRyMPiMk05URHZYZYRUeyGoJeCKX
LwcBNtmTjori5dae9R8fn5G4WA0McPgOxgI72T00NVMtXw9Gd/z7bdfgO9L1K+K4
OT4p0ZNltoUXat76EbPn6IpmaP1Rft962VwvkTaKbrLhRFUitCdxBcmO3u2x9Ohl
uplB9JU3lpbRTDENBqNV/BhRjKdsZ9wTVyDkAbrDbeUcCO9f607NTtz0hT5xZhIR
mH0LsIw2PSCG18rCKaWHUq+i0oKPAUm6usAX3/gfCuKzjFgIt2qGNH/kT0KvpfQx
I5poKrdQH8DYWR7MBJ3bAZZAtZhsGrH204Xjqhb7YJm1Zr5dsZ6K1CpBXM8caAmT
pbVqgnC06VQZsoRWLxff3KAJ9r4ST6s+3dAVfitXYDvd7x/dzqKHWkqxbJrw3eOf
Muu9KKxpDt4y6KJHg00a2xzyiBtcRluWWQshuCNKOeCe/tNfiYt0Ixbj6VrGnrqT
XoA8djIMETThQIAXxCzb+9vC+pqtDG0xQlEPGMAWO/6M3PUBzq3boYKghGWAX29U
caKHqE437TP03GJsJjFot2JMDcbY+O79zWKfTdMLIvcHUtlaqdHhiWCESZrl2cyE
woVzklC6tD0sbVByEhwBEbLO2e0UxJ8mZZTACBIRuc0DHU4X5qMqbj6gpN8Iq+Z2
uHfET7Mf9TjIBTk3j5EiRFz4oAATPFsjqMcZK7QunhATltOzCVWcKZrlzhMbrjwQ
bSmSnY/pY56gGyXgIqT8jVBadE4xV72MpVJqo8E+NsQ92SsoJQIUCIt+q5gf0wLp
ce4ipQii1JQt8LEt94zeDhX8CG3dTRTdbq63agQuSbCpWjHlILPTTrtr/LeZenUg
YFoqakcOrcs0i/oLvxMlx2E4L1jodBhO9YhNXR/wJVAqFMnQQdrAZrkVGNGZyrrr
rENCMa3Mu92t8ymtEJ0fSm7fnCViTXJ1eWf9W7HPopRVzSYBFuLkw13OqECPS9PP
meBG22SfiBXkpIwXvlwNsfQwi1sWY+oPaljoYMosusYCVRyQiSYoUrYeTr0HWtGs
gZn1IqF5cVbzsZb7bz2qn+bpgEPJV2HiWHUmsW6u9LgAytt+24OpaeerMP4qrtwN
dmGT/RTLDQO1ULc9Hw5Lm0iBLWC4o1xOKKhNsN76wMIo2DbBditoDVW96uXz42BT
Jdz3jeEe9+DevfRN/jPKzCM1oi0Gqy+3ld7/CBWFarGCT1aPY9Vv1kmmcOZinoNJ
ir/Ru1KjQ6IVQv0UGdCljOvCGFv3GkT+N/U8op+77ge04y/NEyYv+5xTh2HFltuZ
O9FWZ5y59+EVM+zYy5EjJruxYQAVRUxT8Hgso3EfC4Wf2bpeQp2rUTEyZcCPi+Me
570ioPzEfr7wpPSs0sSp1eaX+seOyGnJM9qNiw32U+dv8RaktjzonZTKTXvb3sFa
0lLnfECYCgS9greB4bY1OhX51WYllBdZ8yFgaalBl+Wf3cDM07BAy6HeyCLlPJmP
QXSRTz6rEHfjtS2dESKJY6GwE3iJFyHLgx5gPLsT9d5iP5QDgF7Ar7XqpIJmYaSN
eX4u5HehK2wGjEQIFD+lt5Jzpnz3pY5Y2mSeLRRIVz0bSQ0z4cSv8GO+koYCt+Bc
nb+4uWVAHyp1dRZG9UJavg==
`protect END_PROTECTED
