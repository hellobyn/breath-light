`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6CyHO/3xRb/iEPY6QogjvcK4R2/xDZ2Dv5AMG2iam2U09BsZe4ncBJltaYV0YTC3
jf39Zx8uCOZ5s91ysrIp+2tM/KyC5qIB/m4PZhrSpUHKj/rKbWmO3+FZF/8Bgbnv
by1EFg5DPcgfnSpxIXMFEBFUWMJcfRZeOYvem2eC/HOfU1B+zEYFtqw2NX2wdDLI
OtdZvZ1FGR2NCukzp17xZmJP9hBW0LGwjQD+jJ9AKWTs3eAVlfxCWGiepjXELemQ
4Bp8q0e4txKpmc9+TmnGwVPimt7xEDVGc/iQscWP0vPz5ZjsAhesddVtTcKpXS7w
sF/HBa9FRBMkjnRym5wlUNNeYXIST5K3TWFALHpiGDcdIuOxfttyPCzFaePMWUrz
h3BBVLLS3COoe+f7vH5p3AmWlI2X/PV2NEpRnyGEAsRPrQ+wfH67eECA2cgYqKlW
jUU9iKtG9zE68vkGgkf79Yd5Yt1mK2NVisvIL1Vt4UD/LEz2PhEKronCBYe22Wlj
mbQk/WNT8TEdXdTpwHfbxxnbrAMu/GBJ3eu/n8yuiPrh5JrpG9d8JirkvKx4VE5N
mXkTzh10VTXUHxEZJAtDZbfR9Ag633L7J+J1FHcGtA1/Ri/RYjEIB3a9rtey4TnI
9F2dRPYQPGoanq7EqcX2fMDjfXYki/fgyLJpPjp5gsvRUqyP6XPUTy+Rs0ZfSoXz
NKWrIks5zSRxjXhLHFW3nx4UA+7bE0E+xy0/EtaJ6S7aAXMAUxf9JRzwrclQslpW
aKblOlqG5h5UFG5UD8Kh7E+9sehjh1I3sW6/QSDEZjQ5jKQ9g8uIdwerXW8c8/GK
2u65W28+ymLqInzJxlu1iqe690tNzsDDgr7/RszI6XvCjo//o0HNL1ftKpEMLJZW
d6T+CQPFndwKfOgIY6KiBHdBSqt6Vz+mV1SlNuQnVJ+Eczs6KuCsU8IfHG+5kzn5
YCks169pyqR7TJXxH01okR7dKIDCZf+2gm2ODcqcrRTvXQqcAlAM0zEz3V9pp1xy
1ZnL7rLaeIbgk8oJXEYu8wEH+IcR6aQE0lkq2sqPAReh4J64KRWFGmTaRmAdP37R
BZWMZ6TO3Ue0R00Fnpiftj9dBC4cLmWYmsLoW4coSQ++Mf4pKWog8Ri9EjhRPCeL
VD3vafOmKJtO6v0P8RrTpdoW8hWt/jtvJtYucU/NEMducnS/cagi5wJ+niqgCrqO
aKvjk0xYSPKbqnD6FRu8Bph/B5fQgRRgYA1hrpL4nBQqCfK7UT2mBSZ9YSHjG7+O
uqmZSpJs/jhgoHCnIri6AqIpvtgNpASiTZUGZIZMufZq8NoTQlK141IIkrrQQRX4
c86IMWkyguy/FuaL5whh6psgBhZyJbteRKfjUuau9QmqTCEWhm8cCGzp11qSdg14
zlw0E61rgzuwgoDK+AsHHEGnF+UVQ+nEbI8v14nMlq6ZJcxuD71HBVAY/ps2/CqD
t/FrS2kuglXFkSrnr7z+JWyThr+2+zdeiZMElyogRNm3h2L+3tnALUzfdwJi9xPq
5gOt4uGoPzBng+R25Esc+B2+t6CqczswrdJJsKZQchmaSzzvRBlzu0VgPhiSmI/8
w9PEb/vRUhFWpR2fSWObS2qhSahOE9W3hUudP4EsfQ+yEYFi3Gee2/omB186jcdP
nvw5s7x8mg7Ja7PpXiwCBhFMW8rqFVBsA85a2LIU3eL/X8WOjxwLl/gKj7q3LEAX
ts33yipNFv+5s2WyFLilMkR3PP8aJvLOTi5awSe384S4gLbD254ZNwAFDDKSSC89
XNjzRqkZt0gyZCLnsyoywd/PMgXQD0s4sTT8A6z/z3XMGhu6QjGJ9JnLjyrn1FAh
fjAJopwaGQqifeSXXJ/oYnmwN/LxQm1EpcM4ZcKtoYIwXNBoyIuVZqBZygCaBj9C
2TwddyS6wgPq6h+wGQHswJj7UeQ8n59zyrWvVEGxS3hga/IzBg/EiWbGnGYAdP3A
/VFusjT8JBkF/G63rseS+/aBO04emzyXhaDqc98X6A+dYjiVWfTz+u1G0xrOfMsi
AF5WoK8Ty7dmt9Bpn4rzwrcrwsIxhItevz+KtB5s5fhwTKu6SMG4sfw32KQCwO7x
h+mJKmO8FACPSUgHjpFOvCKcWLcd4uDITCgbb+vDutX1JU0/4jbEM6jXb45I6K6f
L5bFWQzkgAi6KhvwevSIGBu9mRe6syyEYJMBZdj4Yvqyq/y9PNCvc0t3Y6DX+acD
kr6hfzFkGlGQSjHiY5Myiw==
`protect END_PROTECTED
