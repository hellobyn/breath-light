`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
un6DROUr9hSYYQ/Zu2FpPF8LZTo3I7z+2S1T2aM1DCtggIcs/VskSGcX5r/OAbk1
qowOpuo94oCNkN8dtmyup0QNKqJAblb+5aI+OkubJ4qZC8/5Ze7M0hUXlMgzVhzU
Zn+XUH8a0LA0ps+vIiYASFvMNT4IsBL2oawlKmTNtxGMS5yHwvLxDXRucdkiM7Qb
SZwZ1xmwopNmZlTe3alIu/zA+WH/KFePMR/AUeROJK0apKK8p05Br9xEtxd4QQ+2
J0FUOH4UjHGtlSPvIaS5K/oq1Kl2ApqBuJi7KT5ggVu92fQ74aQNtajbn/u/vkDZ
X8Tpsw1KYv7YweVfp6HwPJAUZ1S1CMLPLECTq/dhvJ9yN83I8xf1tKSZNg5tOTJc
Z9aqwnnw9szXEoA4/m22Ya5yTpbUswUGnI/OTDSAV58gCxzPgS75fbpDgJDS0ZtE
jOafoEHKpFTeYPSaV2RPyBjgx4fMEE653Ot8bfZOgAY=
`protect END_PROTECTED
