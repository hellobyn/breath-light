`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnAhOMW2hKzUOocXq0OZBWvqV6RPWh+Rwct8Q0Uye4UWx70+PCEPY0fnEoS1Daik
0zljAUSbhWz4q9EeBnGSWbAYifbKR7osVzbkW5NXG2Um9Mb32ptmwbVNh7M50PzY
Zp0P62ZX0ONE8we1ORLRHAA0/dzSmF1N/1AKnWGu5ZtVN/L+kRN5pOFHO20hTc7E
mcYygwpnPNj/fGjSAMuuYJQ2Gnl+dthAAGiK1dYSkaLFFytp4Sckoeci3JCnu+sA
BNcYJfGkoXPQTxk/VYrcYeH9zx67HTI/0R1YtQN098laFTcX/3mGPdX6ouEkkngc
kQSM+EwS9hL9CfAGkqsd26G5xvpF4feBjWXbWZc4dUUEGkrmYAkG55T7+Aw1PtL4
vdN+JT1KCBBjB9YF8gpUIkr0V62Y8S5zwut4U/mRtdc=
`protect END_PROTECTED
