`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcFYgioS1O14xEzMfKUvxLOMzXPkdv4U9dU2fXnZxk5iYi5heXK53XhRDoD12WSe
RnVsdQS8Gtp+fh7HB42yRG+BdIeVtF/1F35DjJB3RvA2IPyl3gOH2z2u/20ewtJE
Aj5DRI+1yYVwznhuM91208XwORnxBuBdkUyMiBKTu1ZBVN4qdSedJFI5vx7j5bnj
Io0blRPjVGf8fVyZCoOdOQRcwuULEfHnmKtN3Any9qNZ2QZNgIkP5bfnYbwGI8py
Vy7HhH5RUjA35ZqLDgnC8I2+RbsQP2PgQCQ/h6QqmrHebua8IdShpyj+/OBMRRFl
iFwXNVY3a9YIpbMbPrUKPjveGNCk1XKbSOtsSv9JS6EZzpWt66DTt7hqIGn9LMBg
29x1bnr1pyAxO2xqnvuEugF5ogp78zebSEkfbRiIlVeQjg271YIM6qMknvi8eFi2
YLwq1OOiNxkbmfTU6UicSvP8HJyYhuUuNyMIjpbdROoBdr5fsXjV04lpjdtL67hK
Ne6KCmecDS20KfvGELGE9HoSCvgGEtD8VMtUUXqPhu5sqmc5x2mdRRnTzvrFiutf
fpl+wD6xWA2mfd8AP+43NM4On5mRraM1tpKZfsE7FdUYFiZgjT8p7WzRb4VuLLqJ
cSGQZ4QjhWE+STOiNXPjuGb3B4Jo2TADkXNm6Jb0dFdJ00wFaU3tiNscf1P4Dxlz
Kp56rAuyWjWBefqH1174f0CC3twhLZIr6frpNuMIJn+x6O/fMSYwJ4zHkprO7IN+
mYt5zimcFiW2a3gTuFUtYvuDVdSpKFV9X0VQTCVXJpq4NJA2TZlyN/TxWW1bWNaB
TTr9S8YPsIX+hG5lJRj+MSvRpWFmtF9pVid5o+LJYzkkZZuMy3PUeUux5Y1eaTR6
FZaKe4uhN+eYUJnXPbH5Isx1Xb+uLIQilAavpFG5zLryT2YPlEeXK3dfa3AH5OmL
sXTKRaVxy7JJyedXVtwZCJDcogCPhssMP8qtSNBomavYPw3v1iw/E32mMLDvh1x6
2FvuZyZvL6j1ZavDKkIq8yfLcScD5PTbL/gWFyRVGsBggXlLDga/2kDNpdXSb85V
Kl7BHWCytG5NSSh+1v/cw5wYuoNx1/Ns+h7pOTe5rvS4Sm1b14Hkr7Y5EvSaKnVy
KMvANsLroY3Wunop+IcVVH1caLu80bs/gMMmVgpUF9Fyvp8Byw2cNo40vOrCTbqZ
j9InNdM5LXuJMTSje/OBoGDzKwlZorP2VcT8yfLTIUSDGtxg/hR/unHa9kON6Pg8
K5FlXPZV2upw85sAPp2TQOe0AeznLp2pISp1WKcD79hK7T+MygP10PU8HruC36DQ
iFVvJYnqSWncq111sU+EH5/iqjRDSwXS6YOIZHOALk7MuWyyuHAKXJR55H6PcNJ/
u6vK80qjNmVFk8w3C53HGBaXjWgg7EdH/qHtWQRAj1eKstG2dymUDpqKHI+ymydH
B5gh3W0YASkOE6ucha7LpmFu0EmE1k8mSqBILdWMnL5nmHwdDR1LLhdGWaAJZcnj
IE9+Je476AqRpqUqoCknQSBz/ZIwQgu8V42DMMslVT/Dw3sIr0OoKDuO9Pbdj3z9
0mTPQv5GzaJBBq7FojOyWSMDn/KC0zxLr1up8HH5VkwqlaEe0mYZUCUZVKVxsw3j
yV131GwBG5wmlDyCXTZk9Oyff+qSiWoOqqy+HisMfe1p6cy0WoS0p8IXqPgLiRrm
Hx3SHGD7qjyga68Cmx25ciivs4BIrVytX9piQKSbCr/g6erQd0G1YRvEK7KUcGH+
Xr6Mpc2sXS5GHb3rLPPwSIkjiJyvx02TzxM0u6UCTbLTnwxhgCQAG77rjfol/hm3
JPSabB8+VgGU2hURo24hqvX31W42YDzykfifBKjYrHRv4AX1c33M5dSaGq/kmr+C
A0ThmA5gqiz+ypU7bfK/M3c6wfizZkQdHpZmv3KL4hV8pMwmqPSFYemIwdDka0wj
vV8/K5iq40VDaFK36Yqw3LpSwZle0NtWTc3Kt77ZrMJI8laT1pYU7V9EcLhcEe21
7ISywDORaZgniVQqS3jZNb2D0W6BLb7zKt2gboT8k3LrvhvFh18IZZRC79Ycc6ui
9rERKWWdrp+0WXxL0F1gFm1rqM64y7j39hNhBLs/ywBf77QsmMWJPltSLHDfS1Sx
5P0JLXxR6qYFwK45kKLcGMsj6bHAk7LcrHhzufzTFkieR7velPefBoptJc/q0BUN
MYp5Dlms6y0BgzthG2gOwAlEHVY2SmwTyCBnFGQRsJep7aYAsT/L6PJyNxXD2wX3
ldNFvZw0mIAUTNdVv8ZeVC+4C4rpQUISt4gWRAUn0R58rrg/c1f/h+pD4B4F1cEU
UKsgB/DOReQxVES6Pnsx/TRdE6hY5q+6W+GzfAPoetqhWuzCUKvHIJp+fUWZy4Fe
u2CwfXq7pDBNUBL6nOma/ZGGTpNHsHpZqDrP8/QkXBoGl1UY4RmMpgNHGFUpr3FA
14l7/RtbODVolkH/ouLt+4TELboja35EEnMarS1XLlkz7k6ZYUPYXiAi4ZX+Oobz
i1HsMvxEtHTXnLygCm1BMv1Udfii2VAYdr8l8URRuCgJDDgSSQb7TdVW86EdEBIs
JTHtKO+pGBh2DBtzIeOR6JHAFf63CyKi5BCxxclpTCL5IvSzTN2ooIW2dutpU5GV
HHYLy9QERk0UgjK2IHSmlD8odctd9EAiCo1tg880IVUF7GQVFIbdLZ5TFBbfvrU8
q58oY1rBWk2005ox/q+4+oJDio6tcFf1clPycmXTXeQpn6TLAb5+XYxhqb+/bwz1
9hhlloQrPChb7SalGnO6kJmxNPDueybD56qP/apFXdoCRoHsfvaW6nnwQZ/z20mG
mddxrWSbpqRy6Unlp6SACocJgzYt4r25vpEsbrMqvEbTAJHNC3cP1ELOEUZ6fcot
J6yzKRW2CtcWyTsQ8GgudQdmydodik5V1FJIOAq9AWr/qnU2wNf9RsZMeQ3o0N26
7+pVCpTZD196z+Nh18T5s1k3//B+RX1XGqMsap7GLFbO4Qh2FsyRISDHyTB0LFvu
9ZtKCNgMMxQR5JBHn644xRcBxsn+Uosw+bkYKpZphQIvSW/YWla+p1jN5RFE+r9R
2HWFBeb46Xg+haZFHXyLifXe5GCm3X5/E8Wg7bxdp2Ph0/g7yyS3WA5BIX572xwM
bLkz9fmaU8HMk5qvrSFJDyqmlZzkqzDsUI8MEJhAlKZHdziuj74iw1Ivub1TlaVc
DVgUu9tgvsU8cpdT5lFSIsx2RRRhgJH06r+uuaTi2J3/w2KqW3LdrE/xEhX8QNPf
Sh0S5R9P3VTq0mT9zPMyZfAZq35QNZBV2viVa/q66r0DHghezmDgBkufh28JlbdT
n+mq9eFxBpSfgQ4DOOI2ghrNsQQMVzHLe8DjSg6JTeGB1fwm3VgfhtsybeHsZnn6
hP8a1y43skiCy0HjRnQhz8jq+51JzU7vbrddcc6iOWauYtrMzMNf3YtUkMhj8h1w
rLWBEPt3LtH60UaWG2ujvyQQXBa/FB4RqpbnlA1b4mGCgr2t/yPiVuh4vXjzYqNM
zekGN1azeH/pva5qvMOIz1e8mVJkc4DGu4dC0PbjTxgr+59afQ+lgP5LSnto4uEk
LQ4/GElPXcpKBULZlSuqCQXHJrjx4mZfIb6Xo5Cy0e/cUQhh0vIUBz9Os8t0kL4B
Lrz1pnO/V7aQwFg5DXC/n1hpX5OY0pwcZiMlic4u1BSlie9ORvR/xakOfN/E5J3Q
bcsSlGs7pO+jIKw7GaSFTkMPsTMaM5HYU9alOBCQKYEgdEv7RnVzQvpmIU9zHAO+
xWPF/v1+JkhNGbz6hWz1aPFAY8jjO1bfEp75CpeQrtXH0tRBRr1H8kKa6IN+SwRR
q52v8PjL13Hk/OtvJQeYK3Vm5ev8yZuYCdQa6+IBzGQcGIZHIncz4iv4W0yP1OA8
+5BqspxXLZNFapdOFcZ7vY01CFjT7p6qJqZcbLrwjILEGiY6SoAcEE7YP+bBq9NT
EdxqNN4/gp05Iek6crVGwX71XE2qYZRutGK23LwfseVmhbDzSjIqBfhLHo7IXSi2
JHQ9lH4XGu8Ztw+AMBOTJVoNYcW8fhrOTaTHFrI+UO7jqa7My9JrLunn9U212bn9
DE2IakKthIMq76EwsgrgEKp572uioOt7x3ByhsoKu9U7g2V9xbgXltbbtmOUL/2m
FngQqE/CYuMYQk9iyacQeMCB2xGoPmqgAkdEpSPGd1e7XhkM5xf976N1ZtSbYp19
7N/E27KGPLId8hUVM7Ds8kraaRdXDC8eeFZapasZomb3Qt8GcuRreGJu8xiehJ15
4XR79J8fmMsvDp9LsQSHb/1CebeHSIQovOt4LdI3P4VJn7zufebd9WCN1uF9GKsy
NR2EXkS2OVOe46XSrQi29QZT9dsfjrp0cSaohzMwGwVEieCxDOpqyz6/yRRtFIQW
`protect END_PROTECTED
