`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HrMriHEYBu8KCXQvo1jL+Hso87l+Qw356wvgHSyoWUknjze3lbzgE1b2bex5FcE
nT/7mX4nMqKNB//X4odta06okf3YWRLNPcltWjqIGeCJGUYloqGvTMPjHhku+eb+
zlB5nIZPOr2Yro2/RMqT0yp6FfWCPY65Drrj/2UU+ze9rJnJX0rtrELsSlSZDB2T
0BVJGcFb2J0YhDlnxMnQImKvIRfeJ9hwgddu/IVXqKgZE/9a7f2kMMqU2NZ9ARBI
7hdgsUM4xB2UQpu0rysX3GxUUlav96IMvah2wwUi4QG/EZe4eHllR2y5CDWc7AjC
3xmT2+HFo/Zg4gEkHZnVpTiUlx5y3MY3ScHWDqMkaOO+EVKTbeZdSTxk8n5Ijaql
LoCOskNbpeheAwHLNfWOYWpqQgAUDJ/b9mUkOkQFLTWouQZnoW8YGSsbrJ8P43Wg
T1ftvszyO6brzWaqJSVWMG/Rr4UDft3hf9cuciPYg943OHrold1rMisrC0IDep+Q
UDm7tJt9KHYMWu9wLsd2V3XeQK/U1t/hTESl4+VvQooZiu78BgDED4Gevgfn7uJA
231jKyD+uyU1LnnbxuyPvk0k05XDDKkVh0SLKWY1yIcE+Y09RmNkPdRWZ55aaA7a
tXgoZW0GpqQEqmB66c9kj1kBYpZvCpooluEaUyGqHi3Iwc00S0HzDMh3m3+E9Mli
F++htTxB7Ijnl8uZmvm8/Nohd3zPNWYvVTKo4GyD1gPSdHpMo58+5SkJblgTAFYN
AkwKpyXG2YQXE0rWvKK1A0325+zgxsFZERRWjaxunvVHHgZ/RkVoOjdf6UExkwqO
`protect END_PROTECTED
