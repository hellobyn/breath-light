`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlW2bYjgH+GOMguf1cuicxGKlBG2DSMxJiEcTcqzGrg8fCdoSweQOo1W7AOBvXLs
x2azAoaDBTtYdqPmRUdwX+nt/6Mw+QdlRawSkmndq8uJQehZTB1Id/Y1T2ArhtSL
Zu4V5NY9P+e25Cxdfwlaf6KW5Q9gn/qKEHE1QgcKpeNFKIDE1H7dboAaA9vJGsfG
Dm7NXoQzqcdkoVjwY6bjX6Hx7ZVJKtwJy+I76pYNr2WqD5pNeRNxaRJxJvfkuCVL
RJJQjO2V8/dcop9tkwv9bXyBymOD2J02cTHM7E7My11imZZ6+utyHojcFqeO5NBx
RDizpGobpJSxsf4CYnY7JQ8HDSv4n0iTrOLzIWkosyxEErXsjb6BsWhEVBmI15/g
FQP88bY9XpFggrUb5XyNdgHlXRLJCWExsbHZTkyQ3KthA3RrToZo9U3e4xi1xv59
nGY2zYeNj51CW0fum45mjm6PWSv4yGYiBSNWT9yRbI7Rr5ZiaSZD6FJiQg0OfiXw
cOZRktnLockCzvGmzHC1ILccvT8y4uwu2fj6mFv6j9TDwAVbZ6kqsDwh83I2/Dcx
cDDXJSR/grGYYurJPwXsnFnx5gczF5z3sVIKIF4RSSUi5oaD/gRaI1+7MhN1NCAA
MaZr1xwSre9qIjA+0B4AwOHgmKpPnXAJjC0Ol1jqUlEpf6vrWn07EW5piqXI81DU
SZzTxqJRBTvcaFmNWIW3nWEVa4X5yozb9+C92ktC9sqaZjFPDAP7yAOt0ua1HR3P
OrrsEy2meI1EUVRHIr/7hIEjCLuCV/+pFHRL9lkb76VQT9qQHb6d60eiPhfjU+dF
5YUpm8lBpPtrapECkwwhVHsAJzN6Nj4eKWvQL2yJGIjqnZKzi+uXwPnTwDEgdqD+
Q7uHs2gAThGoc9QNs4T8aR+Xbwt1dYBJ2isaORd7hqBjBV+HZNB8sJnkVwDO/1NG
DWtpG5KEXNL9Bx0j2SyOdoYyMwvg+S5ta4JNWiwt6NrFg02YB0uXIiGLnmM85dus
wD8yu75LA7x3NgNNfC5/W+SMwiWHFC1eJl5JxdjTjsnZyreQ1vLloy+eJ/saSYsP
nBBMOYlEAriNS9Yl98wlf+xMW/uMs5nZSvSGmthN1A5PjkHq3lcuEWPHKTxiZ0sd
t3sDQUpli2+tNnv8GCBcRfJBR1Obp3FWXvt3Mx0UEaeBWTYlAdeXYz2YZGSV1VsP
0jT0dk8mOVMy2DzAxi+yRRywz1N/bvCX0j4yJqNq3oaEn5CjNgrj+M7ogUZp6wMf
uoPXNtW/QJNl7B2A/ZSqvvRcRhosiEhXR9KlPGRVdgoJEMPkcMT0sw2nkc7CPKnB
irPFIzEmBS5IFOtmRxGH56OJOcPUPHD3xovJWGC1ZxE9iVWeeCnwRqUjnPCN09Bp
dyb0ZWmpvOTQBfeOBabHCDiLpeq4WUzLeTnIp0WFOJO99Gcs+zTxWX5kvywYpk/3
P4qZmjxFLN2xN+/DTY9LlMyPHbsCbdkZO1gffj5b3rtxF6SSXDqIXsTaELlDsJMs
Oxarny0F7M3G1R2/rYVO45u7s12liUQcWgFv7Onpa0us9GGB98CNm5KLlM0K+/RJ
HZVpFjM4CHfM2mhZUjKnzismbKWYDvCg5NyhMRXAY7W5srCiAXmSKwSbQJ22fDoY
kSadls82L8a2484EZx/Rum2jDDi6dbngtY7GR1jiPwT3P7d6POyggzEcg39btZAF
a3LpWmXT1De9yjUIuRnWqnyxQyEYxFKt06My+CgOO9kJy7dxCkZLOTkDnC0s9sCO
2+LXfIu3KpL5/YY9WgOmDLJiooQaJt1WLbw/Rd1ed0qIDLm4FZ9YGY2pF6PW+XZi
ycnyFFYMM7fgN7s/h38eHZBT/iV3aw+UFqykh3A2IKo1c+pybvSIAGLIki7MV91p
5+HgSGALiUxa02G8+i1GzXj1UUHj5J/bVUMDO7vGIT4FWqX3kvosA1beHLluSPdn
zswjvoi8/0moZqZf2YUAE333GuZc3RSdwHSjNR3aLlmYC/uex5qDnuysbJFm1jk9
EpMoTjYLRDI0jgsLpax+qnqIo0kgvREgloT9yNapQxSJroZHq9Cm0CE4CQhljAH7
moPwo6HQlOMTh59OlP3y54/c1OK76gLeiJ3gmh+UQxcw9DLYNmQ40PwT84A2AjTU
N2Cz5Ug2rSKdbDTGJqhw7zivsOAM6XJunE0OiYj/RGusRjkEdXctyc00j5sgsF7b
HcBgLYcN7+fi/vFBLCkWQ7RMNUvCq6HTJdEnWbaCwZBDHzKS9UDKXaAE5l9yyAfX
E8pk/YM9WGBPsAD2N4FuqpKiJDCLLr84375kW4lqpEbRN8N2i/TCx00WZpmsbuux
QV0/ao6PuIaevpXzeEZrBAFydd/egTX2yhsVeS5t6ricllTVnLVU3BFGU1asbdlP
8x0x4xm+sdmkKiX7vSF7X/SVQNwc+eFLhpspvu4/ZW3xp/qWPClO3v2YKEyi3lDz
Ic4TIIkVEmD8qYwqKL8APeQvO4EMKDm6t9Wii5rMYZj9quaCzCDSgHbBZBhkRUxK
Bao+gfJDzSy9jodC4XctUe+8r9w8je36DwLXCj0dDS8II/9OFPxZkFrCXuHo+ycp
jKJi/lCCBZDg0aorbGtPBmmaILv4SezszLfIZNyhKJiz/4t18k9ZkATwOZNbvXZU
mEJeuy7i2EuMD2ti0+kO+pFcLL5V6H47aE9XujQ8NTycWDD2t7sBteFm1sBIg/dT
6sIytz+OpQ5a5arBoVU0598nlmGllWd2QAdiDDUvVZSf6eltCVDHL0VzhgKfhdwV
lBlLHB0R+w2QUreZhMjxrvf2Gm0uOOY1masFZIyDQ2G42MjJuKYP5AuokZOLn15P
LJrZZW5opm0i3EcGMrPN6QIoj3urgQtfAbOa3kLsd1YAahU0Wtnm/YDslCa6hR8O
dFV97XD51Z1t8SpaCRN0iddqA5Ij7ko4vDnc3+HHUE+y5SiMbp/xRdSbYZ4nIHnD
8l20X6ZgHMaPaSYoGqz+OXaYgwNva/XNhS9Srebp7XXgZtzepp1s1qhXtdt2WXF9
5bCQWj0YNyP84ZCAYDWBC4yzHp40CaaabHFbPqn/5EpzWSCQlfyEsoYF02ceqfyi
i4o/6aPoMwz7CxYz6Asj7V9t3epKzluFavSr2iPkaIj9SkofK+xoa2CcenV9CFNi
vrVpnFsUlwEBLrsX8tk6bUlc+b0/58TzjgmXoWkK/YPsNH7HG65AydMDILQqgDG7
BPQEbGvVSLwAvHZI15Uq5vcihMM3WgGK2MswWd3GD13gWvgEKUsl7przKAKPV5rv
UfHKGMc8p/5BU3FQXuGXYaHuI3Ce5htM4doKkzKdE4jZVuxUSTzCKbkKgyxKbi+P
kbdJwli21jlD+Je8UX+sh6NvhMCtJbsh3NpUnL6G8eKZp5ekQf/3hGk6hY5in6ZF
6im4V9sDC8Zo+vo4r/AxW0bKYzCsFu8uDBOb+D7m6CLcWaSaGrl3/DvZvXhqGOrZ
Lwa12IPLAWSvw9OInQlLJQ4GI8TUG3O4SpgxG83N0yrT1mlE+jFNZB0Y/7uovTwL
14VMr+V9eT/NZA+lpy7iQ9LZmRaK8BFcZdtzQuIKYnjmTbFA1P8BPIoc0WpbpvAy
Q+NuFxnveFRglIvjD5zYLsVdIuX8Ds9h9rdMp0iaeaWTc7dguQBH0QKkYkEPpD+W
cA3UT+VBU2r8hUujL5fSKDdOKX94tN3MysH+NHWCfTvVsZCBRMGIeNIHfa5By2D8
8ztOKdKmTndKKzOB8sBwHMvXmPHSLQ6cmbN2Kde2Ql+0Af6RwNyf3voIkaOzWuNg
/aoBKanqWd3jh9p/Cnop2/lsb52AfXAaHIIviM2AVzq1prT8uW7cSvbmZSSnDPrn
IXbjjz/iOAcbJ3EqGaaiv3w8lvGAtrF+eEeKc5Z/qrnfmeAYmwbIJmOHJlt+MYH/
fudCrx+5nbQASmKBbQgfDgfWVBd3V5yOyhyXsrjkev34CAlXBo5TQa4MaX5Babnw
ume4QzSk7XIPx3FpvgBgyUuK2WpO6ANoYJU25mko2+eeqWJhapci+hC5ezH2c2zo
OSVkjeXPulHEi4YeXomswzG9emSYSGc6a9vuMeVV5Q13HmCO42pU0uEk0D9DhCoU
AhgemQSnFAwNlnv9OlebtAAbCsbX9LCBSrARR+7//9WB2hMovq0n5MlhFk1AUwYJ
Bdb2s9y2a477q8IcGpPPSRL/vdBzyiWuE9PbpN/CX3K8UXOG07YqClG6S2PQzM9g
N77yU9fv3vWDqzOCeh1EKA6TW+Zp/stThVAOKoCVdCjNJ2rFMZDS8p0dSgBGrSgM
Sh+TqItSf19hbrkNfKrT+CgA8AkSpvm46/or2/RASlw3kcnl2ffAdPKHsi8T7gjK
PFL0K9+yrTd8RbeFyrLmfOa1pSY4/qsLZNN6IugAwJfd4BjQjtAL+1bMsU905WEa
pFQ8gcDxlfMQ4Z1IAnBdxPZOPqKTOCa0hJeFCP0+CXdEJG1MR5IN5C4VVg433pJQ
zbEeIrCATiFeED4HnKI9bvxCToyGWTdw6+csZOfrNovuoqV3L0MCFLR0HlYWAjPB
ET6iQ27Cx1G61PmD47fRpo6yaNNSUtVEgZo7LAaagrbtWc+n1SuT79faWXPQYbtw
f2ZvnhDvqpvMpIhsiZ9C4Gw44E2zfW3EeuM9GAcaBL5IBQzeRjgj3fffG7Eh+fZ/
x+ZySYZz3X8yAqOArbIjuCQFqG1T8v5PIbPmTAolxH69HBv7OjJ+Kyz5c+v6ZgnL
ab3+Kbaejufxgn1eOsbj8oFX6b2U/58vqRkSTlDOqqeKJhjLbLAygbgSchky1A2g
Rp5/3sXXbUswmkWotWXwrLCjjBnAtBFC7upQWptwgY8yRBcsgeIgjI0eZnIg7lFa
k9PFB17m/FQf5u1c0igcBMrFRGCC38zLiPpR0euBKyIX/zxMjtRwZShy73E65Pyx
DFyAsXyuPS2UL5n75GmPiZ4BLE8vWfbJgZ39mzUjIudXDlUZizmmSZR3mH9zKAL4
0e8hgER+FvMWmH6Ep6i4OdlS4CLhXlffGIvZnQKiSwazmTB8/CybrEDuZIEDBNDn
WwYsTcYrXfradIBK6GCY3/rON66ykWy1agZC92fFiqCM7mZRg1KLAhDirQNfMVfo
MY8IFCNHa0Uiio9n2agAMb6w5IzavPI51/2iiEyr9WFRxoiDndcosuN3ulZI2Jpw
FjgZuCrf/GGjWVxSQah6Xs7Fxo7kJgxUTJ5pcIx9fE4fqDX2SdbkZoBexVBr4QcU
fMV5CCFbseVvkl9oNBmypo4AaOUo/obxjoFhKWxgdJCYzop8ASVpoNf7UJmCoJj/
J0vV300TmZE503WsScTKWok9OOGnYvJTDR8PqTQbcWz5x8EsdGT88x+xcvG1BT+y
GUbJMuKFwRjkALXJQeCxXmgcfzDIDS1G4LZ9VLmvtqiKkl2gI/o713mOP8DY2DPd
LDOmG6gB8+yBc4fTXFaxwarxX1XWMIWt0JMmiMrJ1mwTPpayA2H2/XbYGSnkJXq9
KgTkY2wEQFY4JCm6WvGursbaWU6htOf+yGCnv59xUCyVopx1CuOF8ulDfPJwMe82
+dmVqJofAHX/DN/vCkAQ8p4eS8YuNv+mSWhZGv8rq675JQKgZrOP/PoGR2wks/A+
ViFSZpqNK4ERRvQZT7OdMdg3A9reLv1wvRcT6ncITsFggL0jhec87PUF+kqAFHrS
4vbBuSoKJOPlIMeHtAAfG0pAFu3ob5m+31oJ4nbqju95ByLIrvYMH0LsNiq/QM/l
0WAvkj3MnnkalV5BL2eaQ85xNz85fdfjWM+a1Wq5eOxr9XRdCZjOnCv1aDHIU6N3
Qo/j18C0tcT2sCnlBHb8z/oWj4vr0fD/BWb3RUVT5n7WmnfzdXP6u18MNAHnp1gn
2MKbuut4v0mJM5WKgTiU15pz2p/+8MEnc8GGWN5ONaeJ3gJIyqImag55RxMAKoZn
Bc6cFPwMjqHxVEJeNzXJi/ewsvQe3tOV954XhUFaWrTtv76DBdROsD/c/Lq1H2rF
jNiGuLHvAR1McCP7W0H8PYjgdGTfjwrZqIWyjxmsytvZ3wHjzvVSQAbainFQ4APY
dKVjamqtcaW2CilGW9mbTg1KEYAgWPEA99bATG2y+807+GukpeVM6NqawjiIj5MJ
ZedlHlfCYQxtFrxbR3ftmFpnEtEvHXdQi3mVo25wUD4Qu/QdyxYob1o4YQ+MGbG8
X9sdnudAb+/pOY2AzK+tWPb/9qUOe4jdCF9Qh+cXZN7zbUCxNzgVU4nMbjLCdxL3
pixBtDspuGdpU6bJVCFIIGay+19IJ7zy0NHYdbBn3aJ4qgf2S+omgjgam2IsP5Et
mi9+J6Klqo+p+GsqsQ3XYaO4PfWItetjIjqCFBtZvPVDQgMjOqWN2Rf6T4tJcz2w
YrDzeMITFpJxQ8z5io7oq705p6nyAnARyMVmebirgQpFCZpZ3aGTz2qJ8HolQvvu
27LddMJjOX/W2abbcXl/CNc+HqKueJ+d0YhMLCsegiWRmQPNx5orNVz5bjYxpFv0
fdQqte+J9ybetwZZNUEJySVDU+C7g6C8+Wq4j4Xf348JwurePSW0Jxm7injBxFI+
Fk23JXKqaW/variskWtzEDNmJxmxXns4MaEmVrF7qHg4gdA+HOnO5FqqOTmB0xIu
mErUhC/+ZwIfMR1MjoYcpxWoqRjQvaN4v3dszxbu+xiN8wwQaE7zWeZEBDrbbzmi
gOUclYYjpH5hXTg/j20g6F6MC4Ti+T5sE5mxl5gmth9VGJs/0NGkmbGJZGL4Kp5M
G7g8GWnAp06n6PJ4yC3fmSlqmYKlL8+3yhepFSY1h6teRB+zo/JDPYRsVb5d4cyD
v7zq6GWpe2Su3x41rD7tZ2T/nYpFUt3N1tMwEAaJQEtOGa8G8uHf949dUB/ljaml
Ym37wxjGhCqKUQ+shaCYJxWVhcaZSWq5OBSN4y3aSE4NtAEeDsDDwg7KpjW0eOhS
vR43FpWehbEFy/Bd8S3V59xkhNGS9ee9zBWJQ8RL/E5eCtqO2lNIsOBtnyclIM6z
wJVIgOBDmj6OuXBXD3tdrN1jvHqSg3dSXnrUOLx+87qMEe4AJewpaAAS+UTSk2JJ
YPYhW7jeEGoczzp2PGkyJzZHYB+1/wuEAcht4GtDYCl0JbU4/GoePg8QIO1Xh8L1
MSQTCqwW+czdDUwRamHYmPzYJsCFpIsjzOlpWZ4I/7vgTwNV8AZYH3ePxjrEHoiU
JNRLedlR/wA1Vm/fNBF1Ste6Fk15nJy8FmSE71Lho7SChYajfuY7xdwlDPES+oKk
OCyuGzbpl72lhleyPHfxRXO3/sYeyANMroFvBeDI82B/K8XnY0RiLrXE6oWHAvQ+
M2eREqH+cWx6O1wWQa0WuaMUczhIMg+vX/uiiZuKmF/y39QE2JOOwkeN89O7c1hN
jXAEW1I48GHuJiRkOkAaRIF+q8rAILfQns9HuAEdsui6CfSUxctGgf9b7WHvjjI1
z+ajAzfv8NsS1MPIAL7uOs8WvqhPqK34Zmgqmc/EcCuMQfEkhSVMJoXtHOqZJ/wJ
vDZhruTOgcd/w+gpMr29n32GlvHm74CtD6mH52Vtn6WilyD1I+9yaWXM75oL/TIF
OsGPYtIFdc6h1CxlSPnz4lFIyNUaDgHt9XuCbFGbPXWF5xw78rtLcemsgEWX0h0O
TWKVaPq4oT+i3wKMBCDGALZ5cVWa+H3nuXOdZv64mH5Ps8dmLDqoEJ7eL2M0ZrGw
f78PVev8QJZVvBOCdG4HZWVIPQHn8fS64fJdYOOuFOhX1kPlyedYHa+CZUrGPecW
S/zFFDEB/ah4U0ezdaXrMy0WV8ucgyzV8XSqNcQ2dAZ1uwAOMN6LGeo4o5nQvmEm
S5oXCoiLwUuIm7VHaan9rbfl0kycuLHTA2RPwkeEKU2VjeqUSf8soqZIZ3TcVj6k
9V9GHvjeupco16VZaf16wWbPIv0mvLInx0pJUd6xbTjvBc+J7M9vx7H73ndrCuKg
FVTJpLVu4Z4EPt1KsJs1ldJQFwoDTnslDdPfs+AZhGRrzPSghM+MiL5/2XcfHiZl
74RBx3f2qhy89u/F9TGlEJk7Y721qo2xwTRs3FRfgqJDai+LlUnGYFqUa5ByKAxa
FXKosemre4SyhG7qyZXi7Al0nvvpQoWxt2FxxnPsLdd0Trrs0JrzwPf/ie73GWK+
U6rkiU8S18WmxEiWwC7YyZIrfrzLKwZTIexgiEE3QSYYJQ9d5TnRlhBEky0S/S21
PtolIPHQjBl+Yj2Wh7BVr/bOw0xyES+9w7jaTQWesPDRS77UF6rofWCNdYg/43TH
32PFzd6aY81RMFewPYWLsG+SvpZxLpZej+Vf904UQS1v6q06IvXLa/Pyph2QeUCz
tmnCjmHckNt7lom1mCIghSyTsaIa/zhwkpDO49qA8bbC0taxt5Q5kzOAoeAuBo+K
XxmpBP15vW2s9zesmUzXdEJKr7uLEQkP0RppPxegJbmdYJIzDVdE20Ca9x9j76Tw
IDJeKd99BV0i7niyThZKSkTHGc9BVs+4Ssj32NnlYSZZOfiDQmkx4sQOmsykFfvD
JhutP5bfVSghB89giK9FvoGNXweFHUwwirq4o2ByZjl+x3hZEVpsY1jdhVb8h5WP
nPW+uOgiXdAL40M1cXv831LJlqhpKCEFWJUM1r8Rfd/7z5vjPbjxgzhRaGdq2rBj
CCz/LiLrHlzg9UJd5k8oS5WyAXYMHVBC9rgJ1zplU5HikaJLXcUWnVW0Z2ZELscr
doc8K5WCVb9KlQKaIpkdcyvuUFswokBGdCcA3+wQKMKxM7biT0r7oU/iZCfvhxCM
y2cPYoaF7t5m+iAXL+sRIvQ4AhRe9UImZhYMflNW9ak/ZPPpEldJmdla0WiUx/Yp
uw9b469ZwXRWQv8C/4/K5LGGDx/ozoJF1B2Z8cZsMG9MVg2YkiRdKp0Ispuz+XdY
5ncpQJbYxShDQ6nPnZaBYUzh7XzyyY4qi7fmil0Ih/6N20TwN/AkDHWlt7RZhHlH
A0WfjLe2/hFHGyJsyGuYP0T1LMIEmIrWItN6pw5kzzdUVWhGBe07mZYaQl0hwxXa
H5C0+4zfnlLFDRH3flTgXqteqbCA1g6kltW+j4CUMaM8gKZh+Pne8iKYNoLsfoil
elU38A1y737MJTU7tL4okhUOF97+mo+Cjck8TDPDQhXySgto48aOhP1bhN29Gs4a
63ea753Gqhpj7JemJpMVL0RcUI/XheVH6oqUxuiOQPeAn1tt23iy8ATyscfqTlXw
qrax9hMUV6ud/nEQz++SKJEDxmt9MHeOFIAi5UDk1g3Y1d95oDarMUMwNKge4MDF
DfN/Ne4kxGIzTkDWbzVmyXjEUYSp+olJ7yeMCMxMMjbNojmM8u/Ty2702RxnHM2w
MFR2zGIK+gINr7/ea4bnBKllYpUMqspRglx2qqlC0XlF3EYZQHk2IwIxJehLqVip
vgjRLF6rLGI+wY95EIlv9lIRRvx3iGvwJfh3A/EtnhjXyubaMfMc9YUuUK8ULHYS
7hEhd5iBTBhhg7NfmQD52JBSVf1qPLU1W8UkWOibbyweE8o+TQdgtHwBmpSkA5cK
HtWwu7M7Gwh+Fpwcc3CHanTIxhmnMT7pBkarGKWeBsBxgW49p7AoKjN5hfZAHTD4
KI9YbkVMLJ08yUZ3i6lfLbxRytFXQ+UTJIV5tT0DSG99igmNgyo2KM1iWITVeOAA
slr8J1PMgcuGEN7qjXQXKv47M+VymHEtJkmV0SaFaXWXzD/hwalyijoxnpsV8lJf
H+siZ7w+CCb0UOD1n5ucvYp2YqXfPTN2VFWLMsWtmH1qYmWkVRHweixpStsIWFyW
La84zYCdmsf71kK8RcFLPLPXvYw3ISVFknLUPckMOK9LrL3egRkJnwp/Af4RdN71
69esxXHZidBJfnZ/Us0ph+13/mpp8/8Q7CI7i7jbc6k9dT+wzBMHIr7MHqbS3bsT
1DBzOp8gHjPBgJV8Rv4sEV5ixIf4jxgJo6T1UJL23QpBcBJijQ0podSOsSScXJV2
l2na/crIBRcyE9SV/q1BoNZESsgLSLD/ekycO5AExQ7NfsoZ6CwJcYXwGw9xbML1
+bnB+1vX6w0Z4DEutRpvb5XyvwvfuALCY/OL1yiXTLlQf2fT6eC+gukZPSN3tYVj
kbTMuPhLpfovkyChc+AayKtnwpvpqzt3PV3RiVcryIzWou+PUjSVsOetsV/51qdi
2yumtUKH3jB31JA3vQteFqB9JyLe4pHZ8L5IO+wuiJlPU03okIfNsjFcJ//U7Zwx
YAdampAjrbB+0nm0KTNIvk2QKO/ithJ+PqYK05To3vQlZVfwgo1Wv+qaP+qdEi9K
B8yPUtnghLy+n4KYEsJW092FnIYaR8KgIzX2uzK5RjZD+aFxmjPzfTYrT/KefkzL
mJherzuQpUPKaRNBQOoKZvqt5ccGLash9DU6qE6xGGtmKmNna8TgyWDwBlPTJfXw
r3K/ZEWFhAHXbU/oiKZeQqj4ZO9nrFXOMFOE3MA5Sk92KWcYMmoV9nH7MldNWvhQ
IoKmecvWRHARAxbG776ju7SEJVLc8DuyDsKOeFvzGn8xsdE0cYatXhaTWJMoEBsq
0TmuX9V02/QyGe5NCIDbRA==
`protect END_PROTECTED
