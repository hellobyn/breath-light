`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4EjQsksj6MpiR3L2P8RdlXQBZLGYu/Vb8vjOpwMt6NAK8hHbH4NRxDVZ4D6uEkz
E6DOWaqDi25GBQYkbeHJnV7u6G3cUC40LIQ61+HdtffJakhqLXXIDSLdO04y5BvS
DJ3ACiKFLpplUPkDj/gobvtMXeQdclID59GVodgA6qla0BILjK8sumyPp+MzdvsW
puoJoFw3KVDyhLSzFDzWLNjS9abfJiv/sK4e9MnaFJwZhXPudoP3eZatHzuvlyRS
yYQBGRJKJH2rbG77w8ivW1b4KOL7FjiMNTtIicslGWEpxWmnQvwHF+SHybqayQpG
Po9HUDEMyQZ9crlNQ8/g4nVHm0vOlADKCVUUvNZRlTR5R1SmncA7tc+6yJYh8TeB
xsq1J+qbvW4WiruXuKaEovXVk38s3jJKaHH+kMX+uHyjwSDJ4s452JfI6NigyRKQ
8uKwRBdyZsuvEAZhDLgDQ29/CH4Jsf08IBbsUupFakk71X+o1cHjKkUDjxUR6i3T
h+qIVAJR9+fZaCIRoFICM2a/l5mICsZ9PDfy+KfUmzCLcbjFCvcI0IrMqNV0fU+c
n3/xeheQUxkfpmEGo5t2FNR5S3aYw88uZcVYJcG/4Xjuwyqm8VRiCtwCbWfb4hVp
aFiRK2WPSv9ndVmTecdxdC0F18qyqkL9wv+S6OpoZMoY9fM0hH6UM4t///Y/m3AS
3PKeGlCNB7eZO/KrjfEeThDUSZlQBvD8gk3v9WIvgW1EloN12YXCuyxEEfIb51/o
z6TtMbtIXz7Vc5N23/cl3srKQvlapcVa/tl496mGxMUR1Esn97WYzA572yunxLWa
mACc3sFJREagLVo6hsVxdj5TuncZ5PEDhTm+xoxE5JkNNS2cQSM+ify8vZqRuYFs
owFjsavzfqdsCppwgcBv6wC8DF7YjU3Sl9fNy9MYV9IFoh7OoQe4KU5YXkm1bIUN
wQBjZQYLjFYzzRgnktVvcTbBnrCSDr9/2INIDhGxJ6N1/zALuzO4IdF6qoZPH1aw
GzO9zfCADwt2QCXxGqGSAieHu3AHcQ/aQk1UABbyd0KAs7HC2y8dNhMyHLEE2n5r
UZPn20Xj2Gw+ygmfjXojdUhJYso9Hp7zfoF2WZcMVMUDYMa50hD9prPY5dhaLaPa
EaDiylCfMu7s5uIiNrdResG79hrSyN5tkhwML3/KFf7WXTI6NFHLjTXBIadUN8S8
J1+tK8IeMkXzzuOuqyWgQdnZVMph2Cz+daHyZASevqj7E7mU+a6ayQ+tcCIehrTT
KF1LFQYO7k92cow0cOMuJcKAOjT+ErnOdGGy8PIJ2zfLukyAmczuqvphgsDRbLib
ISpgdVQtDSs5VZ4IHm4iKACeZqou8Cup6msUI1o8CzCjyKx0U/vFq91hc3V249AI
PNAAsrRXuamwhOQZpMjIChTOATaFwBpHvMeMUiWkQmnBCg03jv+ib3sMunm4327P
hhxA7KMrKCDrJAkxoI8vzFIHQWgM0YQxpQnwpGxEuQQb9OVtlRlmJrASHB5zbW9n
KkENonrJ2zGNXEhOwR1KYfebgXmcGtkPOTAsOjVSHNqML+bFCgHnS08GPvg+16UL
PgB8TBbT2kgqHs1u86jJfpMykz8V6taXRDB7L/NxxglEd63UiTgg2ol4z+XxlZWl
tgR9Clsz4snRL3IrPXEuOHfWSYGRcSXRuj3MrUJ/cE4ngLMGcLsIj061qq3GDRkd
ojtR8tQGqLbgMvlRQ9Z8ymyKj8Fz70e1HNL172oY/3R1i4uyR+RdJoJgFyObeRZq
5zNOA1bdQVszKL5GhoaBJaaPD0IDVEJ0TmeLjfzXpf78zmj+7pY7pO8/caahNj6X
dRt342Ek+4sifUdDouW1AoQ4P3VLVyWPqgJM8A2bDF/zlYd3DmTx3HtMh/iETS92
lA0MdL2Kn5s0b/tGj4QOq1THNY7RSYqIpAVaIx4QDxKe3gsHR5lZQSFaLCjtq73w
a9+TNkrPWXZMzmFExE94IFbuutxNhjkbNQut1Ik6Pdsb5DpUdp9qfjF8uFWA6KcE
SfPu0g2arlk03WsV5cIn+LZUEhd6h8QZpSE3KlEbMwLERkIhhp52ZCKvTM1jqTDr
PPOvjqQ2gbYuB1spzS/63dljH4EYWiK+CSrtJjRuq2+2LtHjczdPL2WJgKJwHYj0
ZTi0DTwnT6R16ReUk4G3nPfTSkS4zesQThlF7g69cFMq0edK5yVauN8HCzfq+vEk
OMwPx8T7XRUF8gZz0TYeLPlEif09eABQWLvFk+LjQCzfn8eOJD5jsaQc1+mCsFo6
JzF+pIDjwRF9VjJaPdy313gxyu6j8QS2zULa5OTCemK47zSxKmlK77XhwKf0vl9x
rZpS1v9HPB0GS1HAKMnoWH4K7nM5eOJnYeUjASzsenTbGUUPnSlumBh/HC3W0xeV
ws0HXAtUq1jzSqv0aGTRgVSO/7MMcdBf94M01/LETdiqwCWh9kEhUT5TorNVbobC
LLhogbLMXVX6MuYFDrhd1I+TjK8G9eUzkW9W64GWDLFRXMJ+wci1XTw+EoZ0o9Wl
n3cUtWaN5gWT+Gx42AXRuaJesX9l0ANYFsM533iHj2/13X0h975G0k6SU7jUsR3s
LSRaLs7woEdf3fUcbFUNQ0bE7684BIRyOxEk/dboeUvC9NVob5uR6tlS+7OxP9bu
4o6rbo2covDcJm3VBs/Tzq+tyLopaZrqXwKfBIzZ6IOkMI9K1E4+mJWryBNSQ3a3
HPXuKV9vSTZdmEqqKVW6M/SpPSRoIBzwxz6dVfJTko1xvPxAsoDQnb1Yt+Ct823o
s9aW7RNnbGRWEqcVODLnBDYBms71R9bvjgzSdBJWdDbuEPVzNQHIL+dQs/GqI9Ch
dawNmVoGbR5B/n2RuxVWYHQo7wsLdrErSlX5a+o/KNVULGEyph4bV+6KmU/cyVaX
9gpbX8UkidmQCNb2fZxomTco7S6V3N/n5XIVefio4XSQwI6QRG1AdbUpcpOOEEBt
gT8iiIgMBf+5YvccRCLQuEcwLr6rFaAlITXResTn/Cq2OGH/acFaJ/wKE6tN4Kot
qo/apUlfKnzkkOGHcLWB6ljPbzUfh/l6/7csN4Igz/v4MBGYlegdeRt45x63XJ+F
/UzmKAmXOWREdEsPB+s3Jx0yMDcwsk6A6iYLthZIYMa0MeBjLu2+0YkwEaUS9x+N
TOkuzGQboS5WGvnBQsJFTL1PZNI4SnMUixkvk2OtHDArS/l3mt3E/7I1kFokJkot
cCpZSh5YXHOdfb+0In7oartyar3mLenRHFF+ReRV+qs3ULUWeeIqy0K1kfQMQuaa
GREPvMR4jpOfdgF4IbXxU9puGQrr8qoRjr67GCK+S+iXiTn6wCgWB9CMJAx3xdO+
7m6ExM3mWMrMxbZ7Mp82TxnMmuYnaCMjDdGK6Y7BgHkPd0MgG5GrsOZnYSkf+xYs
EFQcUu7yqB684Bf8559tpAnQ5SZSpjdWq/umEc384zMiRS6ks2iHzmEIP2dHXyGe
7Xxp+Hmt3A6pZ0hWvaLLxEyItS6Ky1gm11UzxQtloExNRc6CdicT9xbIaXbzWaLg
Jc3Yu7A29WkkB1pJdAePbU+K80E09tO2XeLkfqohxuiHyg6CTazd9iFA27F0WyTx
PC3uXwMdi+4tnJU8lPowh8b0DAHnox7um6GqrUolkAY4QLq5I20ZFChPvts124m/
8jhfUoWt4kyihtscoXgwVrb+kPqtGCImizSOmUuD9e2BujAcTOvb/Ji3fDdf7sIy
VgcNEQVPFX5PiIrNvlX9edM/Wp2IOIl5yNeZQR10roNaFbHbqEcPY8bZlz+GYpAa
U3vXskm9aE7JBH4bTesnxdh0jptHkryzZdE7QMVKZRorO3opTsK9d0Ys42IlktAC
89Y5pID6libLXzZI8SxJpSqpOW9zDBGQfVaizG814UxyQGKCTfsyI5wHl+3E/gfe
azCfSsu8/olHC/5PTzdCanuaGNz4w/URq6P1UYPtGP1rSn9Qv37ormsqRAOXFB7Q
0dBtKpm/JGtVe/QTAA/MqvFRKEt1uT/ZFcp3Yl9z4SecpI9GCLT6/uq5DL99VLou
Ee2CQgVxGJ4NXtsv+9fvuc3932qFlljNU/d2xUbQWxrfURzy8VAytKIM44wEsKUa
9Do9id2IvXKUoq7XQhwxbtHvobILUpRdMKzZpSzcV4j8UaOoSlyDfRbGlw0dY1k+
wXBp/dVOXuozniBd67bQzlhT5LSZ65EdD0pQC0U+t18Hz6TDLimWFMz2YH8JQ5q6
zFzKgzyJcQ8WtvlkkKjEMv6ExjKSAcT0gJhXZZGhAAtx3inqSyEViga/5Ywvh7Op
7kVpBBf15J+uOOAY4kBN5XChTgQHX5sQE7jDAtz/njw8gUt9kZnbe9fC5wuEtlQw
mvb6Ss/L94XGhrXye2ezge1PfT/wZ5iZ9qf/Rn+ZKHlYK3yc1BEBYugIvkzO2dga
2Kg/nzqFGxIUykdrK62nh16dCmRynaiUwpd49Gp2Yu7kPbY7MuFSQxdgxz2x+LYZ
gBAIZ8hJBId0olm83b6qYUBgLT8omtpdZXVLFiVHa4Jxb/karl+IKL60GFLApwoi
RBYUg3GnpWTThUmh1x4rWow/PyZP2GytD0dpQZgV40F95vdYmOsoJmV5Zk/mBOBl
wV2Ojz7PaC85c/wWIdbDQRpXiz2EferJnL0giscDQOTHOI/Kuv8yFbqRHrwviLxO
QdqS5+piHbZgRDaZcSUXT6viY/eKrv2iEoSNaow/sVZ9q2aw1VwXaDUMFuhl2EBe
Gci5+XwrUppmTy7NNpT4WRFq+Q7XfSnNnVBaWIbfCvl02IPkNKYGylmwlvDqU5+V
Gu3iQliBnTDQT0RrBUPKOkrExKhQMPDQWZ0fgQ5LjkMErg9bFo1C6nC7Ez6Ac8xQ
Vdv9FoyA10MzrCdkW4/qmQ6TEv3OIsOQ0/qRzIuOfIRd5hWr8toozS3xOnEZGwyn
k/6nWzo17FPpbDWGi2MKBTNAsb73OTWm3lGYhzWCxAmdEcNujHN4h0Q8VNVGvk24
wGK3F8QTvvX+8NSatR7GNYxL6xKsb1o3E7ElOBxdvLHAKvBGMKQrDgtwHeyzuGN2
rCYhh3lcNX2BKQYbjDeS2a4vePbAEQnT2terlVSgMXgOwrWsqgQ6HcXqjGZX8h3i
vWfVL6B3RqU7jzJ2+rRAzA4DnDwefbHJDKvgj2bM2I422NcwOw8o6Wx3ClRqRhLy
cGNWmKCrTO/Gqe1QFMA12osZptjCnG0C0izBvh7p9npmL//U6ofyS1aSkRXpQt24
oD+DlDrB3Qd0FK8WWNn5UVIkc0lQE4WWFLeW8n7FphbPP4c67Xrg/viiJlr/g+9b
1W7ImjByAJ3SEb+cfEgKdUQl7p1wwvyjuvwt218F+oCkHeAp08CtIsjCNZKCheGa
Sflma7k4hrXIKEIfEg54Hd+ctU/TFfxx/3EjKrIsrp0ylMT3PonEBtcar0Qqmv+7
mKWHscomtR25j3KcFryc2nvxi5+NJi99qZz5CTO7/svUo44o0s2JxNYfMSxUM2xk
f/yrqQ1i1X1yw2yKsfEYKMTTX2OYwGjQpt2LCnB73RbqInPomf5T8A91/QKmZlAe
BKWWpK+eAaBanyXU3Phn4+TOxR8n4q1DTrgyGN00dCYG17Z04g5cpL4Tn6uCSWnw
2C3zBHvHGkWnliyKF7FblpliywqrF5NkvPaP+hsSxeNWokn2jz0MKJuv/3kB6Dpr
uWmehGgbPrbyY1eXTJ8WkojF3YUgJVjq+DnqdtdAqcrMEkwDtcx9SwcO2+kPA7AP
m+s+cH8AJdscFmo9W0bZYyD72F4UeC3XLZ4djyaQyrzCxy5NhMZeyLffZQDAhruL
uA2Bk7exlEJZm8PRUDrA2jMWhrjG3B5YvI+liG4cNoI0wkcB3shxBJlHWzlP4uEM
dI3UoW00+cbSDhLLdaMBmUd2POInKEBZfU6s1oz4DTZ2uQvuahA6pod/B03qfOIc
5ejy5QXqc5iTyAPLqlbnomPKkSJaC8MFROXVjs/NuYVN0kBbH40MbW4PJqdndeT4
E5XqA0j7gQUBjREj8Cs8kQ4reJ6uANfdvxlfd/5Hjvhmxim8hrZr+yFHiBE19ZVE
PB86OLKx+FwM+oM1IUTuirvwpCgmyHbw6Mb6y8QxGJRgwKATKU4d+gt1lB3+y3kt
m0tKUKN9JxqIF7tBayW3icEdyIP2VZM1jr7XnXACdn4n2EQWFzDV9MjsPGXmFaXR
Ez4bX92hI26o8+svZK5rVBfyZHCWJ2qzi+HF0OCGHiZvAWuXedKBnYEsTqmbo3Xr
C9VEFLeo8Zz0+PtfeSO5lbobtD8RsiUglzUoKnsCs5Ze9KkTCFQhRDUvSSlxe7hr
0lsALRd1Bzp23PjL0R4wVL5EQWCC5eIJBql4r/45un5pvYgQlEcixfuQ4MhH8N4S
nZ0HQj/VQHVy238qtZxJ16O/nSIA2HUF14OEacaAcRjyd02v1SyX3O4mKMfVwviH
2f7c2WsBPq96vpGRnvicUfnXL89v7HP5ku1Tzj1rkOb0XmvyheQz+j5m6Y7qzo/Y
pclLqQ9kdVIizXDcREex8m6EymkchvJIm3G5a37zBSzGeTxLCj/PswDR30kyFXT1
qXra1PNoLfRWfVbC5mgY2oe9BZQuvqK5UzyaDfVIBYXpKVERYVl6AQ7o3ULx0f47
q/a8iBIVMEnyo2CnyBC1XF/yNxHHipmFjBNd12eRbApxKadDjGKiBPydCkw9q74B
b6lOyjH0AwWJbf3Tqa/1r50kt8cA72jHoFDfpH/o1wqveUS5J/PwmwhLMHYIEuGF
fr+1Btm7vY4Mk3b+vnh24Mm5ocfC6O5knpUnMfdcDM+zHs3HufhpwV4cqDS6ZAJQ
+vMFf90dI6cmkk/0JXVZn0fzw8DvHstYQ0p8Q1P+53MVR/IYQXJhYpbM5RRz465G
dXnhWhFCPoShEZEu5az9wtosE2ioEkNvlZ0VMkuuA+wG6CrUvH5LOTwbLWrSZyOk
g+lk0zr2SWNTxqRo8czMQhODhrTVy1OX43E5EHcrnBMRafAWWNdy1Fo6ePDdxkli
3AKwBJhkY1Ua6cIVxRPl6uShPSKsI1wjswYGGBUaKDGF/OpG+8xdcYzhoYxudVxk
WsiegYvxBfqIpujpkxB2raqPllKxCCuniaLhJ0zfCjGNgKVwmlDbXv4eDmy/8sJm
jwLV1ovBQWmAErhzQtjIt6pcDsnwVp/fxxRqqJuNDAfnXCem4/5cxF/rhoPrcvlM
OL777y2kJhNveN0pMpq+iJ7y57ZP+ccyJau8T4vtkHiSEYYNbqsmZebmtEtPJXJc
aarNA8dUUP2FSwUbmJGGE9BN81nwCYz2QPOt+OBXIbh/x1KVLFMtLR+1q/OLCToj
ZdZKAvo+OxDK20XeJwTdrBuffGpXk4nA9kd3pxF8EtDArPFmXxGcvvweXp6yfdX/
xt8HZ0Tu7OBM+0GoDX0P+iew7p7Fs6weIX+Scwwpn3IAHnOFBTmuYlp8QseM79Cy
xpStF5btEyjoYzDso/cF1Mq/ItuhrZ8qS1LFt7+ff+YWUXCCBjXnJRwszEY+O3If
EoLU0NSXNLKBfZ1H1ED66iBvb/UA9Bw5Qpw1TbEP5H//cUeDRvDMk/v/4TTBQ+Iw
qP+FxCdTDnuINZFrcm9wjOo5AG+v5mmgWgA0UKotfEEF9sBXl/YxI3G72AKKqwTb
F8KqG1yPDd/PF8/7tsLFmeI/MV2gIdzw4T0O8dlmXqIFpGWtBosWTE5+KIHzZpAi
Bh8OSGomntFxJR2GeieCK6Wr2UF3c2Uku8JdTSuVMPqxd/KIqHiqpPOpPPwuYu6r
cd6hSzX+GhfxeLHi9iWb1nofEnK2vDdm61Z1frzPJq7thO8xn+PrIjlL57aUk/LS
INE/v3MKeGDm9X5IiX1yejmfF+wJR9AlCQP47j2aERQPd/3HOnHkiIvt3GbcR7Oi
UK0ZMazpI6QbTCVn57ZprOFFFASpxn2YS8DoMgJWetJSe+g+mghQsfaaw3VCCNIy
8rt82cCS4DSOn4GO6nfJn6+pu71F1/xA5lyfhDzsxSck9brbCoORE3BIf75QGVcc
+0za0U4KkmC445NZ27zTkqmwsHOiYQH3fMlVYAMfOHaY/9RZ375Mzho2r6oZ7ol6
tSpsWKi6N0T1zF3OFZlzaeBy7X4uql1wo45SXmc/Own8FJzw3AR58C9lpzgqj6XE
RanAhMCcoIYzvqO4nw4C1F2egCSwfHgc5qzrYvCSHgF+03LHilPbwDFd4lu6ShR8
EKdzTvSlRgmGyJwQN8mlfF2ptwkNO4PEihk0ZfyKZgndPIEAIU6dTlkItbVReLVv
pYYgRbxghfm8ag93CNvxaquc0MFazx+OHdntzC5UGJS26hYHdh00toRSEtgVQTqJ
5FwVVugUJMxWzo5pDxASZe4TzvGy6fRHu8YbO1JT0ApevJKN3kCdeLNjGNFQGohF
yFFvbFj//VvBXZFR1/oMUAwYKFuvUTfDPSzTbog0eU3VmdHlyHP7HqSPascLfKys
q/NAjaNMvKkdNuWkPuFpKXSIqEn38vE7r1ofT6g8lWKzRkDT4/XvgydhWGDNkDBM
c8AaNVX2jNrRPNHCKFxoPAQkXiRzouF3AVnc10HhtqYLbOUNcSKgAmrWriLEhCNd
KXWqaHaieeMmZKO9uw8S045f188ZU7ImNlbLDCltx/WQw39vYgAujxtOiaproSO1
cac82IcoTOCC2kMcrKdonXQiORZuGEXeuh371a9rNKfPg5/4yJ/IaI4c0iHInm6f
AwYTNzfSpPlHo73UNqob4mVTlNwukT73q6wxCnGo6JsEYXrjRkyuVni6miM5sMG5
gfRD5dq5WO1TeamoEJxfWDOlxVnVhIBdg1zBoy306n8v8i8g2kIxBGFzklcIggg2
BhblrPMoGWMmKinHRdcMBWkkILvb9a8YgDRJcXtRzjhUEZ2uS7GDx9Hwxhhn8KAJ
XQVp9YSI15BjrgaAE74dlZYHgthFQ35OH6gcoEbJNs7yyA0FrP9ZSswlqMiytdMU
Qm85hTpl62zieJQrh/DK8cAppewocmx7WwjWh6o7UDvN3eq5V/SvNhfjXJggPmhe
Vxc5Gxgj0ILz69iVCfrXQAPyNpzjBSyvwo2WvRi34N8Rz3M5cs4uUODu8Yl/3lb1
8SVuID5Elu0UPEDz/VH4Yfi//qz5qRJVg5cyu3V89T8/v3bzUWdpZTlWG52aOoUi
vA0Uq6rYJIA1o8CIaukHKqfBioutLK0xOpCirjBy2lTegvGPqgrwM4lymi1a0FsC
n2D+KUCS7u1W3SP1Dn9RrWYezOPNajPuLudPeuy3nnl36Kf1V7siS7JuTeCeePKk
ACD5DgSRsCtrKcWau4DfowXVAWHpO7X8xevQ5+vKJNN9+28medbgdpLPn0OU1X2G
lP4dKG6ke6C2za38ZPuB3TWUIS1O1u7uNZplOmbHn4bZAJgO9h9jIwZXeBuWLBF4
bhY0cfOaLbpt1vLvNZhwoJRej7jdSc63FpIzwSslY8sTaMPjLdGcHiE1VDbfhyH/
e/x4i/e0k6PtePIUoVbw3P+k9ee0vVsADK2w9mQ+SOjC3FSFToRUQ9NDAOZD11jW
a/pc/GpgugXIHEHxuM4tfHjWAGMQ+WSMKPR2UaF4SaP7d52C9eYcxCeu4qUWitpu
9zPZ2GsF5lbEBMEGNQdUZ7FlpuYJNgLExKiapTdGUyWICZeBg5if+/eQHYJ78quv
N24noxYLA2qSaPUoOpUC6OLBo4AKy4Wj/npdeNwRe/tQBpvRY3IbpvBN9O73TBWr
Tx09N5X6lGX7+j3BG6X6+Clf2wg1qpliNH+xJzSHlP4RaGe7a+tdFr8MV3K8b4KT
D+g01Dxs9EDCZFpf6ETEgjzTet9QhEYP961I67QKEKYHzBswMstpEQZPGI6F7daf
9HGsRYc1xBdUYEoVBDjeEehecVQAPuE3KzyV3NxxGyFmcU86Sf4zCFLFT8BLDRir
uA4S8xJoQmIYlNgiJ/07WB4B6Rn9driLp6czdzE049Bg06I+D/Bc2CBjGeHuATSX
ATkaC+yD9mNQw1/6fl3CZHbFbe+D7UQjXPsFWZUoE1dKqS0ZE5oFArVk01Z+xEvc
u38F0jGfkT2Ey1Q6C3ZmcezyF0G51H2qWKo6DyKoNHYM3ieXaMKqoqJQYgDpIVE1
mPjg6gc01wTo0N8Qb6uiRoCgwWdB99kC8uCt7XSeJEip/Bdfm7EogPnCA9ueGCoj
OJ9PLJeJ6uObMlyGh3l7bkgHFeT3+X3bcJQ/rMm8ovedvqNQl+q3UaXGkl5FCIOz
zPCOAIrYGYQ9nfogR3Go43M8j68XC7+naHjr+ckantO5uetQlykwvaqIOOOT2nDM
KE0L4d43z9i8qY+mwsIe3iXphDNyExFuDAicb5oJujtz2Q97b/fZ6iTZUwh/v2YP
fw1xg2WmP2bZzDWjV0S3p+FSa/lFPjkcxE0RnAShrgpSAvrpqIC38us2RjH2Mf0H
BRk7ip1cXdh2WyHDkslf6zBiP1R7r6OW3q2OVgNM976E7h+lX5z3xtSdMC6WMl+/
QnwJAzKzZcBh7+lFwcKiqKO7HMdvBv7azLts1resHIK6OMHuFdB0yRK3i7YttPLH
6KvYiFHBF6P0T5+YVZPs11b+YFQzMJ6Un+Z9ZlQrYEACFtFQZ70laGZ8iAFUqAis
i7SW/N3oLO0mvOdydKOagXThdYjnNdBUN0Nez50vKgSWphvO67YBTFmZFKqcH1MA
6Lk8iUEoC2RsoBCMzd5C8U0Ov46cKVYzYiE+SH4eNeQ0/d60/udqnPtfRv4yPvxE
5JpODC0+YIigr6WNaP/cISnLyIwIjUz3sNb1r2ZKSJ5T8YJIezcn3JFmU+/qkzrW
eSQ+g5EHG+o5T7NpZ+JNQBvZXtS9+w2hk3TVc/wRuVQ90FoN7nVvlHum7dtxfBy6
1WaideB6yKIo/cp2zxVCZOVlW9suUyt37oOVYKb+M7MshoYEoWZKoLPiW1yW37+8
+qd995F9Ewr4FkmjMMwWteR+IkBv/awSd0+VQWdcRxVGdfssfd6IH2iCaNVqFve8
R9qOxYc3PRuJv9jZozWKR1NZ8cjxtQS6s6R04yEZiTOVQjWmOKsN34+eKZ6CJ6SB
zj/z1jaKpR06MCFTuHJlEqdjnFFPQa8MY2RT7EP4fD5YxxtP/sntEOKSm1r+wZuW
20N69y34ObgU5t4V/4afya28WaweHEoO27RBm/z5hLVAvwonj84cEBhM85ZHt2NZ
OTGWhYDjqnRnlppusRJnsmaHtmK6tiDJKiy7CZRo4H/fjVuy1RNX7C43xrBnNcgT
kxEEoL51qjXUHLJoMFeW474k2uT2VRZ/KqRgh3QpreG7jLqYESe1r5Z2MWFiinEG
hQIYxZEQD2wTPg9jWwvEk4gFXP1LcJddv49RxwLMc6oMbVCf1zIxmqlEV+L8+Hqr
BwN9djpisL+UB6pzHHkP/Wf5cxiCclzAM4QCR4IjfEqVdzz6aQ66u2uIYCcNM+L+
/LHRbVTEHLBMGzv3O+KhAi7ZXvv+eYZFtoaq/FmQBIS1+H3nTCaGUKt2XhoozTSq
S7w2f6nakvqd7qBXyRxVRuMtzcsvxymTg5o0GXeCid6emIbMKA4RJf9uVDojpezy
5mM57yQGPSGnu/CekdBky/GClvSbxZgaiy/HrOip8U9RNyO7wsF3f73XqIUVVNVO
FUqNXGU0NW3Ikx4o798MST5ehN+u0EHu9VCMdG4GMCojg1BCWXVm1hb/RHsaJd5f
pc2nw5g19D//LFypKzk68RlSL9qCt9If4eKJOI8Z6ayYkQCId2+7nQT9+QM1WstH
vYY4n1STmXiv5JjDEcXCwcvpHXPl6q2jdzcstvlABXPSVg2PHxupG9IQM+NL/iKJ
VrWuGoIsmmw8fm/5KKAwTPOiuLo0ADPNbwBKx90NY8Kx0S3uVTW/FpvbcLn2FeZh
FuykVJQEmQsF9JG0RodENV5xjpVExBtD7h0kOL+2UwQfYktWfncXHwq2LPML7UYF
LlZfDGrIbrKr7v1ZhnLJ+XCUDsFGrgW5pSkyPqhnAvZqrF6/cgk59HTXClwNnGHd
ghETxflPPD942tfj30R8mqwCBsKOXgYDYoMcfbW/RHmsbZDEPhyn0iIkZHP5dLeX
3tI2TrpAFtRLNtnVzL6EsUnnHdjrgICtZEps4iRrxGecldmXUHc+bJt9YCxG9SkA
y/Tn9Twe8F7GazBAliFzfOQzlhdl4UU25NRcfHIqubH6oA6BdrlHfj1bi+5fdFCj
K6isWDYuA0BPQqanHoBwILTPlvZ6b35+T5wKzpxGZo4BauPTYb1+EAe96Cc3BXMm
BBJnaEa8txb0+zZo1VLdW5PCEP07mGr2FBeqyWpn+1jvrXaVbuOKrn+r+sW6qnU+
/jB9C23YCJ+H8K2dGmST9r0EL5m2SxJHu5LGS5VZ1jDOaqKzVALyAnO0YS9JnGAP
ttqvOy3b/Hiqz6MwI51cFrGENOQq5edgPRAQWVWB7kOISDZYFMY+LYCFfwCMD/HI
H2rsPqUSTcpXhX16hTYKm6Wwk0X7eY7v25GJ4+Aby6B2NqzgJSgn+C7ZtfVH8U/f
dMO5//wx04iq6fm8/shYMLV0Fy3I4iiiRipscJJQ8/aCVvnBaJ0q1Cv5DKtpt++u
GvuwOflfX9SyJco/+rhbVQ/gWNIdJRklO+qcFXPz1j0/O5ZpRWQB1BPazO+igmez
QD5EB9GMq62iGNPQrygCNXBkG0bxsZ7wt/Lm/2eXSeJ0Qa9neSP5N3IhR8bBWX1S
VNHottxGSF9u81kau3NO0x7QCBWM7focd7UcSpTRceIZyjFBEYAs5nvuS/YF3WlY
FKoOAmMkpcwKa5a6gz7ErZMQDEbmZoYBbd6kXvVikJ/BEXqWdtr72367Kp6vQPer
6LECXxdMbiQWkuw+a8t5AwFCVRoxuHuj5dZwSA9zHISnDWyNNmnHDnm+0su6IY6C
VddBf+prxETVJsNR7NAaoxE1+Sthxg7RFGkZwCiiv9b0ArihH5i4Get+mcM4DYx7
UCIDnShwkgPeph79DtY7/xLtt/EK3fqpWrPv5j/EFU6re2gT+KT6+qf2+uF1Wak9
92B4GdDpqvaN/sHeg4gQYaHvLd4wHK9lTn0VktmN3uQ05gckQCeBcgZxs0kFv2qu
o1RgsATeSvlVxMHfegl3WiNjxer+iUCu61WiLS4GlO+YjbuWmfs3xPJpqH/YSpqa
vz/ZBZ0kvTjeZjFx2vlgTvOvqG7ElEXOjv/AL387uktCCKB3lL25+6AIbnPTxxDd
qRnQTpOloIZ/9J/zzJosCugAS7AqHFrmFMhkOeAC2hnEC95EtjjPy0FZ6DKuiMe+
C5+n//o5/KGMt9AY9efQ9cslu8i+taAeOAYJ5GghJCkEp7sW9hvaZgEFoebLS2n0
TOFlsZ2O6CCZN96/DLRGMPth0JGk/Ji1o5gOZ5dQIk64MmwxZIo5axYVsVrFQ21Q
kPUOsIzCAYBpBQweIYNAbdyZHhHgla5majLU9MDYPzUEVHWtQhKiBKFD8o9eUa3Y
8da2FNPgJwmyEKNuxr1M1GXx69iVoWfu4kbhtggnaM84hVyAXOgiDfazt1u068ut
pt7pWhTDoOaKRHaYlLFJ3PmGRsF4gUpSkMODj09OT0wMSA144TR0ajkyU5f5LW2p
ogM4Fnm7dUNKpjfGaA254ZDLReS4eXE7L6U8x9Mi0dEYHFBdBZFW7OqEqBYnouMI
x8ZmZLq9GR7y+ievXpHL3epljVmYjR13OTdC1fBvodwVKrQEhhaEEr2iEPVpj5/N
SalJx4SDcO56gHArGOCJ+w1ARZSpjyMl+fHOH+LRA8/w8VkVbxTAR3Vl/Pwh3YZY
Ni4hdeW4NOZtpHiePyNhSrz2YYImyQFxES7rDOFee2tXQRxgABxXdpP6Dl26ayVw
lkptfJzCryXDUJefE4UwRzGO0LD2KFAdsrqeTDc4RPPFCYgQ4XqcVB91eulz9qMA
QNphnOWGlctC3NLWoLyPEg+n8oLDE0fdlcya7tFHe2xu3lBNystqNnp/mAb44ltx
QBI54szv30bvGCMV6r3i2WKScNoZnKEFuBMoQhEa9kRoEx/gbf4zM1cMc6D4qK8K
imAca5aUSabnw6sQalGR5PM4J9HyFK8DD/uXxEBX51LkxOe5eUoNP/QieOX1HCec
qkZiBqmIpoReOUbZbNEgqxvW7Mr1pSp2kPDKI4w4pZOIovPa6aQ0ejExZSQzLWh9
XA7vxqTOQfgY4MxQGr66HGfNvU7oOupQyTBqOtZP4csjVrYLpuHHIp7bl7N9vsJl
6q3XjX4ZiVSSEk/2DaMj6LGVtFzkgweww2im5NJV68kehC2xNRlgBy2Wj+Ah1l31
UK3yKk6SW0lBPTRF2Gv+s2V746ZYogS13xTGwcwg4F8bKowtrEe0WnkyGHutlIwp
g10hKM0mkTqz/tL4ZMHf+tl5n+QFIiNe4iM+VjkphfGX5lyYDUNGXhNieu4CBRGX
/EHg6KlD3zzjfPhd+UCJchRWbbRCY+2hYE2IdCWDJDDjIgLFxQKNCoQOcXhHdfn4
coulLT/ZENHqCGhKNtQik9HyRk4WdXRV8iVnYUJmhHK4KVzLGPpH9ACXTb7eOOBZ
zMZuG0uT0XNWl7Ns1Bmyx//D22cc5St3EmiLZzsz9Qmz2opil5qG5b6qFjo9Qr5B
W5YRMImoEcGe5+JuVoISW4XjTInEaz9nhzz9RL3OlBBs1RF22ie574nefO/KhykT
doVFXkLdoxs8PtMIi0WpMg==
`protect END_PROTECTED
