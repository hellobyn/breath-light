`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWoteedyWgwCWmW9XebXsZ2OTqqyFzch4dnx5QtINTuHyOnzKKitLCzTe1u+T2Eo
OJ/UwpvtfvOQLQs7cI7GDGa9nBOKh8vaKWUYnK2P9cJmYaVTgI1HBwyRTRYXE3lZ
AUlFqOxMXPLmMPQ9r2CiF0v/DHSUJsJUvzUPfbtH6x4oRGRlHqQKIyXwXl1An8Bl
9KnNwEQtb75nBUuzFBkmkHSsNn27sclEwVcdXkP8Wjv8IKM/wcnqGFCxWYu/UiiB
8M7lTq6sSh6JQ7A3eR41W9V+a+QOHh9njDmroExjpyS2xnHh+2nmJqym57+0axCO
DkxQESUhCWx6b3CD1GJrJI6AkCF7ZskQcitmqbG9JRWKF0iMyerzMSkHH1fQahi/
ufx6iWq1B/mMIC+jAq1cxCEo94m3/TCVWGdd93fceeKWJV46MqgJXO0fB5dNuI3V
6tz79uOhfJpAjNC+8X071Df890fjGUcQKHLHhgM00hft1v2KYfsdaBfPG6DPxDn4
hecBKAWL0F0JZM+jqUq9i6JK6Jzr9nNmTQT2MKvmbryLfc6hcRUZglwk99/+5MkL
yK6XaJv8dJKv/MotmX2ZGK3lAEgD4ouUsumdAvOGMQKHLxPCELm7K41UKeGeS0Z/
WFIsRadLyg8R8wXhQPEBj4y6HPOxTKyDChv8hThzBQ6I+hWGQEjh3/fJ0hAYNXdk
gGiUr/KhgpercbnRt+QS0sZ1/a+IM536l70iZjZBE92QaYAOjW2G53ztM/t/6kA5
OZ08TNWqLtwkKroGDzNFcODZ/dWrg+88i7M6aNwTTosm4PMccPEKGO/zW19HcJZd
u7NfYRXPNDtayGdovzOzg22TzrC0qS4fHIuGZCQ/glEIvETpaoQRU/vAAmBdlq+r
eSRQEdlA0SZzJvKPTkg6WXPg5cd3vFh1M+NDW8yR7GsMokLVXbOd9/ajSfC1jCuB
qdyiuWhaL93OLnE2Cdcm/ZWfJArCF0urA9Pm98tawZ17xQAGktVc3RGJLqnRjg8c
n3TgZ3KKzERhbtovfb3+gACHic4vNNJFBUGCQOeHGIIjS1tDxxt9Oiume3Rpla6m
8H6r0NPgH4bqvyhb9dc9BddWwXJL191paVL/q2Pmw5HOOUe7hc851ec0Sven/Gnt
1qpQG4NrmZgMXW95xzNJ1oJj9QsDkUjOk3mzZnH6zRK955DBDImxPxKVzx6Xu3Au
VR1xQ3V45VSvypIeFQ6gw3jwIbWLEmxdy9dfGUnRAULShaHw3i+JvZaXgfynU9ac
FjZmQCsT5Z2Dh0zLd0U4Pm6WYMkzww7ohHs7+3YxFSbIy1xy2KpyMEVVaeJUoBAl
5qGF9GwmDcMf5CF/wQoNCIzHYt0/6xiv9GdLdbdTu1yro8QF7vPPbeR0GbwwlS4+
NWdalLz0MlGBYbBH/M+tIiiwGYUxzcHRuKLPGlKViOTA63TfjSZwtl31/Pyqj+fW
ZXxrQfT+sXDSB7X2jJlatpnX91QDPDRK3HnaP5uyeMsP948dJH1ip3eXVe13elfy
2nB1orbrx+HIQ4oHk4zhsMVh+V6OhCS4rfPLs2fK8chPgljrMhJf1+gWT/5xdzQE
GyemDqqkH+zCFLD3MSgaJa2usd4zYQ+YJmhzvhtoMkaNb0WZyM7Akj2/mWON0Bz+
OO8WYXSwI65/nHgzjbVesuancQuML5H3TTGZ68w3c/6vja6inwX/jvnyDj8W2ChU
fg9Iqps2mzEWTOjI9BEfs4bsKzd/khlQ3KZ7Umso0NyNda0pdZC/qwQ0ztRilMlt
14mQuTCHVI1T4XJtXuv5f+FtWjO74dQo/z3GrvJA4XMzQRIZ7T4p4rT1VXbSw8TE
L4WFTZz6ICMx0/u0maThBTYRxfCyApkV8btr1B9QAYAqkcFeC/rk4SpxTwuS2TiD
b9cwEmm7uY2dJWxXaObwyXzae9FR15d8g8F/B4x3PrN7MpZOSFxoeIC4g37nzZQE
esOkee6r0hxPgghcGu6tC4AHSSCqYJnzWD6Th1APPh9Ttq8clVVLBIguEk8+Wt2o
quAiEiCPcLi/XwV8DbSi6s4p6NzDzTqLjWGxwz0W5OmBTuVq5MDkRRujCLisEq8i
LHHx45iPFMlTNogpfzZ8z9I4XoywPWkOX7v78PZMlpScVc0AIwlSW9Rv4CnPXMwn
L6pO7nyVZP9No7syZ+0Ex3kFcyHvaKROm6qb51egzVFzFFjcGDJ35RX9z281emF5
S4GnoG9fH5sDLQkw4gTqWKQfYh7ViA91wf99P15NxxIeIsP2wRF0b/5ZLXBKufK6
MvKIg4b5lbukgrYooPgGkgDDGPNSCvH7D/SrO7wLYLyUkifVOZJQOgEAgw/dCDuR
w6jJXuVJJijspRbg6Pi8K4EjTJBISix/pIh2ku+opB5EURkaWUT4ODDJayRFikdV
bzXRrnzgd+JGC3SVb/OzcyPYGtCzA2M+Foe9NhN8/MrSDLPscwFnIq2K25wtPxTe
FOxoJSul185mNp2bQTx5qFp58l0PAdGWogt09ndiamd76tCqGprdjgFjVQ++t1gc
QkhkQfNqJg7saLfvRDugmRDFneRlWJCyG8P3ZqvSN5pAAyPjYuGUvmPu43aMAMhQ
/ii+slZUyhcaDycsWfgX7eynJu4f7sMBtw6z5OOKf4MBDbg3NRVKKg4JasB2rUvR
T+T+KZedcX7Y+vb2TEmhwD9Rogo4cExW/DFjrlwtuXH0/kLM6L6yZkbdny1cU9jK
CS+A2zOS2Naf469TydwJ2GArF0YiRTL1RSrm2DCx2Fjn2w/+qnC9vIkar5LAwP10
jK2G7iqdpkubcsdRPuA/WUtO289VhF/gKHJ7OzTod/Pha0JfIrp1ndSk4sdnRMrf
7O8T4TFtIfQcFxrFBPzzqhjy0xpkrDmQhD5Up77t1NgQU7GCe3/AaeYoiGeWBQ45
dUMOy3Hrsy+EFfecPrmqf2FP8cf550kpsG6rV6Q/vPgQRn7YRvhTQYPn/1scUFPI
siLWMFZJxofMHoSRpTxXm+KebLgMnop0S/mE8uruTnpvdo15Bh4EB79hmht8w5m8
kCmAIHCxzVGEctHekmBXQo5DqawCJ3z5yAuAvl5L/6xmwcneBTxOZHvkrinymmVR
1QfVEZF9yK5iGfhaKvRQTKBZF6Y216xuUr1+3vsVjVux3aD0tGI/OM9HuLvppmd9
1yigzayBNmFQHtaXpkdNxhG4+TvGHcwacPSsojWiRWlZcTeKrhWHUDtq6u9xaoNc
2r1K4Z+FYd5SlWozWzJy4k80DdZRbs0Awl3SotUWP49ANI0D/lxw7QIMEiGOWP/1
OCMu1nTccaIPbiqRuVR6T6omNv4QwNA/qKp2dkynvac+5VKzUYieBFOIbrUjDAFi
3a4OpKhxk+h7PXU6WVXa6vbvUU6No2lVjK+M3BdT8oU4zkjKSF7jJh4hN1o3fkLN
ibguaJYSs0mpW/eEBUJj9Wsx+/jSYcUErNTXtZ1OjXNtrxsF7DZFF7wZT76jx7zh
jnBfqPM9aLnTaPQEFA8LqkGE1Q/DBb6jCrs/dAvVsii1s/IM2HPqA6ScSitFXxuk
0Hd05+IL6fHlniw7hGHOK9KQ70FGnkL2AVSGPf0mgRYdX/YP4ETJ/WmPhNpVWDBV
fnBzvNxB/c7qr4+gybSvKNEHiC0X45lMNpkZMl5SoxEVPYs8AZ1ljSxbzGdLa85r
lh7V//7isfsoIGtIZ7rTBnTtK14+XwVFkCC4W5zCNS2T7YfPe2vf2faFCny5W7Dg
GwqZ2OAjT7dUKMVeHU2ZxeTwdVqTpOidGJxilSnoZMPJZGz/ZhdFalIY7yGaJ8vI
WhXkup879YvpuwUhA6HTi7UZNJ5b9DBf/tCb8+rntxKAmmb9TZj3pglecnjVFmyZ
SrNg829CaiXS0kpARxwI4QANA0FMrjiI2b0ZZGC+AomlqGp83jIUFO6qiDVrVBK2
vg+lCFqMYwAvm1dW26wVUDroNYTjir9SZurLVtnYIhae1e2kyyisKjrPXsGGqnQQ
NAxLclWbbUDNCVkhvfkAAGrz05N2YKRe6zVjl/06klrOhXa2rDjGqDd3+KbmKYhj
cFfMyaGn7Cms72RIIAwQfPjoXKHXrTjUeRlV1nE06pcRbZmiQS2E3MVMrbT4YY/b
1VydcW/FZRZabJQUta4XOY3JHjpijVAIhwWG+7vQB87HFSk+pGf2I0Vma8vTkfXG
/LmYNfoN+4Vo9nx4C4d6t3ooCuW+DxcT1pFXnLgh7og2dzy5RWyBb5B/QXkKlMrb
UJiTR1psX5hEMYB0g27ecWBXgp5RyChuS+eJ5/d6KOd0EhYWQ6IJ/P7Ju8sH2u1r
2CzXrjFFgU6eDs5+lZ5HOHDk5Q6hfkJVkg/qYG8k7n4=
`protect END_PROTECTED
