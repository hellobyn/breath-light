`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvUpV9Lj4KjFbk1H8b6O6oSqdOBcoDng6ekutWPazHh34BrUtGqRblSQaUhL7eAb
WH0b4mtT+dWlYB1L+d4mDbkolxoS7940EhpAUlyp5fCSzveC5y2KbYYoGUmHoBp/
U4mJ5Dv6wWefobweFZbkpxYefGch3mKBWuVrEgB6E4BUD61/Ig0MIlaB4BTaDaKR
2cTmv9AGjaiPYBdU8wwtpi3j5hp4zJj/ztXbGeOapSgFOU8i2FpCH6MCwlLZq7Z5
8ZBeq8OixKZTTGMRhpArywQpHH4HA3nYxQ6omdmjbOeZ44DOlEld3Q8r0ME3LCJO
2ECCmX/KJyLqBqm8ci2i1Hn+OwGnqTJgTIg+Yf68UmSFEBp6DYPrrMbeEoP6H1Ih
TwOxx2b20JotsE0UrzoiJ6qN/NVt3VtDhgNsxOKKSL5Wq6yGhEmJywssVCI+EFDT
mYWgRfpRdhOABGimp6Qne6tZqmbzYwL0V2bVQr0QAseVTogsW8aNbkKs5U38phRT
EKoTqGmK/WoejrklezOAdIIn4sutk5jW227WtWcXckBJODmhE7G34MLpGRbKPafE
Elp9mth7N5uucPK4p5YjjL8fqn63xmgJLUFNkIWU9Io6Dbtj5grqxj88PbERksAa
qBeW0mooC6TpAFnmo39Zwff/TnR4gThGIdBtDp+3hYyCdow9kD+TdX+b3qVkrwHJ
GFMN0Y+Em5U5V1+OVl06KPHKI0pxR/zLoOal0kOUjTMCWUU+sO0mriqW41RIjrWc
EFq7krzn2Ktb6AY0Anq//BAn1KkTrSCFsARE4xKWI7KJTjem70huVyN2QEw0gFdA
osU5HyAdO972ThZo3WF1r8/sM/1J7YnLUk3YCkccP2G7ChGT9grU0HM4zuscT3oy
UJ/CZFZoBPpG0shqjVqHFe0zAngnslpJFYwbXKmoToYcmQBxl4iR2S37r2jRRqKN
VxnvXW1k+hms4ZWOFvJfzJjWXwatmp6R+zVb09B0wcH4t+SfmyWn7wxjFnNrstvy
eYXOHUPYeIOemcLIjWZXLTxqmFx3arfnTkcXBs7fKAc3rsBb88gjiM2LnAWpro/E
kjOhIgxnEBFemEXl1+8Fv7K7Fu9j27xdVzio1J6aitPo/A0z48FOxWQQs/LyBrRj
LLdkEePyqlf0549Ezq/hFYbsRkZaB61IqL8B5DoXbhbtqNuYhtsgHiBuIFtAhzTd
htPfzWnCAh7W7rJfs7+gNDSgp7ZGAQfP+HS2H79yJqrr+02F+GvYRKKYCvYYoUlT
wu+k4XIKBFXwF7UNejC7eHIEEbdwu+fKxnX0ztuFaEij5hm6ETO/hTQIVZNGbDRq
HM7P2pLC7PPxzMF0bfoPeRa2QRrzke9NLxkK/9VcfZ8IJdKan0zI7H25FZjt5q7f
YTLu1PHLRPdbBbRVYGk7EqCD82cGkMCMtVlTJgqdGSHVJsm6/E8snsWWiuhHcWXU
UPKl0HyCEFqTjU66T7QQaRRs4w9wf5nQHtqfQx617wA2aus8W6mxjuncpDXpqBlw
k5NNAXFSVs/v6wCP7U6InPWWp+Bx362QBtx7AAl1aGtAReRMvyckFSq3P/+suh7+
jLa8dSC/AfKKkZ9aKqsOpgPbqsJrMg76EvMBEmmPiBxpxAHmIf2qqRnNWPpPD3x2
FvDTyZ7QrWpZJqeQWaoTu3QCPb27t08SSwPt/azZnQdiyaCGHAjcQHeaQi03xalA
rTik8v/JGtebIJ+RQ1kg+f2laKb6uKCKuLlvaKNpX8XQMqZTqasiSKzvTRGYZ3Vf
kDIu1zifw9fHDleAc6HA1o9Bd4KAmFxLe4WTaiq5lMzwV6gJYQGepNXU+H0AsSkj
qXT1FYjFud4qwW66W2Eu+PneV4iiL7PXSOFV7uTRl9uhYm7rcJUNwi25n/20M2ix
uKBChvn2OSpAD2VOfDSx1Jv0LT8O0lS4+UIWo/+4+vgSd6NaDYygePf2sQo+KQ4M
vYNB7mfhusJOhvPqJoszTbqhR81EMmAEV+XB6e8aYmyakDaptvU2T7NuuoPhZEvi
D9PwSDe+nhcEXFe9e3GjJ3pujMmWWM6zelNyby+BsV/5whw3/CpMo4Rrs4rB1tqw
uf9L37ZfCj2EB0RXK3zXiQTTiLeROVILXF3m4p/7yYgihNMyjOgeeqHpDkaCivCR
QvQo0ljMiCD8f71vAWBSRKclI1Q3AlSMW9qLN+mxdN1EWXRY4LAU+LvHwVIwSjS0
mpHIppYhZVdgVf/vsAC3OD9dgoL726EziB/0FvtOIxiiXLUY1sbhHeGJZXmzVn4c
c14YU4JBDSlmCv/SR0kELEr6GP1aR3RVRZDLarWQOdicW5MUP9clYjsPEsD6C3Tj
UFlHMtO81wH/K/iCo8MvGavowMFadAr8xVO05lu1D1Y/22DjDdOUiobweTbdlhKC
Xac/xf2+sL7HqdeT1ggCx32tOQ/gsjDYgDYQj5d8iIETDwb/EmxGjKLabEEzWcHt
TOpwHsR0iRXQlTQ5nGMXZ2669nWeIn8KZjvfuj9/QFr7yq8U4tp6EgSkNLu2pS/c
CB2BUqwbphnYOBeE6zipjQb0hSQJVV3t9KsVkhimT8MHYk2TK0ZeZ7pYvStmP6BM
G9JgQTvalEipijiexsc5YD22PvS+LD33qDiKlia1r6hLRHO5eQgVYSi97I8WKUUp
nwoYoXVwuTpnGlPnTalOQFDXLXsERhPi50sT4tzFoyk3e0a7Y7V/yhUrnprYrh4M
WeAdz+qTk02XYfzdg8c8nBs7Git4aYLRLph2QKdpAmC/RAqHunvw21tCdNxrWWyS
+5giUqysN4h+aJ9+kyJuoaj2+DUNRxaUgoM8Z/AbsoWl2z+vHSwB0NXAiDcjYdXy
e9h2JDpGjCdoy4i6Hu0XfZucUt+SBOS3NN0z1DTu9krkSNMBUcg26SeqaNWVEKbl
IU/85q5F3WIqHBjdK29OPvAwfnWICrO4mfCntkf5ITXnDEmuNcODjDuKaobKZWap
e+2c5jUH70n9sk/bHFNk5cwmgsmQOwy9zBagZ5hSvQPQuVnCr6Lx4wNoTmHvDSvO
KJV5fZrOBBWmztxDrbOepBWU8QXALAVYgU91a/RuzFYPZ+PO7vGR9Zfb+M6MU/+D
pkgTUKhUv+4JEbJKRoNpCUdMqeJpXs2ya2Xaf55rDkI2asRSrV72QwAZXehRRL0K
2jrvoQLNnSMro7Zqx0UGSYktQ2D49fqG41xE2I82shXffeFWkGHrAMD2f/F5sZx4
ZIbZQx2AYD0AnhDFbrjDipbPl6FX/4wRfRnc0RC1w5nTCehopGQiX5J+Zexpv+6f
+gBgyTEJ4bVEJq5FsI2YBJwT+ptbanb0+HPeylUsTEC73VifcFljyk/Zp8HgmBms
QC8NguxScmGJ0N0iZieGMYzgui2RDhsr+KArRQ0PovSNbo7zaFyKMnXK5m2ZLvIY
xMQlp/t72GpmW3c4o+f5toweqD9ox5uOII3ukQbbDVTftdVRW3l6Yps2yPO+lIU7
sPT8s6HFHhZXIsI3XT3MiuTb2TwFgpeZCa7kqzmWXzGUanzpeD4E5qxtfsfvOiNp
gR0V4QJvbHDWInp0rM9+hfiaMm1Dkq2MmH/VcBGSe/0wf40ZPyVMrBtKUGn9BH9m
6BjiatPZsGV8c2soLy/7bMQu5+AmTbWvrP9Ifrq7LUJYQAra9540CyidJawyHDJJ
m+OITrOzMnPG9zeOgP49HFxKXtG0Sw0agJ9eg8uBz38e/aMdRgZgjCf9/+iVwdJP
9wMO6VTp/Rfqiur501aynO1dd1yMA7+H1t3UyQEKZwpPyR74G7WoffkGLOOYjud/
P1nhr9PVEzUtNMJZ/zE9BjFwUdVz8G/WJBzEAJeX7VvFWJ+zRsw9X1Bgd++QdZAD
tQsJUJVaiLIKldNTa6wmHETik83hGGNQ3524FvmTAOUi7R7UjL4NcjdXzL0J3FZR
Nfrzcho6INKpaDyR0+6bPTFYuzHWSimvfvTtOMfG3ErDpnXvX22DKXJQcJKi+lT1
BuCNKeMLvWr41miKpfQgVGa/zzRbR2Cf/8hJT4WT3HqNATGuDtGiyBc+DiYmSL76
H+G3k9HD9VpVsovUXydUwMJXP0Fy/AC05Wm53oZPg315nSV2pJa113IHKqiJNVYR
sttESMoD/K2tnyV/OVczcjue5qBErMIAPBuKbfLvaw+J15kmCZ8ig1ZKgxeKoNSb
hri/Gv6LdZVhYjfi7L3p/ebTMHCjQM0s5fgVnr4yRgrNcX4l5Z/R6ZdEH2s9nOME
VyYMYxV7icOYbdqX7BAIwuwgPySJYmFbnwkh+t+fuTAgNXeimaQTu4Yriq/Kgt6h
9XjflEXd/wvoqcM/LGaPmyq8VqtrE8qiZsq+S8gK3kE4H4m/jEkT/Qlh/B/5K6nC
9+r3LNqcrBEX6Ed4+JQuelIprgNUZF/lQNU8O/djKEQrP6gTSblMV1ovosw3hBqz
hHNxjEh5X00LDUzltuopeIBUGWKYsQMOYP6fC3XyTz7mO6FfWQeA5ZVOOh8gHbLx
i2+oDt22KtdsQrjkLVMshMf97tCxNucSkncY4xwiCfftz6j0Jkkek4+ZxUsZGcVH
k82Xfj8EyyXp4ZlhNE5TAFsaeWFPHij4Vh3Vz9CC0Mr6tEsuAy5jix6HYmIVKa3g
6gtat07ec6AVItqeo3c1cKRteo6clBq+PW9U6bSpY8Yw17G3g1DsLD9/J9JZRiT6
VDx18m/W2/E0S1ysu7FdV7JrgBPM/gqZHdwcRx1CpMAuyPUmYwE1j7WXqATXxHSJ
EtCA5uL2v6cLbYh9/KYGWZZ3Bp9VJg6kKotDAP+4NtklmAYyyK+AczNRppGjZZcH
sFsKKlBDYYKpsGr5QyacIJvFMA6jsm2tUXWKyRvlA+yMsh9G/j5R9ubCRSzpiK+v
MHxy9GGarMlYTWNmEdObZvPaYDWSTgU75NZWMGo86RlReDUJCtmVZbrtjciB2NxP
IIoKoA7RMef0/Y7/I2415DikWS3RCeYFS9kv32wwG9+hHwZesqZAkhnnqZof6Ael
60AI3zJYhepswNkcZLaRhBoTRjkoprSsBFwx872Rq7lDnheIExLfMhKYsg3btfO5
/Fv2i8wzLnUU/6G9LJ+8+cPK5A2fwMTB+gtKHXh7GkLKOxO2FHX7ypH8pqFbhZbA
NAB7zG0PtFAiYxTwkhb7wV4BlJzGAgsUkM9dSLoPQUCJ07xmDBtMJ0CFnFX0SRTh
haXLqMRcsi7pW8gsBckYamsBcuEgwk8NmZwga3NffcfgRSZrHJIxv+RjOj+w6/PW
iD5yFyyArLxnrA3WV8+46BM85EPFLNZPi8Q2w7Swn+BDrBrVB5fTb/I3y+7XIlCP
JTF0csbKQ9Ycnn21sRup9lE7KjvLN1SY5THSXZPFIgKqn3ipmjW4V0z8vLIgZprW
TuFE3w1hgc6iUN1KxfDcKpDVfgtUFjZhWAIHUJ9YB+fg7vMRv82sfr/PYb62QgX6
+XdRDJnSd04YQ5YwVndCjRrTq5rn2k8xUU5B6g7WLS2o92lOJdAIYp9b+/BbP0Mv
hNLxjB1s7rHkFfUvqMkLeo2PBDbl18jPNqyeAwzJh0n1nyDKhjONJNefwJOrIydy
zkYN9Pu5ZKEZa/VqqcUeF9REzTFpSbPEwriz3tgXeT1MwT+uJpsklWV7IoxWTX+N
GvcI7R9Ia/2Q+HJ6bcSHwtwMLg1O/QQCnqt+44pQXKS0vB3y/VjZSszp7I8iO+M4
GREtO6BSIJFAbU28TbvCBC0szJaBBx4f4DJglUEonQPdl82ZQ745LG+bKs+sMXdi
OVNdiEX11Nvq31ifkcBLhGza237dDlJavh/zyhG3SJODCpRlCMeNuGA+ifggZwxv
fqWj+GmNk5E6anxJM08hgg85XdeBPTel156942p9ZxCVA78tUpgnmcW0kskxDtyV
oBX5D5G23RqbJn/JFpPRpwBMWSMKmwqQpQ8+bh9HP4rY1Ev/5YYaoDNbKjTj/lju
MEIKuWux8qL5DMb78kxySoJ1ggdg76l83fzREuRFGZR+AAHzPe6uL3Z62Kj2Npm9
4qzkFP61ck/jdH10bM4ud9cCmxzxdgdXATNjmYQHpYDXAdZJzff5r86Slz9ublL7
hzXLXwLFAY1F8i3fKs1FdrDtV+pwJu4BgNcDGXYMqpnJowT/liUNXDSnj5zaOFLy
xQt3hAFm4EDJVRhhgwrnTEsViHL2r+KgAnHdnt2fK3+hDrR9h8D31uWDKa39m/oy
LRI3j5srwG09EdmseUQV0pIkjIKG9znpXG1EOEILg1UTr9+YQgafdFmDJNMR+Lja
mXDc/zp7f7sPFhrpfGcSkwpb0tdSQojddgOjoEq+9V1YYRj8fI1pOevzermWuMA9
f5323T0FBtg8KB6Mu+wOmABdOYanExlILqCfjlm+b2RE/oAFzgpBxRAwha8Pr2K/
XNNRhIP2GrluDzS4TwK1Yio/JVgZdBePWps0uNmQOKNQm8qGf9yI4nB3Yqa4tJzA
kzR4W1ldNSZge2lCalxbCSALRs+0idZ7jZ7xzhYIu0AbuY6XXSHNVhBqm1VVBDpu
PdQgKrB66UcOMGLr79Vf3/u3j31idGWDl3UMlUj7voGSNY9MeDvQnkTqOcWPV3F1
QPdt3HxDgUVlYIONqnaJn7GmzFrKxX3ohp5yi9gagdKxyhmJ7lYvrtuEb+H3P+Ti
GYG9u0xcGaAvGegYkwhW88YhtrQok0aSrOB+SVBXwpM6IQK2dfgBx6cY7vvBwgPE
0vCNAKASmc1wSRlI25Mcmtg8R3GWSK65Bjg73mpsEZ804cqt8rF/lGUpjBe8PhzW
Q8sFp5HbXPjbvH3lc9Nc3BOrckK/lrlnKkUSgEeSXBbvIoIqWx1PE1jCP9Wserqx
OISjK6VkHEq1dkRALiyTV/Y9qif7xUTopj2IhSSmL97PtqMvEaU3KnvWNa7z1a7C
lqcJtqf6MjrXD5ftMivqtCwoMgWf5ei+CVFCuHvMqS14yxL9fJLpqfdEw2YQSKDA
AxIPWoFL/dm/3yq2XCkt9eytEdi4BVTu5b7ENzFTz5S8luDOaFhqSz4x6ZB677Hs
VNda1MSW9gNW2Y/DhtRzQ8OkeV1+qBLHYI60VoQJTJaRAPWZzeEHeilshnQKrfp/
q1HR3cRQZqVPRt5O4zQMNhSsFUOCnzD1/BCsKqTvOYXxa20uxs18W52DrLG8BfNd
pin7TYkzIwMdkjIMJeFBQPjHQdldNVisUzfV2wU33S7KwY1rai48kzHNGjQ3zm8B
mMmxv7sliQzp50ZpwISuAGkcqWJrm6SExTKLdk/yIk9XBAMzCNqtHde4AiCbGriF
ZROR4dsJlxkUwCp4lmDBtO01iFqR7hkdVbHQoi1tGp3zxmoVw4jQUX351KU+kEb1
gpmr6ZgeDF2I6QCOIADtXZh+FU0hh2I21sziGtodMOH6McUpQp3IGW+WRORyXoR4
JO6k4PxZ7Eh8AJeFkpW09kWWw57V7AB3aISF33dInmJAIvN1vC+13u1OnVmALlSe
fJm63M0ywAdNImwyVNYMMZi3FxC6k5b/nc8FURVS074GV77E/PeCnbudAM9HPZwi
CjF5JwENBl3ycUH9uv18RvNvVuwqSz6Q1EhszR5kQO9sBQmed/roVtvG6SJTchI7
kchvUdeDmQI4TT7+5YbEn23FqTzKfC6iGdHZCCkalNbOYVRxPnfQzsPiv4vLu2x7
w7uIM0EUCHaahzvHaYwvrOX32oIx2EW9dcIE/JIZbTXfA41OWANlSKdaazw1CYC+
8fJEsve/DDTj2Ct5VB9hP5kZOv4NDXzNH4t76FT2fnj8u0u8IDSoKUZqpMSkVPpB
LhG+EA4Vc9sXuZA+OYMqmznVUD9Zm+fhoQrRt5WeRxceHAuv/uzt1eQWVacgmZV4
qO7JfWlRnSnZCDa3R1v0878j2gAmmJAa5jggkhhL5KEORm9d7IXdUg4DUOfpbt7o
ce/WSxlKDbE0xii03teFELlwcq3k52LXAtL3LVqfucO24T71+cyZOX9VjDrSDEIJ
u1BTZ5MDEchwUc5LnJFtGD8yVSNQ+b0Ho03bwvqjEdvCjdnlx95muWgUK8TLWtuQ
bRq9FVdDT8Cl/Kpd7S6DHXLLLmZByRh0ANSQUW1Pn8PK7yQyd5l6KvGSvWB6IgfP
pPwcbjKuS9qPIRC/zwKKP1OYdGwqjaP74w3ykpLdbm0npBUoqDIuFkjxWYtovs95
w0/ybNEnCoWrRKnMYwl14/2/jHtqVTDpqjfsC85rv8ylh4AzLEJkh9d4fIeI2eGw
LJiz+8jt0Y4DqNwBJFuObN7GaNNiQZb37iMv6U0/MN0ugQu2H1XzqVRLAscgiki5
U1Dk7uyg5O+AIfBza2xTqNNygqFxbrjE648iAWkj9dKqz+ALAjy5e3w4PztMzmDe
kcNDK2FYDfIM4oZL0pdDx/gKN70tl53V8ro/LShw5ZXDd6GA9YPT2U6F4ld/dqQx
xI9nf1jDSN5bQawXo1OX4fvdE0CYt1M3QaWdMHLo/I/20+KmsP/rwso7TDP6rRMe
QQ6H8ePnTIj8mikWeWXlFtNa0yit49WN+LUIm1RNM1tw3pClcuRyVmfIjwl9JHjp
AkELJIVLViY/HtmqQFGKBE06z0JI+9/KjjS+amMlTRu27q17VjjpVC06ktVlgeKy
u5bonp2S84ptjiDfOp6+CU63AJUamMmcmD06GaXigaBqv8C7dUDEvsH3BrvFOMbZ
YNX+kVCRs50uJ9o3duHeHs+OiWJLAb1lCd/8Vs4D2A3Lz1e1NCV0yu1QzLslELZN
nrhPh/t3Mh4GeD569GnogVHhlUXDoeQ8CcDRxBIbxbUHeANyvfbZ0norzq8/3Ro6
889RzBPusmJQvZ/w5ClgImP9wcECM5kHWae4aQQff1wiFXZuZ+SzSGrk76wJvwIL
TdErarSrdNrSDoIWqDCsWzvRrqwywuo6XPiPKf9+yEcNQqh3um+3eGvrTgTQt+Wx
XByCgw9w1pFGszB55rxBnlwM8DEPX2Mn8WJ0Ow9zueeyM918Bba3XnK0NyEWpxTV
k8lLf/TtQMmYlaFRnzl/4qEs/XVvrS1+rezoSlxXvnDHQWQSrFE9yOaowvXK8LCG
JAYp9eZTTVzqiGYIPkpJe0i7yeEhWE0no8mdfsFVl+8QmB6E0nDKiGkODSMCBea8
PlNu4FSwNHYRuiC98byKu3vD5N3qw/dbppYCYXSAkZfndt5xdkkGDEy/lyUy4Tq2
83e3rbPlpfXaG0F8MUXMm/ruPHUUYBs9/U9SY5TzU/KAOLUpTGAFck5BctyPiztb
v5qUKSo8N4M9391CyxiCnEjIMz9UV7RXJTsHJnyazuskO9Sa7EY6F043fTyg5N4X
DDeUI43gmfGrWMRNlVJb6aioH3i1PAeT20qXRQlGl4nSM9YXKX1tV+geBtNDp6s5
f0JUtLW0eHLjIRw2uxQa6Hlicd7Ch6FiOE5boT0h7dkZuzKvEe+CYjiGF/MciGca
h+4MAhHFxX8Y8ihF7/fExsaqU7Blj4HApJnvdT/m1PpV4esKRBbAtlX+3ANSE+Jj
BGZMB2HAkEc4s4dlsLzYTRduTfT9vOMwnS6+T69bJeHuLDXlklGedT7/E4VFzpkM
LZta690C37gGiX0dR6dBjqTaTuAjU8TiXn7TS+8/KY7KAOn71jwBf0VBXoHERNL3
rXPIDSgvBa8zdalcVaQyfMUxD2oGGDqKhZvD7D1sT7iRA+agzQyZmMk9r4JSYvPX
CPT8EdUQkbcNwGxhBgxpz7bufjAA5YzpDk2hH27Oo4r21G0NEimc04g7DUgLHNyS
MPCs0S3xmBbKhqsxwlzNk+9o67cAUkKBM/uQ+xqd8zdXHxW/tJdB+l6AWBDadKKj
/rUwXXHmwXxOrH+v0XVJtb/DMIz2LV/KaFHs95EysV3xo96oayTqJkDoTHNmUqAj
e/rsxsb2DbsJIidLz/BYCT1mMTsIsKtS4ZQkfRmTfsB7Lxu11Xu/Va4s4IQku+Iu
5Yqxav1ZkyoQo2FYUS255xR+X7QW9NkxCZEPmqBV4lRsgVF41NXY76qamgJhR0cE
NgG/g6qROl3/zWmXDZwFGlwM/zgm8KDMoKOGR3rb1g1EuBBn3bk/uAIBvpdEzcLl
D/Oxj8am64VCgnDnI6IsUxkMd8uMNpy3PtqCNcINDDqcKfaAAcn3vSiqNejhCm8O
h4BYoRewU6Nic4L9eZy76vapAd8SQDjJvv+yy8BnM6cVxWECYm/GysOcKOzQTca+
LQqfn91dyx1eJu4JODtzUkhYMsddQ551cBFlf8tIP4Dmg23kZidxOBtB7FzjP26s
nOPxx2o82BuX9sHLc2VTXAadysteHVb64U//vE+cf8HEBF9KQDSfk66QM5z8ROCH
cy61kKUMQJdMZamkPivnaravpNRZC5NZ4k8xFOjxw/jzSipWQPvI/+fy+ckAt2WH
JHmO3TikRupTwmMp2BLweohkasANnJ3zt3KMZbn7QgDaHiWTklVmRHYO7d0WT6uZ
FRWkEcs50UD6CK6FHEJo9zi3HKzX9iSusiIhexQ7VvJWV+T3BMW17nN7pq2ZeZ5U
qNlVindFrCYpwmJsGPRwqls6AgpKOBJf57Z6Bq2E4wjIAyVphQmbRXgWlxVpPUyG
2yhJcRJyV+21UswAXaKoeHXDuOqlhapkPfEjg3wms71c1WyMYh0NTzNCP8deddX3
QYHE6H+5w357qqADZo1W+I08AqUXuTf/I0N9r71Pj/BSspnT4jq1onZsXX5Xab+H
hmFqK5TDFuq4VEZoymYBafTTzjulc+/TYgROmM+N3FS20cjt8FhtYXE9irlbhSu6
bUNfCJg3hkeoyBInxPSO4Slq5kwmxGSr40ob3MZnqvHsw3tkDYz4Q1CHLl8BaoHe
P6tb4jf7q+FwY32uJ51JCvYZkm0y7CbxgPufq82vSc5obCqVDYyskJun1ITOTvrb
7kgTjDqcLDgXyp1e5exHFGcyYBCcq8eIktuRTTayfR9H7gYxC+YB8mgHmTSMfjFx
5KQGlsjB3ZvFQFkh0qNaWKOiHBHp71iUPt6YZjH5eukXcdEfeBdigoSpEMH3w3+w
hw9GDgDcXQ3kD3StzGa272yZxCEjGOE741qSFqe/pXc2AAM9wpfS2JeZj1k1uOPb
EyrOj9XGOj+3+Hdx92HEzei9io2QP5yVxSD0k5wC5nmd8U9JXQBnLhki9eTHDj/v
EvRr29bMGdflAHaaEXWwXzYxBQ2Kw0OamulAeEP+z8zm/KTv5jvR26LSvXg/IHyM
nWtfeonliaA7rMzOBJq8pe4DtiG3DUyKZEArjwy8sJlsX4R9DfVccNDjZ/UlInoB
z4TM3avOtN227iEp+WQLNHDd1kY6+3Bi6xpuBJCZiLXFYVw6gYziMamCEqJv0cYc
5Mvta6q/+qqyA84cLRlmRRuqWgZX5h45ItfZBxJylfiZMBc1vxuGuVARwWYZB6vH
cFQgbqcRemxKZx6bcpHHXNSVJgaUEHWk2BkM7KR7FYDbwfxTlv7by/mxY2/bDqAp
c5Z6Pgi4Oq2EuLndY7hPh2KL1eV5l4otX+lO8mshddN+KGwKUIF7FIplw5x6AWCH
s52WX+VHE8nKa81td8i6u7/z+X5WRD20De4H8haB5WcxVWNqWVyjJ7QkYelQn1TQ
NYOOvuAflZTFxyoQqSLdFNjokefUKdagi1FlRk9nlWolkD9Ei46boD9zuu5WW5Mt
pEQYK7lLDtuAaYxxyn12l9+tcgCX0ZVHXA5Dl91Ovkn+GbP5Lo3avCaXT6DQJg4p
0Y6Ukhp4Ple/I5RwxUXp7S9a2TAi8ogsq0OSxdvoF+vDYx1nfkX9vbfSilkNNwh7
YtjIP6ERSZMzml/5aWRQaofHfvfY30o0pW1zb+Rj4UIyhRonvBUp9jZ51N0wRa8H
uhCE5XDCTlBq5LR/hyl4DFE+vMn9+vLfGAYiOdOF3GfRR4HLb9pifpVC5ddqG83A
brjHZHMszQn2lgVk2ZoTV9jVzg8HohP51UKV1j1QHvxG/3KDmlVUnqVPsdCqrZoF
BPTRhPuJPwaQCyD2jqNkui1hXSClCREV0Mst8i0QbCqdreQl9iY5t0X/W8EnU8Qw
lxL4a8gPsA5LngbEVFuIw7YG9LauGVsgqFRZBXEddZSX5Jd6QCEzcDmTyiWe0lX4
3Atu9DDEgMbXFtVcGCraZYjPiAm2JpKpGH3ZesQzm9iTICdGhxpdYG1sDFLMkqFS
B25ANAcarXYX2AWOy22uvjJgnWvIqr1rz7tVyOwFB8JMDTT3L1ss5onIqt/iarT5
E9H0M8L3Byq1WwaCIJiaSH1xIvhdfuzSrWgN4BUKqc4BjhaparX2p9ngXDbS6Kdk
6WGzU6LNyfsela8b43mQYTsLm8ngXVuamhp95uAR9bfBDOVMC2p05v/9jdlFqd55
9UnWSD0aM4xw418Y530WbZjIRNMeyT92FEl5D5ferJvtilrwgwhIxamAHqQkbKnI
e5oyQOs0r2EghXJIHTXo6r6esLwQJq22H017Ll9MM1Vy+HuvRlZH6QfTagzQRml0
enlQ9PXhKKhFi9yXIv6f1pB9ElON0NLUYQyPOmRkfPH0tb0Z/WGzEY2hV07kjPsi
B70q9ZWU14PLvls20W9k87PhfBXqh/WgyatD4cezhqM0d6rrkXgLgPE6XbZkpWpp
WE4VGCeZxEQw2lhCxICk9naQnO9UbAY7cVYzX4SDLA5zfMks/LGLR8JM10g7y4vl
VOuvEqhoU87e2rPMJA1NMsFJDnKNtrrJlooM/tq7dc1zl6+k1NpUfOaMye40jXrW
WRxbWPaO+tsYYX+5/2ewGHToH09y3nPDTaHGL2KLxbSbQ+6Dg+b79BtOoN7SV8x9
eGe5nJ99rCs4T+270RpfftfrmNWQoPb3c1m2HMvQiiBdXy0vAEkMqePt8qPP/8V/
crVKYSM+Pn8xVdJRO/unieWGLxkofan5dhtmBrD1DeNpxuwMY+K0d4KumisKW8Ox
srurgNCDxdhOTdRO+fmxHUdXl2oz2SRUQKlSHvJfr89KJ8SQP+rsugRn9ebTlXdm
/kGfp2YedkgG7RHQeWJlh4MQNGskbpcqENKYJUAirwHuYAQBmEqpyVrbJofh8djM
QJuKjIuG72a65fm9sY1VrNC2mBcd9umFN/VYgNbxkJFt4Cf7ZsNNDOxqYqfgWnIw
B3ZRuH/CWqtXZ2fiqZxDBgxaa8PdE3Wrygq1P/oOBhQubmC0he94AssKYLUIYPil
NGPI6/ci/9JJDOkxlYUWKMC0hBoZqTincxGzAGPAFXaqDYPQrHQ1dT13CG13bjJq
575bcnFDh2saYLqDBZh28+Wj3DlYz/PVf43V5ezdyNsTlkAn8Io9rl3/WlWHfdXW
GG82CHVuy1woX0lNgtnWW2NnrYi1/v3sc9WZNPWZOqqBvidGNdd9S8wJkehC+Yzs
HsWi2LBYtpKAtWSGyGHfNJhFM4YIfxYZZnAhD4oPUZ6ewzTxnJEYIybcXyWjJEFu
rAAt+EGlFULh6FXC91Zz2zh9ywtpmyBTxpX7zwLbY4RHPefKe4UOPPoo9xRylp7t
fBBKVNJ4GVKtl8jumU96foihNPj5+rnkuhx/Q9e4lWdw+wBPXvT5TXAxFQgddTqv
cON2VE/b7JI9gNI5nQmtindrnkaDWsxkPjPYn03N6C3PV1h84i592448DIhjCIKW
5r23HIQtU69XDkxHcrjHJQg8t0FryK/wYDK/NddzMgOmQCSImbYidZ5XVBOAfE0C
6XTGVZPS5CCj1SYiEfyGY+X+5H/rpWzcDMW16ouKUay316/a7KOb9oOKTzVvrFxZ
rZ63rjuxkPTZqCrKlu+q47V91sau2Vd8e6Es0lmvNYP7nJ1l5p/CPqcv7lyrPqlv
/0rMdx7Z1/g3QIIE2wncQwO0BtMNNMAkfg2ns53tY+tEZ7opowXfppLsbO9mnlxH
CdbqvO6v/2Bb9nXZ6Qz11JRe3wUbN6kFj5Dw+lGYecVQ5CvEKYTVWOdpQSZY790R
wgUfprfmGH1ZlMTP0hr3CoULQdPdCWfzObgDZbUCFomqyXRR7ObUUEiaa1pjpxPD
pimaEZV591DEFbL/eDyVdkO61413i3erpj6S4Q9dMIR/M4q7/aMwQMwHIFhNp39J
PyTZa9wLvTABKDvN6m1hNe0JGWnN6qeK6LS3++6wwDhZcyZnyc1+tfboYID2GqyZ
Mz/0Zmpf805P86sA28km+k4hDLMXwEnmrLPDCKrblo5ljyuPWZ/COIgw8WOl0jE7
0addKYKkdyIHQby17sU8nRUqXRChdhqcfSQgRP5Oj84ylY8QyidJUflh3CngNnNZ
a6GaZMUdsIxoNk9q2+O2KG1gfSlqt2t4lnQr4tT/0GZO4/LWrBSba4GLeEci2Ojw
sRuGabOC2mjl4G66gJh5PqVtG6x7jByqCMug82jxxZEd3hFrPstJwyKHPRXv0RmL
3a1K4+MyqHjK7bUcK1RS8onRDlSiHlkPGu60Zu0KHjAVhcbYzK4fgCiq9cmOTC9W
z584A6GntpiJ9Feh2F/rrewR/woOQSo9ETXz1kOPA7YikFL10uj29OCdXcjzjqdW
9MNlwPCsvRGKiLFvwzXSsX7lO+2riRWMKZF9bTpRYN/fhHR+66RP5C5KI6tM6Yrx
0IroMQgRiHrd7dK/PV57Ws7TkcubSOT7UHwcwYcVz0M+aVQv/utJNHA/HI5jRHCt
hNJglL4tU4C1q24+hMW7zx8xCaeb6Qd/lZjQI4FeHi8WDmWsAnvG1U0GSd7/yUyI
4bE5owzh5615qwQxiHc2p5lKMKeuhJG0GRAM7V7klpY7et8f98a3WkwpvT+aS4Hl
s3cZ31wQLirWF+0gBW2QR1kNRySabmpxy3zNWixvgCY+NL/EU2MXHlSY47j9Y/Ki
5sKPCqdOAX5rEIJ3fpPKJ8hM+YZ2ayyBlpaONC0a4wFOkeQ0nCYzKuU3xz58rg+4
C35rlGNlDruW8XJcN+bTAxgD5Mwe78/K+A5eGJqJgU0IDk5VPtqBEHnbGETOENsh
pI7KNO1YhDHVi2+p6T+17zJcZl6UCJIBZIneeKMGOqbF04FF6gtYDfM4nPwzFVpG
D0BsdO+QwNYoOeuVwg0I6OQ29uFUgo6xwHZTEDX1jQHUk18uV+PFCsKXEa+eMpPh
gGfubv1obLBs7Q2mtSCfb3c9GjlUATKSqZK6DVcqrQB0IfTlVHj5Jg5ttkCMbcYd
iXNPk+O3jjPOkqKXO9VQbLw/NQYUhusBf2POZgpCBGsGnwq87MfOkDZn8I/sWMJf
Wn9sg+/4sijEStVYm6Da7ieB1UuWStRQvOU3iIs/c/1pW1OQVOMvq3T+27PggZ9N
wHzZ+C7n4HzZLvzSW/XI/aHuaUic1yVov0YG1yl0K68g/2XSngv8zXdDMSf0lxWs
v2zWAfXJ0/DnM4Xg1XxNvwa/lZ/9953uwV283FeXbogNskaIzng7IqhCwTtovpc2
9RlxOoeiXfvtZkcyFTcpVgFgVhEXtVNRTjwKStdBAy6O+Htzg+xzzPaXs40Fxgoi
s8iDcuPosza7Kpx0FbGh4EOwXN6KmTARzaXMYrokhXoIWZFi15rsDGjlA22qEhSY
rYSTddCCHoKXB+JtRlgxn/RgdY2iZ4fJwY8J0/b9MGyMZyt+c0nWDAslDiRWIEvu
a3Fk9QqEgxSsZo0aMZ0K2xRFAJpv/cIW2He1+K+qpdvNWCAZ4rS+Cgg7oKQaVKXt
MTZy3paYRGQKa1A4yAoPlo2zesa+hqFCs2O22i/MOwGH6t7hRjiU/UrdKjfpDKyu
OzVgeCUdX2L49Cc1hTxnx/pKxL8I1lAqh0XU/WJOU2RU5Oi7g8O+L1AUSw4QR2VC
UqnVDUDXUOr36RgLUiGaXAfklpMfNm6MXN46PQ5C66F4WxJBecAr2TlLjpII+kgd
++MIIon1gdEUcpcJLf/FxCuP1N4GBNLg50GCR6bs3/ACDr9hLSmkzkOPA89iD/dM
eD/0CMhHFSgJsvNneDI8OyLd3DNPL8GXCpQPa055qKL2E4sxe8HbZo4z1wiuIKJ8
OCWFE6BqofyN3NUF19wGk2NlXjvGBxOjFBfz/APIHrGi8vz8AaXEKMLMdW12ghZx
suql+rhNEMiUHAJaxyC+3ao8ZvRpeunu2MtjCJSVEYX+hxQT0edBkfch7DmCsByX
poVn+jQ1ud+yKXSAdymenJ8bozd+JpW7iQNsGAcW6qCWTda78Ikqdy0mQMdV7fla
3nV3mI8hgyjpf/flsOK1tduYCl7Pdml+KivMl81OBh4sleNv4/FK8b9D/G0Md+PK
jp0dkXgYZMpTgjEoZiwUlDM7wZO554PSULHemSK0ALQGHJsTtVKPXAR5zmbEWk47
AC3RKLc/zM1HcBv7r2KZ89LLQEzbtRSiC+bHUcrWKiRS/qHgGEUdcntvbakJvWFv
8/Bq2f8tCG2Cb64+pC9FR8052kJfrOc8iXs14qs7d3SjscyaKUGyi4/RHaEmx1EM
LCSIX3QZ9mrQshYpgVOX5Ibx5wy0GxC4B4ipSKgtAsz8Bd2WSTZpReG054Ra6Tdh
uQTRx7K21ExeWCVOo+FK2bL4tnZ04GR/vILf+6fHInYg0uiB+VmW48v462pnl5L0
+PNZjjgDMowkKNusVoy1Y2DRzpjI8TAsyiv9mvhq1mbwBGOx2+OMW4zS6SXi+vfh
f2Nf7+RiFMXX93/bNLGoUnIT1dQxKm6X8I+BmlCcPoAlGu/9ghBe7LNmlSlMjQy8
vz4Dorv+tamj9NGOmonCPRXO30pLsfvRLnlCCERwng9N5S/BWnRjPmc0Aajs3rVJ
oFdER2Ls+d469F44CH1/TdbxymEUhzzoQcKOtldnUy7z7L2t97gE77XNkIYN4LQW
ymoBrJHJxyARMTk1hXlHa+2MOvrbZf16vgrhsOxa5EclMeUz9bIAFkKU38tOUwRg
nAoLrLZ0Ahe0Wy/6nMktQ1AhclCZFyEdJ3nU6uKxvRBAL2SjS0u/fpkdIH10f+eA
CybhHo9N8bxWUuj2Szh16eWPSRuedlJBIGdmW8qUxHVCH2hg9+uTuisIUjQksZnW
8KiIFHgtnR8kkMhdRzzrUKf7EGEYThchc2PO6biPW3BRDZGzplH28VjC2UmHAZyG
jjWAvqsF+m+YMVqiwtwrEHQm7Lrf92B6F3KKEAE2mYuQbhzMUpmD8DTiKAAgCcJq
21g6fiay+Y6xoWC4pGCX7pAw0DPtKP08oaKjbgLVLuHzMszxncOSD5k4lAfqc+MC
DSh7oKUjLzes9MQuHBJQUQwviRzpfhxDmOCG9kwNVqwCCZfUA+f6LHFnwQSpedxN
lSB93WiDs8h0Eq3uYlC5B0xxPQceLqpH7xQ2TcSwM1XaXINWbWPFTgJvyJLBDjEi
zOaHGq2sGNtUlWDWZqUrpcE8tubJeFlQ1unt6b+JU4SETekcIwE1KyCIoViJ+hEo
rBwUJMy00k2Zdl1xHzRqVusWUidKV5uicweUhY9qcHeutqrvAMWCIyNhuxPuzdqd
S1AIBhdeVS6q+2Sa2Tsb5UQfyUZOkXhLPG78K/zg7Dz/AQauAdJRFFG+Y75oHpf+
UXqQETjLh2vmh80j+RUymW4iUj3NuYy9YEg2axM2bRUWEjzJYJrJTmuxTNaiUnWC
tj+NS8c09NnF2T4lJQUR6yPiySP91ifb3o5DCmVB5/O499bMvlL3RkLnfFOL4VSS
fusull2nrbBPHZxmDjDxBBe1aQFiZeWvEdSG7As6ICtAw2BuENBVqT6EwHHWhcqF
J+5ifsGg2YvSsgk3IuKAcZgt1tspucGK1xIOhV8REMU1VY/SnVEgD1mZMwGhhYNy
RqTWpDX/En3x5h8bPl8kFae2J0xTyh8doLqGu/E8AQ0EUx55eSWaI8SzBpdfbw4a
5o9FaaFfWfps3VYjmHw+UCRwcPJx68byyBbACjdgYzKWFY6/EShspyi+LJXFX5d2
UH9COnqN6uktoIEuceFxcFcM5gEV2RNAxloOn1rYvYGORh+GjHpqHMt3JQMQNZot
uJqDzDlVDWdi9TmHb7TUji7l3ETvJqY364qAvYSeHXVyc12lkI0RDNDCXmoGLDe0
7bZ9lM2hFWgUWaK7PUDAMl3/3tgwI3RuQxWgbUpKdi4tnH7CnL75k+YNqs94Hne0
u4aEo0wFo3nFa84nilYMqsquMou6d64JBBUf8qdo/BCCh+hLvBLMCTImf4UxjkwP
njGKCwDEfcC8ksTDpmJ4lTjNLUD4QghDqWppL/GlwX3O987YVSosXJXfkcySpHco
DwGVGVXobJBQgTLubaHxvA4xq0bgTri8u0O6A/G8+9uc1/05QYinZlJ3h5+h9S6F
w+JYlpU26MPpIwujTpSzmepKxQqCnbZSatwruvAPGkIsDzlOAaXna2dtCo7Jub6a
I9F4JXMnQ8P1IlL7a8j+NOBMx06TRB9pNzTKl7eH8fOsPkGsSurfrRLvYivrVgV1
c48s/cyW/jTcBAFP2kkX1/OY5aNb9en1JfVrlj6YIU18jnUOvt112NZ4AT4EWOy4
+lo6CllHS1IlHIduB7mCHg6q4ySA01qCDd50bLoOfFzf0Kb8V/h1YUoi1pgoyF3Q
8KVdjTSj1LyAlrHcIYNPFkNJbjowWdyTYPa5prWg2CGlBgAkEodW7fP3aO7UqiXS
EmKEziW3Z/u8MVTiJsF5HmqheFAuDDOa5hg22Yb2QOmTNlEfKCIwDwScHuLjAqsI
YLTfsaybkM+fdoRG2WSd0ySzSTsxlA8tHL7mcNJc02lSCvVxIR/HCboM6pqKm4P/
Bij+xzoj/SJeouXTuew/ugplgnHc3cbEYH0fTNrCWJn6Z3M416QQkpdAbkIbmQen
rfcuMzxdPHBhJ4omZc9ci+G+nYOUnzqgCzCegmwhfNzYlnYYSd287RcDRQQBXfYT
dx3tJfvNtn1sFEBIvWjWP0jfaCi+hZSMvJwNBy2nmggh0ZNhRu8J40U0BQ9JHcTf
Q0b+FGOdgSoDWc/mEFvh5fJJ1gO/eyQa711KhC0rlJyRcJr2Nciyds538C4+QnQS
t8gmm/XlcQk5wztyWix3ZNWGd+CfKuHiDn9d0+IE4wa6rATTVEtzb9jpL5rg+Df0
WJog7v/tgyDfjaFWgxHGXvcXGBIvhUvRjAqvWsmdAV4GjszwagctyG8b5Iby1TVI
/e+bC2/k4CvA/vWyQqmyGMtxn6aqetO4H/udmYpK5AZavPqCM0RuJ8YWIxeP6xeU
ykbO+iqxyyd5aQhF6TYnr9s8IpsUjG19JaJvXxWkb/wkd+MTELd8xo8H3HdQAUWc
iUJbeLBxAllN/hEtaNEoqzE/ZluxUV84/HanDm1MOpLPC+pZemTZaDWRjt5a9XRS
IbYw3Gwq/ar81SpTw3TPGS4MNowCwDDmeQmCOKzLEWo7zdJddajFB9bjUvHtcsMs
h9YGRMhAjUvvdySxcqR1OA5IX9TF3XyxMtW4hZNxzYNGUwDx9T+89KCtk8gf7yqG
SUWYiJ0TJUzUqwYHw3bZviDMBj5uQIbT9U9pHkfK+c6SBoFmM6KEPcjsRFgC4pT4
XSqGRXjfjaYDj4ypG9DNxT+3BcMYDuuSEJt8cihIgrDADORaYu/FRoiiOHjle03V
OInJikHnBZNLHa/N/R3sB9DSYnkavPUQ8TUGYH+35Zidnf7/DdqkJqysrE01Al/P
FN+IytQIrHfwIoHP+BDGYkeeeQCXwPK9Ku/k73tGt1TdzhzB9tOfUxXteEZRhWBm
aW+8FtvVqdtNoepswubas4mkbMDF9I/C56F68nyJyrdlYqd1X/nLY9pR+LspVYv5
g8P0A5mg8f+IPfpiu6yFQsx2peS6oJ+TipbnKzsPx96fv5k0XdqJkUBMqbR5Bbux
+2xeDb+Vbl3MWBUL5ECWUKs7eenJqqv+w0Qjvx4lgLXPnqHZI7MFw1eHu3FY0HjK
w/EGKW8rzxBSMwl2D4IRXEMJNnxRR5HcyrabfUagkq45ZwDVBx31JrOEClt54VPR
wKAlBKoGb0pvTFDCm/L1Iq62Zn12YACiuDQcExbJXU0Wq2QTpEZOUDg+wyev+xVE
tffndPsDvd70oOcu2XvOS2vDF/ImGm0bdMCU3tiMWlJUsonqiPr+kT/VCoxoW5cP
5SZoyQn/d5F/O2wkyXQjyapqegwEglp8kF7PRfDb+CeCrCa+/NeAvSjpRvAxRmij
eTu09yhzQFDsuyxcmCEdC4xg+q25ZdTPWcmbwxCOnVFajQfeAu1uNdHhMzNXjvs/
SbA1daOsNmw+AqdK88VNiMja34woJO4UXnHMGoLXIU2/AxVYGIXyGevGXDpt56m2
s7mOR2y/APHaYSFG5/O70wJP8/98tvm2xN2Bp5mc+K+/REPq+fPGIU25XaforKlP
7V7r9AF20+iP/00uDaJ0dG++LhdkXhjs9E0+CB/OxLownNk8azIdEAZaz8/UiJh2
CIu35lf4C+hSNO2eL++mnpmPUZ3EBsedxhY1cYoy9JY5T4XkjG0h0HXwbfr3uyOQ
3zqTsEopyB9LGjEdwLnrLgXwSa02C+s0KCUJyblfWt0ITWqH5SsZ7Edfiurrobll
VYlTDCpysfRp8SMstEXxsr8Zvv1DmlPWMnT1p5CPryR6GjnuwwYrkIuL54hVJB1X
MSpV1SNboJi2XR7GJNysdBri+n4pf4ODga5eJo9rLZsSLokeA6pcusaj3DWLkLe1
PahI3EGDcd6FWDfy6oNwf3+D6WAZa6Np5Sr6xRzLMDvydwKhQ1YtnfUIf2WkSo/4
/exeQLiPcRAMj6WznnFBI4YbAkHy+3qvxqncSFKOCXOP+ObJHkIeWXsdv4mlBygY
ZsVlcFujBtveevIS2jO/uDmJ4Amy7LKIrghfc3ohD89NcU+tRDU6OF5k/tgn3LVX
Sz4tK8KUerEaw7gzFzFprSGyXZy/tpbh1+qpEjvB1Fw8m7iZ6H7QvozRXn3UjeOg
ALLZg3CDP3Dwilc8DCwyYfa+ft4xUrNB/a+mP+0LziBLg9Wm6DH8qEQXk0tO6IKW
cFyB5kt0LeWlw1eX/GCu5eOu5Z6irA2ZoHwAJQA2y/0VREM/8KDvPCwqy0qAb0wa
tZq8sj6c2+r6QGmMDRqKJG4WsCeS2jZSan9j+Ctezr1eROkUkmDzDxc93UydFN+Q
I/0j3yx53OWypL28jB5KldR+8j2QKOIc0qHgx73UyyMuiv17l6i+sxx3blvRS4+G
5UNaTvA+J9/U+91M1ehdhHXlYvo2vIeregdxvqykkXm7niMItqS+U7Z1/Ag9hajO
7XOamFZzT0tGo7U0wogCrtkRVfTfnjh0umKofItrMFlqV+VzJi8Z+DnxrDqop1LG
nJR39JWYS4u4+wZBpcmfEXW99xhk8QumKXXcZUR97Xz05usT3cwKuOVQLsbSYpXp
tUQXDW+5GQe2w81z/iFi189pkl4IH1J6QNytlFvBYJUXz2NHO2wafCbK/bqCV2qD
u5FVs3WM5C+V0h19PTVqNdvxJb3RsJPVpKn+HbNr/naAbd/XIPSr260ph2Fg6ChU
cAQVD7ZHb2tbPzIqC1tt6GLN1rZEOvdNfSRNuKrqyrF5/YHulmAznp+XTauG2niD
1jqgkSIxeUaNl9HXTD3Q3965eIU/b1kHOnZ24xaIX7lnV7eELMwW8NcwZl5+WSw4
lNRGZJKbLG3SNp+C4Celzv4PGigTxC/xt3oN8+MJLgF5D4XdQKyccuv2QGK7G9o1
JpBYrToK30tyKYR9i20fgl1dAJOpO5YwQ9Q8fzpgcoFjYz5Z0HKDHOFdZ8OWt+6o
EaOq/hIjNcn/lFnP0LF4yxmrdyecoSYIsltEYMqGZp4XJ90qFnEK+PU7dsYo5FHm
FuDrEfnvgM+jDhcWSaA5ghqId3XX3ytCQEnKCzoOqkn8oAwQ+DyibuHIFEuKxvjy
ff0547+ROK/7kTxBD/Kp8a1tz58UMMAjC8B5qLTbjoSKGGYzQWy8RP8pLHbVzlbP
m8lRyxoWRCuRJdLAatIx9+u0w5On59NEXQ45mxKsr+jLyQQCJpThcwHLU4DlRy7U
ckMYWQrj314fc3+4e/66OZ2cdH+RuE4BwAzO/2nuZykdHC7z/2JS3LfKKV60tREp
McBTZELOjkVWk/1RLzNKfNwFZ7Ldl32QeWl61RxQki6XyA2zUu0jhuNMT+/5fnb6
z/gb2WgfueV9V7ylxVfPKvyziT4qghSngpb/qjHmV/VJqMS+qneSZRQIoE65oeIF
c6Nh4uwdsglYVguzap1Lxpp/4gxmHyYSM5iXF2wRXmNfDGceWSGdFhfXvioG6Mjs
VIfHFycWgb8whxfd19ACiY2yLIm5GZq8XLC6j2euDdpCbctONWQ4NMKa3noej73Z
j3CTDGa8/h8J9lbS8dBkNLm/wugG4PpP053YAUH99Vk6BztKl9+apuzqBPwUmun1
H/oEMl2Ik2lHKQsJHFgSFdhm4ffSd6Fh3xbl82AgcbQow1G6bmDHAnVF21M8spk+
XhZ6nx5cjmaUQ0RZ0Ptu4apzUxrdPK3VmJKIwoJeEepQTgSi3VAC4OgtncfyX7YL
COR92CMwNZjoUyCCTTbW6A94hWn60kG//jEdbupJMZXkavDTsp/lGq5nZyJcn9D3
gU+Z0pet6qsuifLkKGITR1XWKrbHVHAhz5HUvbNOMcmZHtbtj5PZBnqNo5wO5z8q
S72sur97uLYbXSNXiXhFM1kZJ+cnYcObYIFhabLry2jmHWIdo0FWgGE5G5X8qDKa
dd2aEHYwA/Y/Jd+8gLO6s2Uu17uGw8LB43/1SwgZdgKvJ1hm/86/9F1oNADPP7aG
KB2VD/WXd59a4rbYcXjK/B3Ow3pac+avtUy7Ulm/hNGCN2FjbTBkFYmefXUljNDc
eDp8vp/B15NfP+niF4fHYx4P8OMlfBT+c/n6BQfXn+JANUt41ccj99Dlp/CzMrnf
1kDWV8BqT4olJBxy5ECiEOHQ6bVr2/QR/pii8WjAx205T3H2OUtffqN0IxRsJilz
WyvKQgvU3LTn0HxiVkwi/vOHJLgKSBHgcDSbc1YO5FGeOHQFOUtQdlORPi4M0a2D
yqDabJK7xJbl54PwnQtRoz31wS0xrCjgI799CdLx5IZmwkasr/lwDsAmteQfWS+S
OSBke/F0WEGn8ZJYdu2Oc/5YjXiGy4bfz6PGS8upK3DXlUCPLmdc55ZaIg8Z4Y99
4Qi7EzQEEY9c8OOi2P+BVeTQc9wAZL6n7jCOkMwlQB504O8ica025luHjoLmP57k
nJVfG1qcKwswoi4Ckhp3u2du3ftCyLXtj8Zid/xrlxFS7lVFzuyiKD7JwBXxvKpi
9Mb44p4wwmtty5v4fMhKGlAvknJ/G13w6J594CjCghrq9dqeE7rchmZB/sdmVrQR
GiVHjTZjrP/OWTLnhW1bkHIDSn+oZPVVksFwjwbNrhhGc9sSg9X8l4+pL3jxDo1j
DIdT8WaWWMDxdsZLry/wm7htP3LhJXBx6isHRlQx9cVqp/GsPsvxJqwuctnI/NI4
nePJDMlR8EwpC9YDi8hGrpyyNlpR3lmW0x8hfARxEQgbEmplcOb3FEA4tXpjZAWM
Ol4IDGPJy+BZkSQQT3Ekgn9xCwSPaENUxYIZCWIB6gFMAMRFQObM+RZaKjzXxdl9
bIGubRuDHLugENtnrq+V0oAfKaiTxutujWnMF68vvB+n1nltkvIWEYnr+YBoPnhc
JPK1AX5Q/l+W+ursrI612Nj5E+8uhvQxosWAZU2ASCzQuvawnCI1ItoDAMskDPTe
EdhLzMLk4+wfuv1eAZMLx9hdO36TVxgw4fFZe6XM2ER4/OW1Qjjx5uGkIwzz83y8
Sja2E/h2Bndn0WC82eAZ/2Nako2N1jMvJbb2N15KUQxUdqamXK6oVIhZ7TjJEwqb
jZmKRIKgtk5iWIoHwDHiSfH3+V9KEfz1IZtwNeAc94vnXJLf7fFLl1SpkLw0o0x8
56zQucYYwNnzUex8Tth4JhhaDSC9npiPdCmwoVrnb7v8tY+DMNer/Kj/ve5oYArZ
9ZIrWKjG0R5aznOY3i9ObgFVrC0b/VLgYwTE3CQQv9kv+Q+GUYBoZrmakM9iqCm1
dkNk8yXuC3mcCvq7/hE80la2z/BYWnq/CRrbJA3m4Cz3MiS5ZTDVpF/6H/puAMxO
NLuefT0xGR1w523gazOdGUMXvYaNfosF2TV3LiQhK6SgJRsJ3XhnYV27yndP7lsm
iVXImqCG+orpvFVVUHP5Bb+o3tKZGQh2X8iWquXiqtBSfe44/tM6VazBt+dmfjrn
UWdH069qTGgxp/XVusnRbjYlWFDmNiZ6ICVlql7IQlfGFaeqxru0YKZyXVKl6UOo
FAiAqwusqZrqRTrIbSly2H0QLh7ub7WTfln25mjlLkQg8Yd3XaEFdjrrtR86gpRb
kJqhrHvh66v5nDSzoLU6lg7YXoW5aO2xXrp+8YPAKA/Zk4U38WL2EGB+akFAAEJd
N58kOuQU4vshuIWeN/y5QmMOqYru4lCaJcvSirdS9azIRYKjrgHy8cTuKb4Oek1x
zGc20MGs90iRuKg6Ofoq+ocL12L1KDnc7Tf7YmSZct3PRdPad4Apvs3MKtv1Rs4u
IqAmG5MmiXrz4CIqMrH9BCYxr2COjI0DH9BcHnLmeEJkOvz2tsViZGnbaGjwrym9
U3lUEupMgRkeG4zK6T8csgfoPNXgroH+NKBa4D/cDZwY+4ZkBEQt5QVJr93DO7U2
ZPx0GsLbWcZWbMhBnHf9cPoFQFtUFj1vsU+ARfG6//0PAB9niwjdj8aTY47ceV6i
ISka8zDCS+Js36VDEXDTV7ExWGsAIGTsec/quRp1oDQ5jpgko3K5m1BTpZqXIhkN
1Oa//f7QvR0IwEzxn5dHZ5QS3qEpSt+KtEatL0lxgWsl7Q2ulGPRVGi7byzfCAqj
W089JbD4/CzIUqMXRv9Wctm5i8oGaQyFa0q0PXtjtwoiwXcjWM39BD7u1fthgqZK
5n2aNEpxEDP5f812rQ2Wv3nOWl8KEBHlEdH6nECT4aZUVg9odUpO2nnoEWs4M9a+
XMa5kJgS6C9BKa7TEoHUXD1zQZWL55GiM1nj+bQglRxSjgXLSr3ao/4YuXg60KU8
xUGDS6u06+lD0H5BsLlZ5Fc7renE1YaJdON5ZErztwdMU0HFl6O36B+RdKsmi9T8
3h+w/KyoC03q+bUkv7WHuoWjkp7Aj4EecaEgFFSWQkR/ZU/YFyT8Fc/jmw6ujlUB
m/Gd7BDrZ/zldpyB3GG6APXHCkKUSXlOklS3srL8Plhf5WFSsrQfd+9KqRo55b4A
qpp/q5wf6WsszQC/hVOUrxi6ne45JqvnOJYtSpu4hkaChzA7BuSDryfqFlrcdg+f
YjdobWmzKXuhtUbhPMo6uK3LbpIwJQTMllswEWXvBm/Uph61RT5kn27DSLQkWLIc
uNlj3t8bO+jwMPnOH+zilUT0o/RH9FVgfmV2ouzE+ZAlkm2avcIb3acXhDb4aosO
envzJ9OdJZicS4wiH9BqEUdKKLFC74vUA1hzuKCmmKy47orENAlD1aqYQ9i/6KIK
wkwn3ZRoObzZ3TIKgKZ3+jGfOs277WkrHZEbosKr/Plyshx0wG2gagEP3LZVUNPU
Zy8UQjoWlpovoHPYVeDBT8zr0f4bn3z/pmgEXdA6ZnlOuUNbjtICDrQIXWnY62Pv
b1hUwfHLHKL3vPxT5PxChn7dFlUDDm97Du5XQtm4JthjokL9RgUptGrxjL9BGAOl
eIM+a9Xbt5gXad6f3Ym1xKZZmbi3XBB9Q3CEgKCqZfyoFwz5N3A2/uy8FJ0N3Ota
DVR02CH6KJ/ZDgm+BXxW8bn7BNRx2nADmPzjm8B6yo5s2SMqxRNWqOzrXcMiruAe
DA6WibqrAUUZFktwmsoF5RSjLofCWNVfHxSKOzIz9Gg4TXda3ONRPNr2j3kw4/7A
N/xw0gg4pHmbpNbWfgQH2WRbhe+iK80q9HgxnnxKFfJakHD39mzcUxeOE4tNN5H2
7IB9dNwwPZHGtym+h8zjABu3fGpNKOfkcHylXoxkKH74GGiwVfdPNAcwZfyod+MY
MLcrAOY3hqOR7aXJvIAAW+nxDlef6aAWsxeWTZBZfYqAph8WxO43B1aHPMJ0gnhb
RQHoLlWJ3FEOhnhzz1Zp7BrIpH/GJvuaf4Bwvdg/nR8t1JlzrofIWSu8X1d9MLJZ
zq9+xDtWvOMv3wPzzZTS+W4R9noc+J6MJPzAcW3rwAdg15+32afjHWSRY71rIA1y
61A1AoPuDJxhSaN734EqTyx2S7SEDblWjeKVvmxDxDe22IM0zXgJ+bLBSPzhOSXw
ike+DcBzLEgBMNCV7+l3/gVeicJBE4tIajrfpJ+3jvnGu/QJpnR1Me3a/4OIhvnR
c0Fm7ZRUQWuAHnAqQy1jtTzg7S7YzmgQ4WNMMvxcpOLu90Lm5cgZtrdG47AJ/tAB
dgm7oqc+07CFeAoD23vmwUE4z0AJHMbY9lBGfPAbgzxxaKF4896cf0Sh/ccIuYuc
U6i6VweMs9gXm+nTPksZuox8itdplHT3RDMKjTU+CLBkDAoNEmMKTUWYW6NPJu9q
9Osa+v5ofSuXdI6D1FU5L/eTBFxJKY9vvZoh02TkfyK+KN/7/HTuVwrq7R55BKhh
6cd9mHzDvYZoJu5GT3pEmKWnzEOGhoSwm04IMHtVApZg0IbyOZpvCN/5QtHx8Apm
J8nkf57HUHThiH8cqzjtCRU7KHTXnTeD4b0AqAccvj5C1pNtdjVzgWMLmCbWjMa3
ogai1AY0aPfbbnbEnviRnVz+lxFZgLb4GHvYUUvBCnBCTIHmdU+4Lx1Jckbgpnbb
yS7i8ozQbPXYTv1q0hHAiKaOK/azPwIAw2Y8lqQ9KG24deTv6ETG7iwqQ0KbnVcs
Kv1Q44vlyycmCICN8SO/Ha9yDQWWPKH9QrWCR+Gl67aVkPhRHju9QVl3DVQsYaan
RZIXeLsm7g7BzJJoT1jXl4wmOSBc/4ri16i96evixe/6cd1dnlLoyF0MZCSWoEhZ
PeiS4+avzd4jsdW+tMqDuFZlzztxB13H6jebKvZ6Icipb16Xplku/yOpBh8lj6iX
5KDWcg43FzJdUWoVLYDAVdNTUz8m/lPM0wUFUIJ0qCbgmJOOsh2r3LX4ngX6n/3P
Nnc8N+bd/nM5BS34y0WawtDpIrwOaZADwHXvyf2gdo4bfJvZYAv5ozZSZ4WEoT26
2Brf0rdECmFTn1W3Rx8A6MFsmpIJznmMZFDWOu1Yu4rtlXPRY9GfNBXc0ySTnh62
r6ysjoHvZe8YTY/sgWZifTbUgsg2uVvAMCSgzDwB4bm+m5diWBLhmLvfPwOODN58
2ffuIVNoAqW6fVEaK05F13UL/XCxZC/Su7fbrGEgELVN4rQ8f04Ycvvfc53n9IjD
42mBIbiqZsSJ6yMiXQFlCwFzNlR0NDDS8JrFHG2JMNQ6U2EhUmMRuGRot/8i3MyE
75a4yyVAwaTS3UouwisDNQpposte1p/d5KI/5AkQByp/Qtzj0zojGmj7O9frp3Yb
ahCuAk6rClWnMFTKnFzvVDDzBCvP8rGY+deUPnxU2WuRorp32besIlKaR+xLJyHk
vXPUU4k5b0+ulFYFPmk3FmHg5pDVJjFcKPP/cwQpIpqiC8oowyI/ydfg3NB+ta2m
6unfIvad2bZUpauENeb76OsidPXTVbs2fe/8dnYKmJlAH3J/ArlLwMjL6p6Is7u9
NgjWZrOBAWungzn50eo33OCtnmKjtO8ROHDZxYTdGupbMrVfY6Lwd/niSy6isbux
Ok9vlYWLRZczcmOvroEKV7yDBBNriSH+dJBbFT/6Wh4AGoIPi7EF52WfHMnToxSe
iuyeDf1UFKA3hH1QDFViJY8A+iYJtaoAc+YwZDepunspWJ7vRsu7hEi88ISP9ux5
d25OZLnoIMDTrxIIscQx4z3ngw0UdVf/id0YxqnJWEN6zjKEYFhgh9wx8CEvsEtG
dDhvlWF/C50GMm68kAQLOrVnxoZT7Szc14nqS5FnaOFz1ThMRPtjXBGHsf9EvHMW
9Hted+IJmD85eApYyTJTa7LMqikBkwioyK/G2/fkOSzqWOe/iUrjIDABhkbyasRa
5eH2bphdzdVvkuzOEjQ6Fdm2BqqDd73awyBIElwGECxVVcOB2TVWtjjLFxu2uhz/
WdfcsEsTWDrIAMk4tMg4KCkUzXypERBxFXQgAaWnkO6Jd38eAYkHYuMBocMdMKAf
YVQ5QheiQkDsfnibdVzJN4SAwpfSq5ZZU2rJWdM1xWTJ4SdiO9kix2wrIM673z6d
7Ir1AQ1Hd6s+amVhpc/i3tqeTbqNk4eBC381Oa7RN6OCugn6ykYWUQ/Vrh0HUXVp
ynzPbVfI1kdu6aR2NAdO6SKPVEPAEAzAhszUEv5dPQarsSrYjvH5ChbaA5MoQiMi
oOfnjoAZDUOs7Gze+9Lybi7Tn3Nlsmu/g+J6VMg5B5/VE5WYV9ec4ZUujozm/XGm
69d6shXvZtZqBMJMQ+GFcZKSw7c2kK8exjuwEFNkBZu+XXvvtjoB5d0Eq3S/GjNf
QnIL5+bAwvSDNHZZtdBTZZAB+ENxY29LXNk39wkX6phqfmE/IcU7mPJe4MOfdqB2
MxntjrmxMvFx5+CECLlvOsQdGgBjS13a+W5ls2Pvuk3R2GRYNdTgAFrPaszzJ31D
itR6Z8gSE9i0FhV2NQvHklmpyTOsgFDpEh8oKpNLpB6s9/byY3non+r01ynq+PE5
g7U+NszQB03EnDsgnyg2Gj1xd47ZQ0ZpDm9CWZXyQmBHYwKhLEEMeklb4MZa3EKc
xB/kWjYj/cOBeVDu1RBUp9rtWTwDV1Rp3gZ4ci5O7raFYecupPCGNqgkHkBIUqqQ
wtHq9hNT+aHvVqBIRLNmZ6waTF96jScUpiDujFiiPmH3jyaAbT25XjlhGprEsOYa
6jNmysnZHBvige7E0aXg1K4MZQn6JiaXImqqSaZKaDMfSKOfhFKTkXsRf37y7JUw
Pyco1XYpL707pCIvrWsQ1CIc7VeEdkRrywJh40aJEnCH4z3KIMzC1WlVYhdZOgQB
NhDjdoOLlTj7NlQHBG+RigGZo007+cNcYRa6jvPccUiX/G8e56aMJKS1oRPE4ALd
m+Yv2+y6gabe33PiqeqAjUAtcAlV0B+s353OQn+wwk88aodz/p1Dy/R+jllEmDum
Iy3Hp0PUns5ed8fhA335G/LVALY4IOveHifDPYVlzfwuL6Rbw53iB1HQ2lINstHK
jNBS1rGPT+KF7ibwBOrBPFT9NVqm0xAXOAgmH9OnDn5g/cVykHY363e4NYVmd13k
VkTJ7JwJ3N5giULda3TTZETcwiAHzkUU0IMo0suHBLJlPMn1+dyeWUWSaSfYtuVR
FyW+gSrOO6n4D3o8bfrBKgAi3lpXfn46bc4cnZ8pugG14hfp6NqkVImvv00I/uJv
mjs1nzEBlAs8DzNjdTYJlJquKsN3gR538DIw6r6UIFb04QW9MEYlOYzGqs4hbu3g
AgXMasHTm8rNw0bkwjNP5PlzPAZXGDQzJIQBurLYE/udnh0B+HYh6UAjvVBnuVJS
4jwwl3fo3vtZQmXwO1KfiZ3awbreu+WuCY+4D3gHUttvRi1xIJ5CXg9O51C6DCTG
AJchMqCb5RDGI9pm8zVzh+1aFmcASbjDvvpYm+Joe3jqavZ/33vJg6GU3MSk0nFw
qMi5n8jcjrprNOaXyRI08QGjQrlORH0l95Ge8F/yR8JtXn3qpZRLN2Z/oUNJY3iZ
udk4CTVG+fUf5l6mgLyudqM3sRt5swNmX+XbvB7HBHWJW1KL8RyRgX7eCDDxp3Hb
y3sUVh93EyHCN9rjhdhiqJbLb0wNEgQyplj7dbVVF/MAI7fWgmwkTtRAX9jRp8tM
t9nkqK3f3bV2b31vygZqWdZskBj52Db0Bhz9cyShezqbN0Ar5LAND4HxptyQdGN/
HgShRiOHYUEBqOXigxXz6mzg1YaVMJL2m0lfSnobSNHbt+Ftxj0kv3Z4gbpHDPd5
6sM5F4zmdEOd+mVE00CwJ+tYalZXC1xlU9Fe0ROd08mJuYYBVa8G/0+Px4sdo/Ze
JBSmY0eSyTFmnR9PJdV3vHk+bjhxc0vWi17QhuxzJ3aL3yyaRP7VKNgzWRMWocYe
WVNTkxaQq3a024auEMiw+39umMicsc87dHRAwJ/dDwNV50bbYZ/GQKW39EBiZFqo
L97ppPRmYPBpid8AiP3opbXyMORCiL/k02SltJRrSozo52a4CjdYtYT7FpCNPojb
o0icKrS163488O88HMCfclpcsNJMEXaBWEymF4SNAkwXNsiv5hZdjW97V+oLE/Aw
/KXkX4FoVAxKc1Xw341WLl7d0Lqt63mzVSuaqcmYKXMxNlrwLukQi6mvOjJCk7RH
wsT4cSRAKe69FdHeqBYJWGV43ZI8XZJ5BwW+Xlap7BFhV+P8A8YsguUSeLzmWLTJ
nEsw1B5QDaFT9QROeaJoXsj4Y8mRdzhupFNonjANJy5Vznh7hvA6bRPnLiguQ/Lf
uexqdcQ7faRTfYmmcE+IGErwNZPBbHxBz0WlaiyN4e1Z80T+hTQsypa34Quu0i79
EN5HNqfuxkLqqe0Qq9CbR9qcis0HiZNsnX4Nvjrq52gHusEotGnAEDb/Lthn5Hbw
QUTubNVfnooT1xm9vK6t4mY58R8rtjIqiMgpJFxuJhGwbJIDAU1oVu0xtes+qbQA
vsqqa7iXsV8YEHRpppWTR8Nu1r0GG7JsRwNKP0zM8XfZEr0YEs/WybeHdj8xRmdk
IY8ljO+W7Dv4GUUfEqu57ZHhqJJEcSMKhRv75kYNc4Pg7h0NwEcECQqEywoeo2uJ
ve8j7RqOGoKUxMGVomNSXaANnFK3NsNMeo6x9wkTitcBAx32qgm7SsyWdAxmA6Zf
YAp5oe1avLl7SZzl8mf+kxw6KsXlH1fnLl7BZ4Q3KL0kKhpOeXRbAM40mpMWVOaq
pZ/nVnrqUPh0d/Y06unyM+PCK9nMQZRj22czIUd/V8ZOAR/ujS1fMxU4lSylP9Sd
hkAFzMlKtAxb73eF4FGanuanK9/rHfqyKfjZelQcYG/7C2dep4jjPPAbC8HHdJ4u
7WLPAjGV6zGvV0BiamDR3KNN9fO577CVfDl1YKytLmtUc/zP3BQW7nbjTRci6Q3n
eORvSy8RZR0wBKHeFb+VubqGv42dxi+wEj5XDOBGNITq6RSO6eX6AwPhPBQarTIr
nM7PhVCrtvkQdgV2hYKlyKTuBSrreBgS9b8f/wDei46Tlx2tqxqTKm6kRqrjiMvh
qXQB2XnPUQFiLakH5wqiijjbBe+W9zJ35NUNzbkZkWuzkfOGMf+tj97Lv2U2HDIJ
ny/QzEDO+7T/nqQAyERffwvG3S+ThCyXn3qqqviHEV0t5RRajN+0anJUDyT9wkMp
eGOW49xPh81jMrNLXxU3nqZP4PQuPu6y97+uZmJGx0mWWYSxOWLwSTvMM3hgPMlY
Kvrql7D6v0AyuvpBfLLzhl3eEU42r86O3JuFIC3tD2VlEv426BdWmZkosBdBi1ZN
Pe2oTTkjFaYjNR+MRJJCsaxAd3FZF3aixaacOydL4wHJxXQOMEkvoGaGigKhSccb
TY2pC9yPuBWlFBwPVXkL7BRJi0BcD+lrp6rwcjKixbsL5nMU7cBnhWvl6FuTjOXr
pEudmo0iFS19Q2FrPI9I7mcJtFDkSuqF/wHzrBhUIOGdEv/7FkZCr8Msk7COft5H
y294G5tfHElBtqpVEU/BB1bJLtYpXoJsyby+2tZdsoZj0nhdVgFrOq5bVdAJtZaF
io6S7IuJ0jSwj/Bvd5WS5xfXMU4mxd2eIl9kbH/hGJ746tL8fdCuP/2GYzgizYPv
pPQY/9OR5jLew+nFt3Erm3ftEc8YPYrhh34x7Giosv4JcjSt6TpXCxgVIfW958aE
rekexkr+d93AxbM0Dn8kjFqfl4Y+F7K9zxXLJ8USYTmWrKy5abSsXv+i9OQ3lCYL
duoskZKHJk5Q7/HjunrX3XTY5DNVpjXTD59IztuFu1R6XJsxX//RO5Zu3/SF5qEB
K17AgQvG9o5gDN/Bl62rZVjc+9Gqs7NxTL0D7Hjf7OXAPRIg8Qzow9/bGajzwpjF
9bqCcJxXLYtrm26DH2u5H+knLcDzQ/9AUxcXZF8Crg7r5txVQTZwFfECVDGEF7Hi
a7TXx1uDjsdj30TUThOJlUq2kE5s35JSo4EixtOxbsxfSxHLI0Oc8U+/AXVIFMlP
ehx/5eb64XjSYQOJ84INR5g/NrJ3b3A8ewVPeJeFwQV5u+9hogq/Tflmn0X7m1+b
t0kQazOAVN7ZjvZMfHkZvROwu0LqFiOjH2N4q7QOJcySjMEHfwJM4S11+IZ6Kv81
e6fLvgnifnTxmAeNr5fngXoioi3bammpwTO9jKgZZ7CxRp5EPR5nIJ6AcS+yS307
2s2Ebu3UszffibJfOfLjiIc5HGW100PC/lzR30V6KjmWZ2m9VAC02/YkP9uQqi1n
3uP3o+LshIkDd9jHzjXLxwYEG3K4emDgmnZGfWk5QOOi/klZqPn7UpeY0plOCAiJ
18mbk8AF4NLqSLGmB3g+Mpz6E9Q9PCNe3fdFHdF4kqrIdEJZOPjR9dfiJXux5y+2
+DfkBhTCGAZFVCVGeF4bUmCmmqliy9R4dZV3rVR1PZsX4wGJo0SMgQhkptF73jP8
3xsrAv9sBqgAFkPFsEB1EhLzFmmnmOrM0VS9yQyLeWLiASn/SggQjHxuna+xlYP2
L8HvPD5cbc8mv5+bnUOeP8CoVusxKYa7Iy4B+u45+Jb2Rq5LdE7BUbRYGPXDkRaF
EFQaOJ+HdvUQlXlfQzftlQfPEK0w+AF0J/MNPvs/HHqXRXDm0TGUu1QrmgHiNPAQ
iTbV7b7CAw18j3R+F28rWlWxlA3Hzgpmi2Ub5HTuPgtsnxv9gDkzN4IN9nxo0jXy
ggSAAcKytT7z2o4Lzf3eQeWLAt4bPF288nndQ2Ui7mQ=
`protect END_PROTECTED
