`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NcvJbeAC+1RnCl1MJGf8P2ZxEbQEf6va6qIHr1A7L1V+ew10GBsA/KLscHGrmO7
dKyXR9xg3Aq+VcYemUvEgsSSN6Xz8k6bt/uz4xoXM3AhomvPsuC7OW71TkiAASLs
k8MxzkebP+rq02Rmcf8NQ6VYNEkeb5GeVaJfR9gXCOlZUEtuQTDwFcECwstPYfBY
PT75b1qQxSJdjT3HqLjYiPQmU7U50kbqMcloIh4xYOYv5atZr7mwvoW4mbgF3dbE
EpehsiUBJwEwF6iDB2JPwxe6Jt0Z03JVe2Oh3oI2VKbZnxMnbinU47IKer7FwZEv
OEQO15+12sWI9Z75akNmYmd6v5ncUJWhHGtLmamIeXl4XBg7BeOwA7d2ZK4C7eeg
iHvAqZ8IUCSyiFfqLfiFEaULfrfFzu2yID8MVWnul69fM250+FsOn5MmQ35bm7J8
e8ZiPTuZGwrGbDibEyuC5rVezUsSPKStt7F09h0G3ZsD3N4Ay0v5KuKbmWqjWpzN
eCLpVekqQ8DTPL+07OvrDOVQrEOplXZEQSowhLY7/Tc8hhuNsYxNHkgnwRIRCZwL
JOvkZ9gM7YNCWqBRBx3V6TfeEyaBCocMtU49HlDnTOEr7WHgo5F9uagC4SBzXXfu
bC00/Y9zw46FZMJ9npZh4It23Wp4SezRnG6ekksTOYW4wKCqFryfbx+upRZg/mb8
cxTNg99pFV2E1bcH5COX8Zupi1NNwduhIVZoNhCQbIclhuGwSbKVred9oTvR5s6K
sGw7n3j543WcHcUtbtdzHM/Qh2+beve4DCCQv1stHHKrj2FLol2NLNYT45pFKddr
`protect END_PROTECTED
