`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwnrBAAYtrOK9eoRzZ2AQN0gAt1JMThRj2okJ+jOCUdg0r0aFe/qG3Yv/UtiiQJr
RivlG4iSIIVwIN1mQE4aa0hLaDxBz/fEf1Rr12MsEugty61O1UNP5pj6ZNkLU0k5
Is0uTsIozgYpAvj3mgE+9TRxFMF+8iJ+Did5zVXrlChMG2GcNOQdeYIeuaCnmqEa
YNbWzm4Y/GugbBjeSZDx1+nTXK/A8ojwM7m1LxVk+HJgzDxoDbdS6COtge4sfqqz
E+V9brddyC3hJCzg3ti4hkIwfxoYUghH7+/rAH/SI1hxrFU+mCZxiNZD/xYziWTp
gp/kYlmEVb1zTiOuCMf/FVInn1iCDIfQXPNAhGAtZfUOyVk7cG5Z7P5kvuBK/V7l
/cRktc+8pFPKc1U9cq118DDNQDx73UCclisTr+WzzL25W4riPcA6cKHFsLzCRh09
dQcJJZHdskdrLy+H7uOFdv/W/cxoXbQux4XL8T9FLpSpC5yGH4Wh4XxdIAscKS+N
vCf3tnVKgJAGo2BRXNuWR8TieBXrwvS4tPRCYdBhoIrqn4qOepS9whOMa5Oj7BaT
uYzesR00cctu6ipAAYcgss+YdxbNULg+Li5LH5eBlu/JtbcNNatKgusno1wi+LuJ
yRjr9DUpCvELFV0WYeMwuyGNbmwb9YjrgP31A/omgsJc6ywbbYg4kY7oXc3OIpjr
w1dGNZzO4NqSn3I8fvVY6OlLEMNwD7ywZNwbcGzB/f7jJSoqWe/Mu502yTtOlUMH
nmvytKoVR6Uukmh5i23mqw66Cz/UjYP7zztLH4KTvU0BMsdd6xK9Xa+XYEKfDEQo
rMwzKp7v7oEsDeTlxw07Sydcg4G2wMWcHnnFhRzcaViPnL7uecsArcCvMvbxkhcR
`protect END_PROTECTED
