`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofw3OM3nxU/5G8KQqYtfgSdh+7zzVo7gHruZ0LVxYCP0WJ5rI+cCNZ4J6ZxHvmYA
i7BFLxz+5J0oP+y0c9ZpQaRJR7QIF8hLSitFzzWfvLBSYMg7JOlEb9/MR21z+MrG
1y+EEfK4vqxo4uOlkcjMdqoOZZyIybBTGKWzBxbaQ5ihNAZKDUAenNc/rnN9AQ3T
J0nkSAyEOz0k87KcyLnr4iqnyPYlEbTOvAqUsWL9uxqv7Dw78HHhKJbU1Qg4CF1y
sFt32R+CT/RgFZWoiJQJ9bk5H1tFj1c0fb5ikcIJTKtJTYlHu+Uk37nOMeRBolo0
1dDFyzBFMyXleCtvrrt8fFE+Hh7IXysTBDn/YGRXQQriSbDRH7WCbUaR02YIYY5A
GuZFCRNkDM5bRJAp6D6UknLJBwt/qkwf8d6KNa6IroAQ2kM5+SsnAI7iKwAvgoXs
xbvgvB2ANAA1tsMBP2irL1YpNlfqYRNI/yGtkZjRT9vUNkRfryRZCu1xSoaEJyR1
Moh+5PMjj72H5xgiBJdcr1SXCtCkWdQ45xVj/ICBRTBfc5EgZ0A3vobyn6rfI6lL
M9dzNn5+aKe4U/PKAudmLZ6HV6JWxdb5afPhXb39QcOG9bAQfZtZeiomLmRF8YeL
4J4CLtuV/9d+QJWKQmx3sPWRvQ1J6OszMEWuKxYKUo0QFodrs3LNH5D6t08ljYBP
5eC3SfPzEnNd46MSAMt2xoVMw6djvTOMYFYUsF/XCZNWVaZrDyoU+2hRO2hztH7L
y6agAMAxQmeNDsxUYzygv2neCTCkjdE8QvEUZ4hpKyzLTyPR5VlrlE4dqm9znN9l
LAvESCKBy0JrV5yaYs4kXyUpFawSE58SuCqMbrE2aw2RKKktGVqZ38OudIjX9a6B
IiCTbRUUVRuefcscYmSASyOSoNMVklyFEA5Dnod+ttTljhpX/7vcqigJDTv10CU+
GwVBWzKPtKg2wj5LpvOYNhQBDzMLZSTvz2pDvXoBCyYvyKVVJXWu0qieZDoF6oof
Y3Fz39EMfHzO8VnxD8b3rFXwJNvpuJN4Wo4EJ9mYSKEssGsaYsoHsHyx2ERj6jJl
L6fXM34eUDNbqcClbc2MFwAPtUW7PEt9I9sRATisozCvnqZe4msuzOuaVEIu9IgQ
bsz/LQXZSFLyh21rY5+duWlIzwPUG205mFnLq0AEGIPY9ZXzkUAPEtLI7vEoQn2P
E7V/9+XPokffu/18AnIugyE/bgfQFNudnBj4N2LjxjcBw+mtwexjQOmTRgXJg4+u
XiyaWYFKuG0tB8/YHq5M2ZOGJsJLo2cJgcQps2Dy10wpoF/nBFzffKyk1+pqkLFy
RAcOAipDIX/Z8wnZfISw9PElsyEed4JZ5XVYiFU/Y70s7Yco5+gYIG46VRcUtJoh
epGFkUJ5Fo25nllXXpB9NSUvZyiPvaGOBYXbFG7/OZU4jyL5IW6zyx22Dlwdayd5
M4bNqJgFSR+RC8OY9FTR15V1ys3XbqWacfHZz6LAyRB8NrB/t07Z/vuk2DMPgibv
EnmNND43s+2csMHhCu2RciesUdrgUkjx3wgCOiU9Apl1dWhzxwcaf3SlZ+CrEUlB
EykZemjKkN5pR6BEeLkIeMVlyYgQDA7ZWAHooHzE1De8KQqDEhma1KYAVhstwk+n
PASQQMg7LRLhaypRkyJdFv2ZUt87O8tL4wtqwGJZPiRZHtt/tnfKFY5Saq/4nAS2
rZKTZa5jljQSEupQaTSndMZr/LJoxaEt4nUNpf/b7CZybwgbcVUcD8wI7I0txpVl
FGjJVHCX2wgs8J7U2/C6ybHAZMntW5XkN7b+P82LKMW7ml5pWMz4WqKDnRzDpGhA
Qzlb14QUXAy5HWh6mZibxoRni3vYqpByYSveulB7Y3PG8of+wa4xzRVLgMnTR8a2
Js4OaBuCpqtkWrE3IPTKOFBb1tjOLc8ougPlxxHuB+vBIutfbPnQ48XkoghRvh15
vIMccn8964ViyQnWDcoWiuyOMJV0Tv8mR3F7f9AMEI8+1VL6KKRox3fDVATnalpJ
AhNlaVhAV2dwF2ujV4shNi6nKquDUAlYznRxviU14ghQ8wtRJWJdiMYWtXr7lrn5
9E5c+zaxDnBy/B/HaWkj9BLflYoDySRCkEfYVXS4Eak7Kqbvz4T9TkAswlWa415U
+Zjz3/uQx2xiGcfOE0QXJCR+R1IXPYAMU8zIfNVpc6nyuPoc4bUpH7tO35l1Pum+
DIGrQWe3oMtdEZ+aDFIj5MHNX7HwpUhg/KkFbsHjAmoBMM6WIUDon9zVV8Zk5hFx
HlVvNQIcyyB62O0b412FzpZIfh4dW0UBTGGr1JBdUNwsAf23DoEosAamSKTJp/R9
rZU0lVbPt85wmTnMn0Pb04yMjM/A/+592aMsZYVORwund/VUCzxziisIy5F/tx1a
ETVaQwzBjuNL7oLMpJTo5lKANDIjxDJs2WHJqW0JZzozdk7bd+7tFrRgf/GTFUhP
3eXOX4PDE8wQLEa+9NjLqrnIA7zIJqO+4grWc60OPWX7O2ez6WjsUrW2D5Re6pIH
wedGHUCSAUUKrW+/osN2Agm+GCf3f9Py4KGYLcrNp2MwvSA6Vd+G61/HyNhFLgWE
mKZxxlDtU3wCHGcWDUNiGu/4roMmPXmyDq/mPfuPz+5eMTmbh8TNdVed1b/EBcXG
++r16tyiXMJjS7jTAatgNZd5/ltwDGEWP3PimreBuqLIW3mDD+HLTN6UyAeYahLA
svqC9jDw43rPwqbe8OWVJYDljErvMUl//ZnSCdoQEKPhMzIGsUsegmL9c6065b3X
50pvf6mp53m7ml3YFH9ljGFm8YQwruQ8r8zZ4PkebNAbkHLGOypTHqujVAt2WB8F
gggZptgVU9sdxrkX4ncD10vU8IOvrhGdIDaqkdN/0ZX7LIHklzqVUXQ1ViUE+D7D
vauH/akb60wpePaKbWSxeV6K+Y6a0/xLZDAQ2UKzyswII5hEU+j5OkmtkorI7FSN
KHm/zJ+8LMNhtulbWu7FC7y1vR6hACGOSe3CpBylsYWeZ6mGzoPD4LReKTMhVF3l
O7DKH0beIrNsqVU/Fd7AvN7pg2tsiFcbO37XTVQa7jSUYLA21tZQaN057NPaWVbe
/WpVp6sT03Ihi6aAtgp7cLkK9fsHyD8+ruxXQjvSmyY8DFqupiL7sHnEVn81CfwI
jCxUw/t3oumw7YSq+K1sga4wf6kac/ZH/REmOFlbsFRiJS+mNX7oOrBYULMz6rrn
yF7zuVvTaqKe+dWZWtDCQwjiM9gpSC4Uq8Ykop7AP+DiDExvyT88tSZSocVCTDP0
8jtlikBZs/8Cbs+tFRjrvqBqvcS3FGe9ZvGLDLvbYkL+9eenlrdnG8wk0FGkNREP
l9yzFNs4DMctrDUOKRJnSV8W/XodGk9lXjnigj6zjbLHCnxEKMcHMCc/NZfrSZvV
sfeuAsbrFy9OAE2F+GUHpc6oUafWMFwHDxNOdf4BmX4Uw7Hfz9IKGBJ4Gq6C7X2Q
9TRlqvxhC/KKkISOluCyA4W8pVFNGhBjbZxpeRG8mhsaCJkRgQB9ptx+C8OiPjKX
pUdDpGCvGEIqFMOn42okmuWG8i/hkqX0vE+hx2Wnbkc31J1Trs765SaRvN+W5Zl0
rmZyokVpw9oZTyTYJy+8xAUzmcNTmYPb58+8hpF98zprBtpzgKdrkhsktK0sa+t3
tXJQV+WsCSOFTZxw9DLj+uiLw28xqrMp+7QorV4d6GNw33/FZ22bGEBcGnmRiYgO
dC5V+0JOCaqoOsvbOHUlLFY7ivca5zedyEJ9rJOtUXk9+fsRzq/ItFd4VtPT3CUl
1GtjPWOO4aaH1JKZ76tR0DGXYMKUtwJHl16Nli4/CTZvHLywwHhIc0j5Kg5iGJRI
F4g/eGXpuqSQHxwmunFUgkwwTgeSvhYJ51aIrZym4dswPyuAySeJYIzdspTR05Z4
ghTns57tdy5HGJbhWMMFul+P5fuaEF2flpWG7GKiajNZSOVUMDP0xC3XMjT4UGvj
aY/gUGWEcRIuPrkNX0qRYcWpYjao8WrM+ZebkHlS/9FjZuv6FWQnF3RMlzAUx+5H
bxDDUCkMs249ZdDJT6U/cAJM+MFXUi+wVGvjAinYpAOEoK2pV1bSuyVgin7yGUKK
mijYhf4ABoD/eL+4IRIQGioP9NaVD1qirq3DsOHVT+XfQWwFSlJbGjOyRxghuBFo
FyX6xZ8+ahpSlwhVnjGa/+ghLpDNBHwCoEiyttgx3VTZU5NGAayawlvbEVXlOAQK
YAY30YoRtVl2QFGeBkcp/+OAI4Qiqhlvd+nnlifdiMmyK283ZwF9aHXQEGvUlwCz
rx9BFkL+Xc0DnXuqVR065/aK0GzQekc3SVPbyu2hp/u71ouP04aA7R1UuPgP1pCI
IrSFdtQhxGT2tiiHeEQsgsbrgTaTXAe1IA5IMmYnZA/t3GulnlKLOpiJ2VWFuDW9
gkpOIOCfQGdn0qeuTPftm5FsIVt9xj3BPa72O9qkDcud7o6bcTNfEu76zyRPCBRb
wQsZpxsgYCE6h7387O+mvHYiqoFq4iP4bWfWtzk6qCeot76cvdYo1yTz8OCuqRX1
632Hp7fsGRlP8KidT4d4rDwRlR1q3Epm1qY6c8H8jnfXUVyNmaGDYyBlWmlQOTBS
4eZ89hB3nnOD19ReDQGvM2nMZZwwchX33Agr5Wgg/mOIhE+q7fqZYP5CCkK7aen7
v+qeQSOmv0ioWzI0Y324CzLu+fK7cj3uN1xuDgBerR/5yywtEFMT1loaR6LUWvR9
99eSXcIJdx3eN5KR/uHheDlspjB3g0Jk0GnQbaiKvPU9VmwaUOzMeZW8OpdrgFPa
BNODtD7lq8bW86iaXOQAWYxTIF0t5akfnbqZFKc3S6Rt/WyN9dIj1whyX8cOjoJe
miSNqQmD8SdNf+Off456oHKVGVj06WMXIPRDZdE6arxpABQqRP7oFWPMKZIJx+QV
w6xdiZAsK3BODoIDXM2A+qjtE1S2Jmff6Yw06Zj7tIMDKy540cxgadcEDoBX+SfG
LcBCdY9djBJfJUtNwrwW3TKX7Z2GvxONklJfKyXYQovJNAm578fKEBTxaxbML5Q/
0DFPg4aMDsO4kc/Osb3qWMOf6Iko000bUhA6v6mTPj+0WKZUESpgCeyLa9mH4cZ7
+zDvRj+ItP/FzSwwcbYo4ZB7F7JJXn6lsP60etJ270KfdfThRKAx86KY+Jrxz3fM
yKFAIYtY9FtvIXlltKT+ocMPAIYQ2Illib8VVrOVOBoir/WF3KkIlkwtZXbSpryO
ZNd4CzNHBWxSAW+vO7LdV8erWMR60vprxM3CTOD+h9M/Lyc775v6EoSP6gvkE8Ll
UbRIInVpa6c03VQ9l1vato4l0EMnsIAue+CJ+Ds6YGm38iv63gM86sPXIGw7FA3+
9c+SXqQuiwawmWbV/2H0PxJz6ARSRr3DkY+Qrj2dZMeAULOuQ/cG4kJHcZweO80B
gxjBnxtvhTUwWlmZNhxQeDiIgb6s6N+3Dg8q9MTS+TlsHUOzWv05SH9iFurtGBOs
Z7C0VQxyXAHmanQrdpx2W9/IM/+r+jx3jO22zDjjGWhK1zObs0+JbG8bjyo6WkdT
9U/0QqoaWYw30kSm+9IyeyJGheOZo7wF2I/Ac4pc5jQrr4Ra9Hv0TpzuG5heC+56
ztqG9zVP3i/DHiLrPknF7WWkaacO4miVFcVmQ3L++LeJ04bN/8jsqVKZqu2mIrse
kXDRwGGUbWcbVrIHQFecFKavWxIiTRowHpqVA9obMyO86MhHkZU0LxCvSwxujPMb
7IFdkOLU+cXtLUbCtLj9bmclOaI+dynvHAQaPSHMFg3wFkTui0MFLV0I/MUQDI8D
xRi2BOWKxO9sV0+eOT5h2jqmK/o8FhZs+jUkJfmSRRyzjxUXSKG2XLD2DDhfT9DR
KaNbA0r08I60QRupgSsQD84FaemurA6mkypqTnMTPTyXQZODv1EAPs3dLBBc6Lkm
+OKIKUV1NehhsCQt3W1ds7VQGEO5fTgOUXgcV2InIxYedPvb8T2uffzlzI5Tj7Kq
bAyXDp76J7Vsc1E/zpMsyUEhZ15z3OSB1j4KfYe7U3uU4FXUndv5jSj2bxo1H5KC
EQgpX8I7ZVatU4SYiM2hptw+X5QOJxiXj8iJ0/luyJEWhc2CRVFo59Og9hC45D6k
odoGJdIy73vdR32pM+myejuVT4dpNg+kHkos1jVnWkvAOUvLs38fNyjh4UTtFdEr
hTzaBU0I8ntMjexRRzotQ2yaCKvjXN86yqGMQJBr0otO3KUx9w6JgGT/srLyFoSu
GLw04dW5s+ME7MfJcPkPn0wGBe/DXvIby+ct26O2gsB4hqV2P1sWBr1XrrXjpwoL
YOcneNimH3IGzyh6mLfCXOtHPKZCrxW7gEFIEMW32Y6le7J6PHpF7m1VYZaivv5w
hqnEseot7WoG7hgF2j4c/IPCQ7nAB8Hlh0Z0z7/ZuA04J81I/GEAsPfJbkmrtVH+
2wioPBWGs/bZfbwwoC9QUN5S335RGDAbE0gejArwxMsNl4dboOUsxd7KWc0nvc87
8xAV3QJJQHnzflCz04chH9hGrgZkmU2hLm222R3MslBo7jpKj3C5cyErsHOw/k1v
ehoaaonhMOXTESsgR3SqhAgDjdfHsI6QcOc1bCn2+yWuwwmsSUJ3fj9ewIao5vxH
Sk7EMTDrWINEr/Tc4BInaIBaMVf47Ja51/jx4HaALCaYOvKAHZhqXSCjfFgoksfa
ZLficEZ2oEDgovOaK18G3Fl+RWUw9yg9WieeF3NFK8wX9TFQ9yVO++ruOAbUZRKH
w+HyyGtq2jX2pAiJlX7akGHlkMIXCO+FVrg0FzJ8YWHLc4mz43+J7QpBIGxQBrH2
zO0LO9QaOPounIjdv9tNl05x6LpXrlFDx0ekuyKqb2qedojMW/OHvlBSAU0HFgTw
IaFYaps6gIiFGyCnoL/6IBzYEGdsOVLSDQ7ZZEVI8wRqqPvZS94YHGrueFr8iy2A
fki3vLN2Vz92z+pSSPPAje1G4eG9EeV4JGuCKal6iSnmlRdp4Zg/UDwgURpLNbZ4
F+j1xqkbyIrUobQ3P2y2Z5Qn4LPGZ6EDSQEOjuawBS5sER0zjFxPcAHH1iMTLEAQ
UIeOInaKjhsFOUMQ4PJcOSY6Zs6+9CLpE9cpSu7eYwknOIL3O2DnkBVneLxr879/
f8nRa8IKl7nhP452EYI5Q/b7sBOrFcUI7YMFRli0PdAtz2zifN/nDcCETwMQrPFM
00BElqVoRF457oSVDq4PcRh+Pr6VY6JV5qfeC9dQqM6NJWIoi/SpQWtj/55142U3
lAc5GvNuaiUJC4C4lFVGjfNglo5R2t/76OQwAZXCSC50p+6iD5l7F5PQ1KCsRPWu
Jp6d2rlIc2fTee5GOkIpXIk/EcUVZFZ7vmxz0Pufyieu++2gwdUcH0Y7ySS0TD+1
j45mlWwfJxJy2POr5TJ2eZHxP5qnN3lWrLQ9rBAuOzf5gbq1Y5MPrG/asInHtFvd
kvPa/9AuArKfiq5cOkCwbVzKwVn1J1r15qbZGbq6uhSjCuXIj2Mrdu4Xw4/2z98l
1AIH/a3f1kW7QcbHQo9Rz+GV3ap0S0MA1sNRnwC/Z6/gZT30faOEYrythNTiZv9I
VVPbAcc7smkiB/Wg5VKtbGfBlt0dc1YUlIgsmzSTqjMBZm3ujGySRALMiDGQwDlv
AdhiCgy0Pfwvgg2XHcWfB1axTCBMjlg2tdnyFug8TnnlV4IV5gQUyl3cMwLdBAKD
IEzbH7q/fFQahh7/LvsGesMgqbSVZZ1gppFoKoExD1Tq+6dCmMWy1x0hrvoAz9JP
69g19Wp87yGaIxO3dcX65q+FWxOa4UL4zJfl4EE2+CRTTah2AutdYHXKsBukSAi0
OFtDSx2cfqAkLRWpPOfSSLCldeKwEOw/dBkx6aI2GSPXiBIZV4nJh0Y49wFlrIJD
5BAsQbVjJ7HNY/W5JCYtV5Mbg7VCJ+TCkBIy7/fv5u6Do9JubHEoNKsxq3tkIatb
IjT7Hjvm5+vTNqE10g5ZLuyNtmoA2PMNIZ/ocGV3yy0foJx8N0rrQKbQ1ZBDbB10
kOkq5wHbymFOSlueW3URJgP47a6VdPQd7gO/c6GqoGVV6h9H2/OfRY04gqNX7+cR
HnbqXxlALPsHo9wCB35aYUUrJtZ6tsnmV94V+cFqMiUnihaBgT+HHp5eD7OGgU1f
uZjTC5JmUiYuYcZG+lYZUCMBjoOslZKvhTUx5maCzQp7g0vkS1HLVVE2jq8elDtA
c20HymuTJFpsanVELOtZlIQIq/kLCfesLInH3ZSrm7ZSMeEscdmMX0GbHcA0Yi4p
ly1udMJ0Am3uvWFenprp4mLXwx4+Ysw10bH16pgtwZqk/Fmi8jkhRs0Zn7ROX3LM
zhvv/yAgN9h80KyiMVK3tf32EZcn9PlRUedAqnkJZcMKBK+aWI/26Ub7oqI2xSn4
0NqSVKN45YuNCTmngActQ8FjiA7hOwKmVTOv5HowZOUzYhFjVtIA44x19CFzFhTv
Lw/5jgdmYur/AVILUft9IfQr/6ie9g7soWI/HrmcYIlIr5Xyw6h9MbfT6Rkzn/Op
BSLcQQMtxU6c2Fm5cskXN6Eoj/uEgEITM0gVDqgVXKZiL//bZDLhiwmxpX1MyK9+
kJFZwwMFiukzMB6tRAx68g/Q0eAk3cJPOjybtlSNW/N8BaoR1akNdGSJbZAHud4i
agUZPccq+WJEFLtGHn6TXua88Dmg4dkI82hENSKnLSjIKhaD6uf0Su9utxt4AIMG
l7tQEJ+fv31Vfjzh883/AUklznrTIAA1icEk7bTLuX8FqevrM5i+ejbjrrWHvt0l
d891RhWdloVi0gPZz7tNE2uh9WsylU/4FJqJ4NmfMUwisG5snin/kJpwc7SYlyUP
CyhZrG9pNpf7QzMBvTRvKZX5dO0PBU2OkL1Ku5H1s77DNWy6Y790vFmzDVKSk6cW
Qu+auunXmVe5slkNh2K2wu/pbLFtUZ1MvzqMSVC7xPRveRljijdGfMKpLGmvHRtT
HsphJK28LX0V1TGU1g5Pnu1nxAY5JNqt+lzCm12+cPK7fNDazNObMw2JM118OouR
lT7BQw1dNpxiqNnWUjGSkUAHjaQEFwBncq24Rwpo2nio8aRUCjerGfiGBQVwrPcI
TKmjsC9t4VfwKMxjeti0ZRC085Pt/fcOOosIas+dvnk7M++wAjpa1ZSmI+Ui4F9g
KYw78qRVU63BTtOncQ+llRoVgJrZBjdRrPEZBRlQwlH9R2hiHmuneCyE47F2+pyq
PmlH/sP9bVaZpNMnufhm48YRbzVQyA++EVwlaVZrNN6/Zq6nShgzGIjAxs+/5Irs
WE1os2SglIrzK4H/UX7cfdzh8PW1LgU3N+DztgN0YfOe612GLw1dad/WPj4G99NI
paPOMuPOVWBVQ5ofjYejWdEmo7mTsclDflqD7s+Dltqz7RGoS+dl8F3t7rmboccT
kuZPU8zkAIBigotQuV8DW/IRaYg/GtDS8IqjG9VDfyF7LtqDtTaa9DwK02jIlRlh
JHm9QRA+PZX7zSt8rEiK5nm/EgAiLD0NHOaAZpEvS0/DguSnY/3s4X539tH2mXgo
osPyNaXMTTk4uQiAwUSFoh7+p8p5Z3V0xywx5Y9kw3tc+Zy5pue3bYCp968ls2Al
kT/BnUW2U81hI30uZkVEFZoDO/K3X4LQP+YirG3hBiUh5PU8uhVxLetHXK7v7keN
9y5aa+x/55Jdi9KBH00lVKdHQ+xUeZGr5KduI4YjAiHaNV/XZl1/OkrtNn26ZH5d
vPEbIOxj4nwkczLebUMVsOhSKssNY627SuzdNvWpS3Adjht7UrNzmbWupseFLbTf
+K1jegsQGYMeFreZ5ptPQLv5EGkenQRC0aQPe+IJCI2j/9XC0uHAIz7tRj0YXGyq
nJ+rGPTrLXKlfbNhWQtS3iYiEvNEg6kgC/1g5fEnqkZqL7GrPgIqGMlTPJgSz86i
1ncZwzS8ddJLKOv9J67ELZSQZ2+kb3MreDzbhyrJFtVqi+Zs+6e1+sVkMnsoash5
T4VAJuP66ATcavu2hbu6/ryuhFSgixYqFTj15zyMolvut6h9wfxRhD4+mzGi82lh
AwsRV+iA1GKTt4MAGkqJNtVqiBk3j5wjQdOO+GcoXLblP7gI7gHc4i0Cbs1Bjpca
+uq2HSlRsmgdh4RwkOjf3B8sR32pEaMp2hbc7HprgizOfl7YC9bcOsvfSxdzPW2R
ywuFswCBjpA7nwCYHb9aOx3ys4uWtUoB4gQ6nES3RpehSoLgry+AejU2Va0xYmYo
DY1RLlH1prIWBAziqKN/L9wzpwwHCSQsYHBgYcEZ0IViz537nTZO1a1yGcaP93bX
Oklgh2OyLo//ukmzmpCS2P0k7ZKQjauEZusEdgsdlGxNOWstD5ipt4DTFRABfRs9
ED08/TCCtZ8fa7U+M9EGUYYU9U6B8KmOqksY3RphyDOyWxD0u4sGGELtvAG6uKeU
WdFv/cpggXzeGnQby9av7StnSs0HmG8ISt11/uwuEtNfc41tvJCIT8n+J4zTCkHH
l+TjbUjNpH1/42OFGqCiXxvt2SwCcBfm/55RiAuqfUA5vz08gjpcRARPaRyVIdXr
N1izAjQBrh1RsyObBtGCDneiqq6MxU1qPynP5eDJb0sbr8jF0x+WdNm2l5CDSBpj
MSmkIXGm+iKSTanGG4G0eD0tBRg6xuowQJAEqQdVzkbt4cBGzefJwdba9+wD/3Sb
hmM/cxpc8SBVOT3Aa8BL+lU1lY8bhNyUv01V2Jt0+G/eRUrSmGOSlTm3aBEGXAOX
2qFnPEoPpInvxvSL/7gG4RLvSh6GbMewqKRvHU0Y2xkYYci9mnHuWKhs8k1+1kXH
hK0ETLhnKCeMCvOHL3BqWi1MHVEOSHeKWX3VM2HMVpcU4WXtNZJUgmJa/rT+Z8Ge
yBK5YivUtGNOzzl+L77XORJxcgGYlla5HecwqQrJovTY3KfyWt+bfaLn3nD/ncGx
ZbFCMJ3uwLgDtlcRNqobEQK18E4fwEaxc4W/pVyAGvpIS7w7in2ICMW4VZ8H2zUn
9jAv2nlSnpiWR0l/HrUl+dWXZoZ3tH38Y0tHyUghcaghbyAyI5K37CGbY8IFF9/S
gr7rEn/Twwee6KdAPgS1Bs4E0zgmFeKuha83Ok2hJz7s/DI/NnzgOSys87mjmzHt
q9Z7Sn0zFarVXkBMcIN1/huq0wccG44Lm0RHynsz+g6iZ87f8lJuxRJQ185iHLlh
pRAWEei/LRk0eqfChk9sfw01WxW04CA1SA+I8lLzHNpeFaOKLC1RAslkNeg2vt1w
KIKn/or00iZ/upLNs9brNzTKONHeWqdhWTUEjRMghaR3YIQ5jxuzAfbXBawBJQIU
RywxtAWCOEaKHS+JRQdYYRcNQOPUpWU/DbIejevzlHyw1jAWeScBUMKV0Tya13hu
jGFLDb6VcaFmwPBBIk08e9hWiArDv5QE46N6Ji1c72I7MilMCMLlDinNW+1Ux7vb
o6GkfIQ1InL2+1EF249BEmBJeP2UHhmLfunimaEKXHGehtr4kO8jDuwZDwKxmbrc
qx6tV+iUrwH5BJzgcee5R4HsoGLipTziBaj4kEDKl6GR9So15n8MbVPq/ypxkEv7
hyOoaNve9mvz7hnsm9rG1p8JUTLi2s0ep3bvRm6W8BdHtmHrtwNPfkVx+hLm0nzj
Rvi/ZLX/xjzdJgLG2883bcsF36lqQRT3ey9QF4iOZw3cNq2OJeIZoNQzr+dnwgIF
+OQZEUF/UXEb7kPc7YXaLLit52CFfU0XO1bv3YZSLW0PHMtGlczJlv2EeLIlrmOV
3Qb0aHzXL5N/tjyvsg41Pxnd2Xd1oQfFJmdfynjqjBczBGmeIlLY3Hd91M/Vb/vq
sB+lN7Trw+1oi5iOpymr/QyNyoJohmS5m/vAeRtV4+p3d8Q2TBHcQtTCujolBmJM
aXZw/fL+ycN6F5p/vJf3FDPiwqQqRVeQoFUiixoviOeYJXxzKe1rhrS4slEDnkEs
VAVvgxJeou0cBiXQTriWKrUh6AEf6PI1oeVGpOzlZQIK3CjoF5w8CI1CyGpPx2s2
i4D6LCV4KTmh6PVW6PNjHPO9zmWjAod8mVmxN0RraVnRjfZL7hJrtSqa+2g7j7yr
7qZ3VR0zMccJiqx/yZVIxNl7gA74h2ZPY2224Ia9070WOReLVlpnEWAgjR8qQ3L0
VEUav+c+NHwb7D2FxcV1P0nGcjffCN8Hdy4pSDzcTF689C+g92RUO/ctzKZ4cUa7
MuBxFQeBDsYhpfxz+gb7zrUXRzep/WOTOeYbo47Jjf8eqoQQ/WtCF+/FKo1F19Ec
lJ3rAKCZzJQEYt2K8+kXbIdYip8x+7hpRuPgu5ez82saBjOcFOQIk4ga4bBpEAPm
w++r7Ckv1ZXuvePDXAQoQQ==
`protect END_PROTECTED
