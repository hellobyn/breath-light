`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nzy++SAWB1GiVE97KlxsuaxOIUiXaN+x4cuQLmstGnTwazFhN0/ECFrFAY9vWyia
TYoZboL3KHMqkLas3o16BAvcmtsH1XO8lblDl8CulQX/OXKEAWg3MqnEfxWlp3L6
pUo1gC4oGhIvnu7oy+yTdwJmQMq5dqqjV3xcJQGWxaQvXDzhkH5Ls51PKtARMmn3
DyrcnNg1fSb5bAnqvNB6VRtUScKSOMBWTzc/sdN2Hj/WNb0cOLfU7gTc2liH+cfI
FZgq1e0YrBhk9VoqgFGfiIwK6yWvH6dF+aw6aLvrKKb4J/PgDafI04e1MRyiTKF0
ek/No56VD/yaPa8oaBu2yUi2B+bTNRS5KtZ/uR8f4zuIEUaWUc7S0eDLuG3szotY
BygsDUP6jWLJhLA6obTX50Th6auzkSlzwv8UK/sVZyL5+/xmvrTK1RQv7dGM6ryY
GqJmhItLAo0NPrpHQ05CfvR3zLHt5sbjVVDvHTJcwaRf14k9dnzJ8+kudQvmUrIk
+h4b+XGcrMf/a69PZzktbKUh3EKjteQPZL75g3d2FhyPyIClpQahG6xl+LcUSt57
AFpBc5GYtXlCqQB3n+SkqI0YMni6tIRTHKQ2Onmd1Jm2fy3d1L4J4+ZIYqMwUoN1
tBZmvdyf21TxrtRmG6nQpqJV6xGzo1Nruc+6jbFLzqqPqkP5AVKUWTT0zpOQ7LC6
TUPE75dxvEDgZmkcQ1ok5Up/Nx+vzZakSJjRlchhTBIYOT1+/uRsi5rmxMWtkMRX
r3sZxlcAtNDpwSF6+F8yvD4vb1F7GKI9HHwtBhQM9xt9rL4cLoqF+MQtkqqR04mh
`protect END_PROTECTED
