`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSLKTsaPjSKFWCQdEHv74q4chO/UmeNybX6IpBnuJM0r441j9mJ36bwKA0ObSKLa
cJ38NTdF06GLmjA+PvOwnTUOh0uYDEDdsO8DhTmbDDwXCOj08hpO8rNK7zxl8j8z
M0gK715OU79/+CFyMMAvX9v1rzR6XsKkQ1lFEr/I47Oe8ZwjrgHIB55m45TvOySI
KVY6SBN+BtBL4OW+qleFsndNLT4lwlz+vdTjfa5POUnPg+R7cj19/W3tEWks46Sp
gQpeoYwEjl+wBDU+WXXk2PCMUzyz4fh0rVlbsUWokYxnI9b5l9oTiyfKTzrWKL2C
OCAk0nr945PLwxGorGTUyRTyPjY2cBBeYXUexwjNChlteIHfOFpkbEygOrln7dXW
pY/J1ZMNrbShvGYJPXFJZVy87n+BgRUWPe6TogidZcdVIxbpoRC6MPgY3gCkWhij
4VuU6KcpFxi9DtOj+oxOmQWV6EhXE00ojtUOUbSZzKW89AXvbFYK9MNbgV92w/Jx
TctvNGdE9HmNnnDjEFKGNoejeg++1q+19encgKQae0ClQU9iYQydVipTfndmRINd
mnP4owqVEIi2gUymuTK4LS2ocBjX+TlWJKXZB1DIMkgxd0FZxtqpfb/AXCOa2OIe
idQTIDE/I6tu2qArPiu/2lv1JAdnhrgpYrspuToHstu5XACNZ0PDpSXgJjfe3JOJ
qTFfgHlg2xLUX0vNOau5Obs6ZC8tgIOoU9ET8JXqZcV3vZIaaRu0YY4MJChi/dEY
Il59XmYoE64E6qGnWg0aHabp504iKe3c5HppfeBR8Vgw88NG/IXu6TISEpsqFJ6Z
G+RGkp9vWff5TbyB715tz/vKUyh4CzxeT7Y/ZPl0RQcESozsrAF+PobOl7S+oh0e
/hMoNT/9ez/YukDr+ubVdyqVzZ0F6bFTNE3G9LOYQx5PEdqZ+sMMtO4OjulJzkkZ
`protect END_PROTECTED
