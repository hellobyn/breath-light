`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrRlVCOWBEW2aRAqkfFVzx0uToTgXaVslVFAF5N3f9yPTqxosB7VM23L/LLUnUw6
taPwOmCbALQbMiQ8caCcTFh90nSjOOJGYl32RIk6H72WkBPUCczEc3xWgqLHEjRC
q4GfP/KL7fiWqpeCmU1lj/wwOXbiYze3YfT2MEXT88WBwLKteFJT2yyZqJIgKgCs
AhTX+2AZlt3wWRypw+0Z5e1LbBXUwzu5iYtVf0+CkF0ppXLyWh2SU0FE+jckeMd4
aWBps1Mz53feHkUq8gUdVrd4H31mPFNRyfcMuzn4RcS25JTh6IZpO3N0Yp3oM/6q
kzYH/f1zQlKe8Lf53IJtVoDcQ7Cov2dp3m8nKLPCisRsOObnTgh4cGPfgpWvq7Ff
XZToSEyhB8bKc91B4EZdxpDo1FfdiV1rluBGzr04WCkdORu4+l8KUmKGwGTxpIBS
BtyqjW6axilJVbr20m5bgJVqiod2JGMn6LlaiKOCQfYQUnuJWBxBzo9QhaRZ77Kr
NfRFBxSCpqK2MCQ5XxrM6UdDoTjRZ9J4aPblQ1gseBS6mWZmnHtvN5/btj1mUIzb
EokOtbAXL/HlRXpQtsXWgMZZgqtthxLdSd688zysrRKDqrZiswkqk1VvrW74K7ti
yxPk/AEcuhBc2VQ/1y0k2d3sRdCxTi43pW8SaGQ27NnfspcxUb8S6BBMKx26GA/D
JwswX0rrAF6Rq4kZhfCaUR8moXdhLoKdVaqqmsn8sDWh7y4mq8GsXlJyxOW0QNQ1
+sbCDGxuMd0KJpM6Zf23XqcWDc4VOJPRNXmPcsAihzpJCqqD5jZ4+IbZNYbovji6
rWBvrfQx/7ML4vl7MUH74fMgAkg3F1VMsLLSks6SX94F4aJi3/IYWjQhKBWDFP+7
30ppjUbVjjLJgTxBgxNBZhGu25r8pFJNtmmsBExoMWb0Pf79BGJ+VUpvkjiqILRG
HI7k0jcxhKknDNH5zk6q84IvEV+h22BUe102xq9PlbYBPAR0HsaqIsciaqmXYys8
YlHHTFDTz1RbeE4JHBm7Qi1JXt0YD6tQCl7uh7tqZkGOTdGKS0at9xq9zSq/qTIn
ANFSj6jz4B2UHtgKXF9Yp4yNFkpUuQYwCP3IsQL5Rjf6ksrE7uhxkfDe1S48PhPU
hW58ZIAAgDciQATj9IQjpSlgnr39MHk5ae2zkoQ7JtX2dNHx5SFU6eq2U+/yoqGS
NI3Ds3anGCMRKp7hmH072Ty5Ioczgf9meoeBuT2bhuTJMR+nG8ANXSH4UT30X1w/
VUgjpBHkT937XbxwB+f15NIAKMG5HNhvmWT/5dYd7ligphMUoQZVUXZjOdmxKoxi
n/3uedGkT8Xnf/0RAng/cPtPpk5NHvYP5FKKGo2RFH+dJgMtlonZymrptTLFElI5
OEMB0N5gwwMDYJumgvF06v5lnfEhL6iZYKgsgWtDgx9EdsQbnq3Nd0hBU3a44sJc
Pa0QT7mukRb3FZk/ZoC6c0/YUopT7S7WyU6wtGy/vbACNsmnfUDD+aE646q32J3K
zM6/DZ573I1L+EfJCljFG0KC1+oKytVmkYt4h5s9/tEzoy5BUXRpByIWT7ZGe9M2
En+oFG7DMhlGWJddxxdyQyRg7TpnAUgLr37pOHKAX7/rGHwgTg8ial4PDrRH0yOX
G2jXdXNdYLu7+bP2YmqHVi8cjy63tDK+m4c56L+PBVqxJ2HZeDR8j30NsDK1wTXx
TkVZJYiQTVxzlVYue3bl2FIXYoeGujvBj8zoA7AlLyYUH79fW9UX8DcInLa7eacn
R7Y7/9ZnBCjO0K0cwW8uWdvb86T9pLmAB4bqiSw9ZxNovfZjl2Xu/gZYj5Uhyenq
WZuycekz3hXKwIiHQsmQVYfEDg1eQBTaMO61tTnYmlg2bFgm96dIPZROtnlXgxp2
WvCLI4GFGbGrUaG+9d5PbVnEcKRxDsXVm0Z5eVDarBfe6DnSRoSzjJrmNYdT0ofw
9EDL7A3r3+YD3+i5FqjdJTOq6X/MveIK4ZRh/kw7jYn6LYOGyicV7qdfjbH3YCPv
s1GoC5FhHTI17PgWgG6wMmJJoebxH9yALwkdU2wqtdimAW/kSwqByZQVqb9UR1hM
lhm/xV/q1OIOvXCIFLOOwvmNxy4+aQ1DNc14hPpRmcxRuoZy27RAGZ7s+GboOXdh
ngwGzLpEaAUnviOACHrnQn0GWMbElQZUuAP2dHADQYLj2StYYwvBsggI1n/UepOY
0bzZ4uHZ/U4+pM5HuXEdVOHwJsUCC8jgnwQ8VifHXflyyLxyq5qa5LrDCrpwRHLu
AJwLXdoxEzrXP0S6E1DY8wk3J1Jhwx2IvV3z2ZlsAsFIU2MVx6Gc4i4/eWRG8J0H
zlPcl2Nvme0z+G9fDGu9Fuiq/5so/H50EVdUqH1mTe4gbcsqZjpsVWdftdRpkAG4
KD041olekrMOyJ229z9LroWJt4bHnCdVWC11umdePgLH43Tp9IVlD1aOLnLt0tl3
UrJqk6MWrcISuR8FsbvIHySLEhAvJ42WTwXiPNi5Vasv4i0mZNhP9cGtXoR5SXWB
LTw4/YDit1G8Ccu2HeQ6TMo8a9KOkRcWghKI/7N0ZMPck5fEIBvXn+FnMo42Bz2E
SPYWj8s/b40zE78bFX4yg88lfh2ry34Jm3nfsQkzBK5OjjRDWz1h4DF+xvopjk4o
AnUyWVk8k0xD6am6XbCTAKbuHnBANxEl4aA7JnauRUfGJ5PkiTCJ+IXPDKT5k5ZI
l5+6x6+IzQI7T8YAJejA/eV2y8HPqbVrO5Wa3vx31Ox1o3aQyT4Ngg5doAfIvTWz
QBH3kzHXlnRh5xZ+LAH+sy4wDjtZN3DM6ovQCcEMpvXVcK5vuOYXpfIuKV317jV1
BbrSxW+3WEgLgNvhqm3pX+qgvo25OskjXs0tC9M8Kfc4T4ZfH8TYnUAHEG9sr5sQ
2smFEM2XxwF9K1brp8ctGb1b8z6lebMNDbFla4ap3vpXQmkVpYUNiTbtsV3Fjkvg
UEE14jYR4ttmDDRXVpFXO75etyfvOeFDSOkimHq9YOpSPFVVCEiybOXsawda9D3Z
h4p81rLJ3b+oo1OT4SZGc0PpGoqM7KUXxkYAjVYvs3xzYaNVHDCBmQoDeI5bRczx
ZKqU8vZ/ytUYB7ppfvAnbq/N9bxE+vqfgWulR8YEejtahST+cHu/iU67GUeOpC5G
nqWE6lNi8nC+NBkAGR9YqR8lZWm/B7K3/qNfXK4y9ZC4h0YD7pX5fBvURnAs9BLi
GwMzpx1u40NYqr4zA1vkObvgGqH4DgkyUvORiPoPCz/aXVXVBoU49wFsiOlEGvcM
sIDJUG+EZxF5HEyPrACPnGWXl0xHtJKQapTjxq4KnUwF0HYdZJB67Hjp7CYJALM6
aVZkst5H+fCIY9HWVOkqnnwa/To/m31bH2PB86p5DPQC2Oq9Q/AEzVVSh9iFwiCi
e507v9toV8xBnk6fyRwnT96oakDn9jwiVJX8IlADG/CEn9h3pPAo6U2mBEA3gWNx
xuu26K0u2QP0v3tqHAfo7+Hs/zfPxdLFyN6j8migSPbnbIh0GHpljR2QvrSmeCpU
HwEqfhQ53otqoCDf562A0LoDMQ1jCXR1saq9oZHa4qVM30aq7B2EhEwUrbLn7x6e
vZixpfxtinzwGzOOYw1j4vCmcsWUzAwRfteY5o6Xr1AFXp/vlWp2gJ039jAzzVzF
d9em6jFe6FBxxP8m6rkij8Q7N+D6YcZIsmcMmdZFkUSy72+AwuBYCQ1AhutYLwWM
D3sRR/5AjKM7wyX0Q6chHtBQ/mLWrvtlm9BPb7KaFAT3D0aOiIAfDNEEeehUukd8
dvj5/3lTHNWHdXWji1ZzqKD3MCrNH0me/sGKGPvfmD9Ac5rZBl6yWv3EgqVf9LnO
sRGk/mLOjBdyxy0djgX9pu32vvVMdvtXPHaf/PdjDs76fG3WIi0CqjpSab3Iq0a4
Xe/WIWy33GH77pH/eJLgytCuZeAt2pNul1bbnJTd2I29Z4lYLBp+5QFoSZUTGQ5k
57kMDkhCyJ98bSFSGbqWuuyeUzQ6ssqPppaEAoZgmujmLrSeLeW5sHA6qFsaIZma
EoU0HTXlmQ8+2KKBfqSfirZ9LGwJvlttMv+9sCBHyVu0Hst96NUSmWSy5V2oU5MY
vbJlwePfyLXVjqdkWDWIkzxBn0gOcZ9WItlolbJ5mhv5VROMeNjRpGPAJu5VRbB9
phKtQWSgtJdTsyuUz+XOYemh+anjutvX4oujkJFYc9diU4HDxmWNpoThdWK6/5yI
J1mLTEhylYTp2UPpGx4u0Tw1ru+Bkec//f8ENuc96tg5vN+a1767xwEbBNQXD3DH
sbDE0K2qxS+mdgqdEEg5bkaR+z5QRK7kcY12xkPez3qucFNqGps2E+HppiDDkP2W
8Rs40EhwBOvCK/cOf4P3OFxPc35M3gPrcIv6mtfuKo8mU8+JFPh3aam59gnXHlcP
NuLTysD6HmmrhYGidE+j1m+aEtBmsoQhbFh9lDzUf23VX6PA/ZCyH6QHooKW6uJQ
+ZW9CTc31K8uJPkSJLFYx37KjgZ+wGiLofHGbZwlEY2nfBL6ngCWKrobtEsOz/l1
3Zl+K4L4RzsR5zj9bHkZ3+fjv9bpjAoexftWS5mWbXObGCXcdXOIHekXKoWnZuR1
p2rrTXF2ntlBAusJuC7ciF6MZhhyUALtmeeLOTpzIY+V4sBDZb6QnVEu0msel+Mr
qLBw2BEe1fAwgcNKlRC3HGemujVxtB4bSSbRyYGdhdRVVfybRE6JU/VPKAZIRt1u
QDX1YqxWQv5493zDb/nQCmyn3whgztYpGeZMVDHZDuBtmmkTWW0Z/jUlP369SEMM
C0zekDLQhLLljzdALGX4HlGXqur20PCiJpO/uFwPs565zCScw+WPACmPjp/8WE7F
Z9/j7LuEhU0G/CmQ0SsvCXG2thXgiwUJt8Qgtt/WPxon0CQzhntEwj4fMkqAxG+t
Zvm59ecy2wvDnXnzmWrit++HRazjNZxjD8LIDWbHmF87q2gEmbWVK3DNMbFg0Srk
ILOjGteiU1zdXWYm+4dDdKW8uYybA3TozcLG4LTGT4pJegeKEZqEktX17BhjYxUJ
IY0sbAgi2y+j/E+WModTW0CXXxCtaYgSj8OarY6m20wH8qFPJxWLCc62Oe9AkT50
EqSdfKzAbw/nqKK7mVElZVxtb6iQtU8VWo9fP7nrQuty6b+gjs5lgvU6vJfKPm8U
wZyWH7YLCQfeYUjJNcgs3V+059k6F5ViZxorA/i8TKcLz9iKHzyJffjxu1nqhBsu
szY/B20ZrDWsTubBvEhKmyGKud/zq6SeswuAVd+VSandJNVG6pDuwBYjGnXkZdhJ
qRb1J3L2Lce6Jvbnmub3g+53N9sQ/s1ukDn6Ym8P6Lc5x/ZDQYS768o9P5JjSDxm
BdSyV44225ttbgDIUBpvzehJtYf4Sj7+iBChj/icWs2miGWk43piMGc+KzmeD+BA
sdkRibjdfsv4/4Al6kmAMyGCe8Lnu5EpTo3qZqdCMjUn32Zpb0oAhtpESSbllgk5
qGF6nF2ww20TPaQzlaipOqur+SW7+qHp+AvZaKFk7vZDkEKTEA3tiCTP3FICMeEe
gTxiWLtFRuO6+Ab6REy2HBCMwauZeL2y8GjCGwwzW/3RStkrGkiX2YY/BRoXeRgj
z2DwAfKyryS9hUYhczvfU6QshDQdn1FC0RPGeYmu5lqBCZVHv7RfTaihdUjuK0Lc
1WRplwRGT9o7zna5n88cjq12SGXhD1Vw2EisOBlpglk21BlnB9RZUUW/lKg5WUgH
cigGMhtlnTn6Nj3o0vIKkA3iVNOf3DAFsD4zH56bS1cntd1h3BLaQj7B7G2Dt1XY
K+BTKqHNC8M3ffucdl3M+BmLqfnzuQsIr6ugdMTeOFwWYs91Cs2Wt286QQIei1U0
nw6ZCUIbqIgzoufwX9PbFh9UtQyNXIXZJZn7WgGSG1PfMGxrExf+nfvZnk1RhUoU
YnKnqZV3rANP2lOnUMK1E9IqHKDB0HGldvaXQdd5K2PG4fbBhnE962rEI6qjq/wb
+EHr6B6vvzyZnCAg8k3qu/vkw+p0hfR0EBLQm6fhqQIOCe6huq6cRaL3bE91gDnC
YwA8QBlE1Gl61I5ay1LVaq6YyI6HZ4tkK5G6a/un7PgrwupfYi299XSb5IqTY67K
jDQxYbC6hgxHWJKbioOGk/hjIELsEXZxzmNH0UiGiVIqYTdxdocNfNujTVioVy9G
k4oLobNj6+I7wNwjhyw2kq5sGcXJ4WEuC6EFbiB7NA9jFGmTvmY/ckVywhd2gTWb
5KifCka47upYWgW3Et0UCJIjOIPHPyL/CUCBvejHEhisz7emjyyitdf7/sHDRZVF
7uyhhUeYSW+NffsUTq3u6z0dBeMV5MjJyJWUILNjh+1D4RPdNnNG13T6I9qUlB9e
JaWUSnFT0JZXXEnbcDmt4jcnCjoE/lbAbNHLLJpVejLlx/vBW7p5s731Le0mNKrb
bd9DombOM9WZistGD9ndggy1Y1NyaZsfmwW3R5fxR9sEKmXB+zp61sXpHb4O4oJ5
O8inRnT5PN+fexEL7wS42W8JZR8SQ/ac7vLkhPqhmqaMrdr/w573SUeljwx9sh3a
bIDNEmmRMqJh77GQumCYqTshV1EShzxvMsJoWWVtg5plATgMTtYnhh6NamUaFUAG
xhRpVbi5qToJ/8Rlt2+XbVRq6HZouWG7dvEEUkR6I2YFIDPzHYfV+WI9m6lTPc2c
Zd6naMdzbQlgfj8dYS0DSNImul4pwGNOWchvdDn8mXruCed4LopUB2VB3cqkghlO
GfkQui6iDDdJovC65LGVboEkbFYnNuME4jsbSfIp6ADFaryRkwHRpP+a9zxZPOB2
Kc/Mb5KBWng6EVc4kME2Dnnt1IZHG9EaTPQjqia7FUICdmh/91l9ACjy/bHyOOrF
Lw/20xN4mf5TUNpZtB2JVwSC2OcYWT1MRapPritYMerz4Xxk6P+p11H4W9kFCHUB
OO24NKzAXK3KU4n0bTwN7dKReKeVViAbbC/Zt6D02olrq9S1jwegRQcMxmFBSQNs
D5DhjVt9O3GEF6c4sG/spb83N0pYGVvnGLoAQkGGisue8YW9Gbsa/Kw08b7Gn91N
0LIqWbjxIK9ob1iWiP8azPyZzgbRgBF9a2RVPhc+OpGfFrCTA3g5i18ap6isB5gP
FT8nfONuq0TIwfwYcDo7rNX1GrSvzJ15ku33itju3eXGjntksbwSIRGQhodAjzQq
PQi8fsGX9kThlEG5p2OoU2hb5QX9RimjPNQrrphnU/8QZ+udDJj5brjKcg7A9l5F
B9BhUajfEMn+Sslh4/IsLbumUln3OzBtyIVwBux6GCGIsJi5H8AIznVupgvkPJ6s
o5YzbDhve3wa8UnHeZvcUg8uoAeAtl6HZdmPkELGZpzspa1zmtdwsNLejbecVmFb
dxgS3fB6qlaSoEW1PonnhH2daU6hpyoXoPxpPJlbXDnmIJo70/IUNfum6wW3KLS4
Jsdc/jbHvANvtrZsAgRfboQHzD2iov3ap5QJ6A7deOnTk1Njuo7B8/ik4dyR0gst
VUBe9oUE9gOHaWOP3hAoTqDV/F3FgTt6DEG8Xu4eI/UbHc0Rj3j7jKNUVzNiRakd
ZTzkQPRISAVQdrp58qd8Rhp1egN5OjV2wIqCVKsoER17VyvePhFjsPEnJ7OelC2O
pVuAYvNXRaYa9/2MTJ/NUIlYLXiKEXWv+MRcorzCJRMysXkxenCBLXurADNq6lZc
d0CqmnMRGtxnx9kYZD5e1fZ0EHQ3u7GL61+u8rWpXpogFhe4ntexEFuZ+MWJgvYf
oiXrqMpN7pTK/xh25HWv6Sq56Ch3NtAmhQHY5SwWmQjqPqULfJIOQQn2IdGbeOHy
2WIBgG5ZsRNJaWhli/os6XHsgZUohbrKfUxPHr+UQQ/sTlfTLSAM8paFGioeca6y
qE0E0wlLLoxvE1yna/3l7QZr3yNeks/uVQqzP0x4EUnMeQgOarzk2URgphilp15U
J+qabQ0RUJJ+FqBHp8G1jY9NGAuZlPTq8p+aXDVV24W6Yd8WWDJv+/Atz9Dxd6ES
Pi/M35USJqZxYfxchFu34UR4plRPOaShdKC6XkxCWIUEHcaUJ1NVMweYPkB68jHs
7L0b8C1h7+wWHaKVA7732WVlCyUWcwKfdtbqAo7R1A7B89S4livQFkHbUmy6pSy4
7WoC8EvlpGBuIhj4zavQJw05ynWp+QsRpOROyJmRe9QWXbm/6NvktS2OPk56ZzRG
nMryDJcQq3ZlkGReSmhxMrFY5/iRmS657h00VyfV6iglLJrIAI3dQ5Q/p7/1PHxn
UySwqh0F2E16HI0F0ChAdRAa2JEIi228/Lufv9tsWvC6lbjVWWtSNVXCHPaiI/Ww
WVlS7b5GxnpHCIPbNwlDNaZXL5oWipCx6YfqRZMgVEEmH4CpHflLaoSNhc60ham+
oCMtxMEK7l9fmoMMQjeDlbgdqK8V6eeLqpXPbkcNu8SlPC/3QdpkdyknZ0DJ/JLj
5nnr3cHv5Ri+u4DRKiMFZUUB4+OmtdZ9dkgiuWprdh1OxxS0QhAAKIMOD4c6AAtX
9HnB1LBOueuXC9cqwvejM0tavwxO+ATFsEQJk8OcvFcPJPqxwESHT2wrMD1N7+v0
1j06kx3v0vNu8rcCM8qM84zMGLMf3p513uiI3aBbDWW2tU3CT5wJywyH28nOHyKP
D19fK3DSW961XP+EJNldtERjHrXkc7rc+t78UzAYFWRSl7PHb+mHm5N6mXjbPWMq
YAjtOKx6dOTQCg81ZvS0nmaOd3ZJlqDoKY67iVOC75O6jcK8Aop4DC4X900G2d2q
K8eKyOMP4+TLA0Xfx4s2diuz485pb2mBnV4l/s5LlUQd7YNjV9MG/qDz87Z2FmXh
D7m8GKLcE+0Bkck5netRq+f4s/aO+6eoSEmHTph7NWMpB1gmGyvnSFHZtuNQO/8b
nr61TInebe+K8xiMa61Y6g==
`protect END_PROTECTED
