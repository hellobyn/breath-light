`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXFgelFPpN9aZHVBcGZE/CXuQBcclN4cyZ9LHVE4iL95CiScmw6pghfhwbUYceD1
6cIddhQHGRzyxTFIo3LthKDou62xeuh8FMeMX8CRIT2PX7qt+GdcvvFkf2qUCTCb
Zzqxh5h3KYeIwZq33Fhu81xKQCWkJX/IhORue7z4d+DzZ6aa/cgM/hlxwgDtNpQS
CR1Sogow039VlvTZfEXqhcNlGno98Em4JNxOmxJbREsC8fjRTQU6ea1xgcXruIOs
4U6+d/dZpQUPJ9jwX6NQrewGqI878VOIMgUdyUcrglh2F25Is20+DqCA5LMpWzfh
+RJOAhbiETojSBcLtN9EADxUmPMr2q4/B5MuszN00qApFM4iKwumg3wfY9lD410R
rQMpSg7iEeKJoa1h6ijGJAqgGU8SrgyPWZe6QqPevbFA+s3szynEnWdZvZ97fm2p
XZzAGX+gtds30PW4Gqz+6KXyhVVemD0WIP2fzoeE4PPMk4l6E8ivJnkAP9o/DhKB
7W313ztP4I2pybq2XtsMIfFNAdmihuwuUv1NSoJxoDq134/GLvrNLTNyTQaVJv9Z
VoUZhpwkWYNJ5qDYnHqUT+YkMDyhcMnBGxCiX82QF6s5HboBmesAZY+uyhmpijip
oykCYHPCvyk/KZ51Plhfxxqaxr8vL+TKyF10nKdPWNLquKDVKn5iixj2GyAg5PkZ
egnlmNkw2A3KHNRLGIrNuWmiS1cM1nCGrEyv1SwwIycuzWPzmj6ORaz1OPgwXtvL
Bod9T5pwg5Y7D3I0VRPRCR+2ZGD2uIxRbR8w/zKMKPym5luNrzqme0rfCHbiwRyf
IhRJvNp8gyMffcm0m/miVj26ldSNFD8CHD+kEMQh5P4ZdT4ybGTpqdcw/fl2Q6vE
bIprn0MC1hVklbOQ/x6Y/FXkLyTkcQYQuzOYZ1w3AwL7+k4kLjaf07T0zmA16tvD
CKfDVHUXerldu7GbiEhT4aso9T4666LJ26DKhjI1XOJ7EEjsxc/hnT86oWJUVE4Z
dyKTrNkCWzD2wvd3+DJTaSjDWtbZuvnDS3XK7z4OxrsQA+dD2/TXLVsCzG5eBIUo
PYOfx9m8qI2WslQB7IehL/trPRMjpz5EpuTrg7SUOuT0D8JN3rbCcvm/FL7Pc6+1
Tx7GnUL+oSHmKM0xUeSFGudztALloAGgbbXATqoSZii/S8SaWBsWuuQQeP+ZgVXq
SZ45fFeVDQw6pbklvZsIMsDP3e6TJcnRQChYu7rEZwTsfyafbHUxVzN8eLLquOpt
ANUAqehv968N6lgIJAye/FqUTDwA+5oMQr5TfIsKqOvHfQ+ITopCQtpkE+qEc9Ci
WyKw4pwpV6p7Mk5EcWuFs8eAYvuATCPs6SXeYnwr/bpV7PjVePfRbgyaSYTiV7k8
mtbqCjRi22EOIETw9Mq5HZXUje7Ct7X/R5wG++nJcr05YD049wKvG/Eh4TlxteYc
1MSFWQvbtzOQtUpyWzsQ0Muh6fkFHgArnJFdZ2iZN5cqOizQxccvmW0a7hDgDZ9E
esc0AbH9woWTB8kOXFQ7vibiM0fKd5adAF+NnDEYha67L1jPbIe+m3eOvMIBH0jO
189T0ephOvZ8jtr2gZTs1VPJZD2nOOEZeSeipjTkh9SkQyAUA6iEU1hCI11ljE8W
at1//4bf5BHUOw8bSneQ48rchiAefgGpSWK8rrefe6I7V37gyCRyxe1CX9mSV2T5
Ko7ZEVENEbtgYXtsPO0PAOLjsFcx6+qgj2icCkQ5dfxxZl4z30VFOWoXWtdIXEFZ
lY0j85ZiQfDUmXrUaBx4X1qIQ3Ggw8pTLgasMxG+zwl6umb9PQKFgb5yaB5AO8gb
XqJgFb8RAZWuDSfNGgSv/C4qwNhs7DYZoi0qqZ7fpHfbhdsmX2Vr+vOGVD0L0Esz
SPOw8KVzenEDfMjS0bBEg019Tv3Llg9aJFNFRqL72MxHCVWF1o+vTEa+GP3o0BTZ
AM1MEoJQz9fCy5S0CP6FJRIA7vVHhNDka/eVtHIZYzypYlGXpzfnt887t1HeeVW4
sXWWCZ5hT+63qqrfwpZy6MEEzk+MnJfNlBwjPizIQE5a5gNpebQ7k4bArJjZ+5kj
TMrdI0Nt/2Dd2yIeZyiXJMdaNtaleIqV8Xg+7bgCuzHnOw+h3GJf2THKQnNKb76X
2CIoueIzyNM+S+j9fjpYV9ajPlVaBbv0gh7VETwagbk06iwIuv2Xb0wbKFLeIkiD
QToCtyiupv9JCE4Vfj+X991VnPcKdM/csQGLZo8DG5vEtlDsjSjmW2gWcZLuiPRX
RbkeAWoTBGzGpMyG2qQXCUS9o7J+Do/cklHsLeternFh82viXTwlrNN9YvajaVNw
1pIIv6yPGVPVSSLP8KMZ+t16YmQDq4J500ZTAMccdGzp1yf1Hy9xPbIqrNvozPIn
oM1JEb4MNIK5Z5us7tRZXma+Ray2ooVIhNiovCTaeo4=
`protect END_PROTECTED
