`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RI9aV3xTLJxHrhL4mmsneKzpjHIu6bOIc0b0xrpQs/PMMtW/dDQZUx1/XACFTacL
jC2g5rBSeMO64GEtx3Z6bXztUGwUfWHST3DZ9zls+G+v98G3l5MiRJRuMcQaF/gt
CJJ8XMK3lCcZebTb0EOup+P7LupsOBTpppHQBm9IzXIs0ezlW2PoGw026kx0rrYI
qcVdBNViZsQqARoFjRwezfrlSq0lKafroD7UGVE3HTtU2Hj3opOuv7q1iAjdS/Na
EK8W7AaGZv10v3sPbam1mjEB8tyNPpEbh9MQ7axjwpAA+9Lg5OrtJVV4FfDr4JoK
j2j5BuS/N6q7+Mculq62JauZZLAQK/3mRbAeWjfsGK/Fu8wuNFYWy3imvmmSN26Q
b1hYTXuwfnPMionB+E7dxleC56DgX6eyReAbdFWyCmHr5fpAyQQVtthlTOdDTJjK
16VcQL2BjuE5W6b/k0scGWOTcDTKABGcBtPJbt1IUloQOkazs2y0GTvpmS4zwIpR
JIhuolUy7hp2ZcPrXR2vo8/7vehJ4Y/TAd/XJsqTW1/ETNPNvJSFT4Biw97HxFzP
bPLJJOOWfjo41XtDkUP9E74oYU+WOaUKSoIPvX5pqFX/0Jzq7wUHmIj+vDihYiDd
Pm86rbkyLez39FZPAMIOivYqWIG0Pk1XoV2H0XEJVRPyfL6f1cUvBgM45Fqxj/Kl
i/zqHNvHNouQC5D2Bf4VLTn2JIGNVY4ueBNyUv9innfnCIEYuijaDhMEzxm2AFv5
dEeIWps4jfnDiibuOXEIW8WPP1i7i6oqCpVRHS8nd4UASGVVl1H6BB8I6ClsRHdw
PliJmnk/DiLsZ+pMvuRUzQ==
`protect END_PROTECTED
