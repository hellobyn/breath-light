`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7W04iSl2E4ozOztxagDH/ntWC42H5eHNPJ6q7Ssn7idu3cz9nPcFkzxTd2e0hAp
VjvYkcc18gtU8bG52KIZheNevqfiETB0SkHSv4ev5MJ2Z/z8BvIdL3bj2iy5XQi2
ZZjIFLt0F19Ys9aAD9qPLCYxO+U5RcD3M4Nh43Y3Yi6/JWMOuck8G7Q+A3fDy+Ls
99pwHksKKZqgeOEdllEMhBVye6KmFyX945LhWgZOkDgtYUTj6oQBWkd0P5vycE8e
9woNvQyeOJPLUhbGhfYt+rXOCV09W1J9HkSO1u3QvkVdyUQUAgbfb2EYCqmuBUjM
gg9kRv2dSDn4Wgeh+kqvVkaesk4klHIvdr6hUJcxgBYc32EupmZdMvFIk3hdYCzo
xeE4QPm1k8rzsQtPTL7ZlK+t8rlZ8dHBC2tupHul/+u7WMhFCBDf8MM/JSGDaBYA
cPGygfatT59u5W/jplNC2KDTnp4z/833luXKUgsVsChUKYWa79QO9gqKa+jDzWSu
AyavLzbNe3ClQ4urigTWiC5tyH8ouIYCJof3x3T5x0+t8YzhOI0OFDagIhHnSqHA
gNIrJgEt41njn0mzlIHmsrXTamsGG4OB2VvDmXOdMAz3ay+fqDbFOSZzVVLxUWHE
kPghvNZoILi3s+WjNjnkExEH5gqq1JHJAxB2o6tFK5xOTVFmPFnX51MFAMapq6Sd
0+Wt7bocInPECsspL+o4SiUt3b33AFQKyR60DOYo87rGvfEsVjKspS4kZu8fhWb8
4iHBwbmpubHvh0NZg1L8yaySUwXpPsH1Md/sER1lCQN42z2MdFrAy3Cm/e/mGaau
CYa0RRqzTaRDx0X4U++UkNEqIwI88JN3SlHhLW70Tv/Zg2I11hOpDHCSN3EQTTsN
7ERy5UTPryrhZCcT6U18vRtj0DVfo20m2QGxtdaEBwOHan9Zxg533z+yiS+L+92y
`protect END_PROTECTED
