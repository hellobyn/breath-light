`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RntVByIyBBlWD8oKQXEbva7NxFHlwS6hz3Ogvnm91FgiUT7SogED0kbchfvdeMOU
1exktx6N2GxzRpzVRG5zeykL6jr7InsiaC5J+RbVXBhPFKa/N6lhA9Ybi/EWqlbJ
CO0jZlvQlzvayhZq7fxXkjR8ztqNY4KYdWufGkYsrnU7d16CgOAaljDVBvs2ZwAk
mxT1uE8ThfQnyhWqzSRr6cdHz5pB1a0CJjIINTx41oCT2htcAG+vGaB1cG7Y4tNC
wFz/UTgD18DOT5oVDi0msH4/QCfRr3W2z7xdZV3BqgdiFnbhsbcPhPDfBuT6UJy6
s1PySGTwsTw/ysTiqteaFIiIqPeya7d8OCgctJstZV2frSSXVpX/DNrURDoW3/Nd
O13FUAwdlthBXNTEf9g0jMdDGTeqspQV80Ke6UrcSSbGC+jz3M1kfGInvtAiR2Fw
ZTnkPXx0wDRZla/5YSSVjp77I5AmXYRdofPgtd4GJ8E6k7JRviFaemYm/Mi0jFRL
YZ5YE1NuCnxwFyrQqjsTJX0+S1g7m000CSDe4BREErQ3SSoVeWoj8gv07zOqk+m8
AU2HGREg9anOM1g1WBqdrF/i0blDVsl+2s3fIK6A2c3nSPevuC3e1DQGRdH3qdhg
bTZcbXt6M7eNvv0xwS2rS11yYETWsBJMqlctfM9R6Mkyk/RIWmdkPA0WGaxXzZV2
I0lrQHzsrC+IbOjaCAivEXD6vwEL8fG5mQnyl0LXkKifTtTYAaKC64EHx+7JRwwk
i2sMvmkObH23VhcoKWAqfeOnWYH9KjSMZr7jTbU+a3fkWZMbskfQINjm7VrzU/sG
olLYz/9mNexykavLQwRhZFPlM8TWRWWC2CMCdU6qoiSfIfYQs/smOhTlgZW7K+ge
gSS4NLNy3/JQLdX+iRL2z6j1VK9lc6iMjzsIEfRirqZFR/U6EeigcAgtx1a+BNlK
l8epmS3kJKFf8UvBlmDY4XN1EoGtxoOE+dXUOiEYAocTw9fh7qM6uJoRmUTyauh6
KBQ+E4q967ezaPqD71HoMRm1lLGzyj+Lv0of5Xj+vBlgfuL+e+VXQ9hVnsX/tqER
wcQU9hxjd70nC89TSIOLhAKJ0LpcDhk6mg/TLYpvdev2uV+gtPYi7L4+NFWlt8SA
rqlVQEJkVnfh0pDmRaHefc0hNQicgwV1P1w70nRGVuXMbZXfyHWEH7IGtdrXlOmJ
zogNV3mHat2NEzGfvFI7VFTDmQl4GFTbNANZFfgxEoPtU/tTG8QjA7oWXL10OPCd
q0IXQUobPFdB9VhFK1lzMenEgmfUjfq1D4biFQdFF9yvM3tIrn6CyUcSPEr07Zg3
y6RYG/YRu8wUvZdXHLS0tWWSXO1/UaK8DnfZDZ7439WMc9hQzCJCHCI9xs7iy2iR
rSjo5D1DoP9L65GxRaQ1PXtFpvQ6P6zSeIpCwLUKfQvPodpgXwMGWV/HIC9JZI6a
MVxKa/mFnwX2sBqMuvHGfW8ySGt2PY12PWsVfz5DLbrBvqUDgeb3FX8j0OSb40J4
f5vP91NMHwgTgndtQ6uRM0X/oxEUzPri+joAC3w7TAruyxEG06w8flOpW/stbMug
KHmvNkZb4Xzi+ASFQW/CN63JTmBgq4afoKh7ixMxVfKnMEt2fKClaFIBvslnHnsr
zOpGDvMMLXHADcuvpK61KumZCt8wNdFLKQVl5zMmOCNzxdaJildR1ed+rK95Knk5
vi8yXFOClV/Yqi61grJl67w/ulwm9+K9nzkR7Q/j0DCTWM2TZ8Mx40urdrz+qeZ1
VVr/h8XeOHWiZTM9QcksM6nFjRrdda7Vg7ZDARGkUuYBiL9VcSOxLOPNufrlZ18u
sZRB0WQayohSH3IDNXw0y6SIpE+paJ3KX+CD9K3dGrT/DxCC6J4dvX1T+odIsWEm
0ntG/XCDNQ3oqX1rxhyCTRTDvg9qjf9gG4/QeNSFitFrZfriNyZo6t5jA7Ty+be7
mAqkjC779rJK9vEidW9dbRZ/EQ8OWEP9UhXm1XORQwd4CC4pLk7+Fb3i5nfpRO6s
ISvn2SlG3T9VkkkTGKJJ/v5rnpdfHUU5SEaJ3W/K/NR8C1oU9qrjRsZOGf1iM1xj
4Mv9O0Nmoea42PavUzO5NyvJ98FsNu4l5ZA127AuQZ+mT0Gv2gfXsDQO0xD4826L
bchihQoAdoex0sH3U9jjr3woKxds4trwMuFNE241PZDwH8iDhA7QUufItHYCPxuO
swQERgnFmBO4asurA041PvbgSISrluB24kmSJSywXL/ch3ccsC2TY706BzLU8ITR
YXBdrgVOm4pM7D9K2GeVvuCFQ9KovlETIdcs1V3QfXs=
`protect END_PROTECTED
