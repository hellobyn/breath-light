`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UG++y5qJmd8LAJMZJPOY4vfmIOk9QP/+cMrNiLBYHK/bUjgTcHyDDT890L0o/Zao
4alUqqz60DkIzy9HRM932TpWyeNYIz0p5v7U7vhw7I8IanDbv5RLIn9Y8GMIlgFl
KshvbNBN0tlpRtEmsLrTPR2boTngqaGJtAOq+ZclxbJaQmdagrKmjIgoYK9MGHE5
vcKq5dXncUe46YPo/L1aMHGwpXMzm4SnScWSdDO+7nI3vkUmCY094KwZaYrum5zs
wH9fn4MsvZM43cqE478V85Eosy3oyUQT+ViKoDAOK/2tP/Bf7YgXkTjKungW0RsL
3oFayuPbwQwIh5Woz+2B/ZJn5KkYwivPf30xNNCp74ms7hf09nxor4gOBEIoWglU
ML0ak0zYeNQHsVaFxw/3nFEOE7iLljImIKJhg9fteLF2RFqxMJ2qV2dChBJ1i6da
OMwN9bafKYvKvpbFYE+m2VqFUyi3IznvJ8GfDjeMVt1N3fn0FRnI1yLivYBA1OgC
v8EWk+DrjYpn2Dc0jvmQRTdYa1CBX9SawzCHj4nWipKvYP/6grQ2jUpw4RaFKDSY
zvD/W9/BgCtPtuMI9TVzuxbYnNivVSx/nwcIePxWy/fwFGIE2xatByghQl1Y1Kkp
hbRBueF7UUsdcbYEgGtF4Yq2im02SbXlyOTSezs9kBCIO4G+OnYaWTaPreXffQYz
RJU6S3dxEg7odzkisYqmgolqZq2AHA022OvlBNM8VBPxzkVTkb7UQ+Vw6ZAKqce9
GMbr1vkU3WMCuqrTEmofBzjQuS6SFNPVp/KYLQ3dUVqxIzPWY/a/sRVAkG/8+hAC
SGlv9eo2aHpjwgS/laYbKeDSYKfHT/qNLM5Qlkc29P9KmsGafZQRJjlnQqBjPl4o
iugCYuJTZdLVe7J/9n+dQdrnRc4e6Q1EM4nlCKKTxYhqixnyXBwQGttgiCAyaxi6
9RfsGGjypIEUnc2S2ReoDbU6yMiPmgvPT41bMYpHFzQSPyhPq5FarAB8XcL9eATy
oBIYe5XIZvgmI/P5EVqXarDTluHDxOL8T8egjETUmuZzjQ7a9uMKNBcoI1CZixUD
6w/e+iriDPqx4jHwG0sSkfHAEq93hCQxYqR3pv0rQIu0ajbT3LRM5wjR3E7W+Ty+
wddEZWLJglNQgXI4ZQefAmueqGau2trkgaV859MovF+UlRJOXZpcXCGeCxMKdnr9
R9JMzVuP1E9y0pb03ax1U5MReZV2q8vrRTk8L0i9FDj7c055iJN5+HtItH1ZVoWr
d39NqmjMJE53Iuy8FMZWGaftsM6GxnEU5xpDk6eLixV7mr7qgw5SFVYz2YmWXx3c
+/S0Cg68mEham0FhBzpnRtslAlfSCQVbdHiBjr7Dqsxk4/7W+zgePkL6sgjNSKZv
xrWAnaW+z+R2LvaSTdalXXXb4klpO+AQZ3aU8TXr1d2+vpS9fqvfr9Qn5nUYrvLs
P3OWQczv2p1+YoNAbjlBaDXzy2tyD0xPSdRCJmXwcFnhgJBlNCdt1+zkpy+lIKBU
Dg5TdxuzsoutIGmH61+M5Y2rZ49Lvsx/Gt6NPyHQeOYkJiyftge6aS9Nd3S9uLbL
/6AcdRFfbG+aI5gtyWvI4ukLAsYelgMhIP59k2O3pLQNUj0WULY31//5CkeFaDB+
ift0r6uJ9AKsQClY0JULMXYW07GXvlF4lFHrl8thFl11QTRO1aIntXwhv3CocDh4
5jjUkzwMVi9tDyj2VUrl9k0Z2NHS6P2pcc4C61shFtjhAeijIvgnd9v3nJX/hb8T
xYacG9VrunEayw/V4ItbYcb07SGHcukX5RMiyNSkcOWixVkHprbVlWjoISTpxtuC
qOyoGLBvoTmQyAD45o5eqetHk3BbgL9qqWpas25ceI/bEVpua09A9EHASPyoUnA7
qgG5zjjJm1XZXvIjRIAeSXpnlc++nJErFLnXHDuqAjCtFx7wBhCK9hJ3i1bSU8qp
ip0a/Vm/4nRpsvxa5gQX/cszLqzCuM6qfhiNwKM7HJDvogy/rZRUeyDI6+ZdANqI
kHUc/4xdChsZILdYnkSDfhCt7XMdDFm4188T9DinrhOrPxFRtY8PwbdSoxXh7Nr7
WaoHhdael24hNyS3fAl0g0aCg+AW/s0a5WDLwy5Zhv+eWfMvssqg/1RjYf5yiuJq
0Uspch9O2qxaH2k4+fDtInA/uBCjg7BRr5uGpsuma6qv1/x4/JPSDLmFZGXjnJs5
Bl4tWfBPzXa1UI0coBf8DX4cgzz/U5OyqSlKUp0WvjmRP8r/Rfv9wQZ9EllCrikg
bsAmM10qHLeoGJoJSFwtDdsfIse8Zi1gN4p90sYjfgYXvmxOzrWGaxy6RY3gWwvS
u3pXJekrxHwla2dA/+PyPwGZA/EXKgT/F0IyAv1rPDyww+yLA+qe9QtigbGHd4to
yrCCXm1LS9HswVRBV/hMKISCDaYEWDwDN/e4SAcB2lMh4v5R2je77NHNBF6vmzy3
lyR7ZSUkpBAjLWvzEhi3lbEiQsKl8Aq3fq2c/wBLIPNUX0N2v7A2eL+gl2BqACCA
PIZmCCksXdTtia3xW7Uv892kg68wWSYmp3ffmycsG+VIykHC1veWnnQqsEqw2kHw
ciskELJEJrRA0MAuSkIgL9r3V/i0fFndduRi1z/pLeHXenI88k7FLCUjVe6PRObM
MuA8kyUfqxtFdHI7GTrozT+4A2m7ljovA48srHXWXI4c9hoSipCM2I8CdUf7HDSN
VmjQgb6HL0e3Y9XH5fVICQwSJmvKtPhWaO298B9hvl4OCbWZkhTYCelPClc+N2K9
as7joDZb2DZ23eEGT60ibDVodaOzvWqYfk8pSoLUsiM0SPUnYbh7ROyjNAFwL/tZ
j4aKnCV6wPC++hjuTOQkJADtJEOmOJwu79Wn37ZU0fUKLdYpAuDmNCukmVBi0sQh
4eygwrNmUYQvR6qm6uY+Jb9lb4ZcdhMkhIb1Kb94ZalXl9L30t+gmkvWaM3YkC7I
JP+/DBgO6YRTPq1jVcum6Y7kJb88TstC1zs0MDC6U9KLfsjEo+dIHZJnEtV4St4i
IRQq4CpJ9vV4r0IvxYwZNHZSbxSjTmNLtav5GBpgC7Z8Gv6X2iT4TF5K+dU4LvNJ
vp/i0q971hZU6eRhhWtIe+eAZGYi3WsIwqBpCil46zeEvAJl+Cbeje1gUXFx/0A6
wTr9uP2QiGS5BHOgy0149D8qUbBCq4IE/dRQVjBovmJkCVmW2YZrUUA9VpiJYRHt
SWM1bd62zCA4CBngBu6UNMie0p1NgDLkME5kXXS4OINkZuY/jgg9zZznTwo4whrv
G2HvRqKc8+dWcIcHtmJboxfR6KWyk81xqAcLuy8ktsZLfYZAbcgII73ZAiUC6b/a
AE53y4Ul53OYfXw1Gi+uxzqgY+n0hLJYoiheZmDX6O9NrTxsY9O9FHfxxkxowjWk
UTNNOoX41MS4NQzCaPKIVAPIwO0AOyW6HhWmc3DNDRiCjN+z+u4wCJNuNZyWhyei
apYuB1aPQ/gfl/0LWJofq+7sPFu7u1rt/WlRiAo5yC+kgZa/+iwKeKadWgKfDQmQ
/mYDPWBR5bxg75IydNUHoDkREqyBPpZ4+AeN8hdoqh6NAs+bwPloCo8fWEMmhVce
k0LSMuch+LmNmQhpcBV4nnsCBlBH25JJhTFzIu36I2yxmg4KO3iyFmN/7+LAvqmx
nXSjMN5tpDsARmLsxEdiwSY7q2pAY/jNwRPGKoT6fgWlFtHRfLnyT5CTscdQvNKV
W+LZcSS2SwILJy2a5SU9WDVkjTqcDA3aO60CaDn3k1T0mjM6iuTloFDR6h0rmi80
cTTH8hHCTCalDLWIFC2JNRSOK8m0CcsKZbMMjLHD2FlL/rkzrX7KKlcl7UxOx50T
THxKEsK21NmexGBxSSP8Y33PzWSsMEYuTznTwaaXSdx+Nlwe6QTNRemFCKHbv2DX
3lGidW5EKamG1B3pzNIgknwcj+bhyrIeMQYB8L5IW1L282/E1Yf+8fkdWQLz0c0t
0xDAUfUJZ1u6qQzPf5HYXforNicZoWVjbNqZaT/n8sbM7F4omIpLTyBmCwQQKhcC
RAioULlBwxZnPeD9HWG6cJpeQ9mn5S01PbsjpNI7NeSE758kc35taSnK8EZc5hD6
EVxKLa5h4qoTlVHflCkj2vvK6GRHIXZXMMenuXpnz7mw1kOpBg36ydbxfbUGXpb2
PsaTp0QOPVukUssxbjcJrRNOvZVHcV1555CyiysLyjH46VMxLtS+gc0lnG5VMXh8
2rvQGLGZ3/N8sZRCQZl5vdKsMaEYUyvMjxSZ37Dq7xyiMY+Bp33LIKyuyFcjT+jp
3EjJwYsu4RY9gcJkidZGVX2sJKASvoogXg7jPOVhZcSZtNOxpiO47n8tpj9N5T9U
KgpuoxXMGOLBh9EjrP1yp8b4rlnlcq9aMnmDZtfxkwjh9tLlX4H8kR16mNtmFim+
dC0+uOYbSAzbNW7qXCWovTmZXeSRDLgmpXS6t5Y5WA8pnMHWMhUqqGvn0E1oFmsf
1xuB3BUA+TLVOJQselssfI11hg5WxK3hfsGuGvY1MKVuRL1tC3wpBtSqU65XLO+Q
49web071nCtqV9Pa8Garu2ica8ShyorE9bf03BJLJ6/Ox/7MYayeXdBH+Ma1lxbS
Nt186cGh2RFve7qqC4koSfG4mKXpjERTa1IBiJhsSxgcxEYXmZBHdjhp8e7Bq7r1
wZrMqePa+wyZVtPgeW34KQdcauaQzclnsEZ1iXO77lhq+2HDz9Zzbc7EHM1TPBLX
3eWsA5xCkNxzFSFedOV7m3Kmld2xSmT28oK7Qt4yQqpFVZljFomrNyVuXnSeH1Oh
DCV1b0J8oY4m73rj/WW3oOowNxRlWqAM6Gb7pUxdywISmgiNKB6s5ae6QVkos9Pz
TAw58QrjIvMJggyWONox12XBFQ2/FvrHR0xrUZbN3Hpml9L0YOFQ84z79vCufjYX
5zvnuS0kPAYhnY662AVebHPMlikjO+06berQqggbxDG6fyC1LGsxu0z4pjTO2Uzn
aunU88gOyNOW7cQOC5FXfa2K+z5o+s4fwLYi4zJOuBsSwbzYAvECEqTzHhUsqLKL
3RuWEyIOuK7UHy/I7nC+cLkWGBe63cY8I0VsX5monxqLt4nF6TzAfh/uQPR80U+4
XgqbghZZ1yJPwImRn8CogjGOXoK3AEZ1HfMYoHCdepsXtNAX+kt8S5CavomPRbzy
5IBHl/pKFvl4vkE2ROjuKP7BIoXch7TOPoUHkb3EmKJhNNcbUPUNa4lz7wkKIHGS
qOtSqmO0HvhmOtwBorRdY42Vf8D+4pGryzvCOzJc9Sl7xLiPNDiZ2oprY5FFRDaa
9SrYqBNLeVapSMANuK/Mv/MQniZDTQbHbRKZMGyatEdtrHMnE38174jy5tKPz4dA
5oBjltlIJ7nT4Q0vAzfepKvdoTQL11j5hwmOX8QvFGfWGUCrIhwsqp77cH9AOoXb
IarYQzeoVbizs1j2NgOC1FsLcJy7eksUBeIuiC6tbbbK9sRb37b1IR0AxU/C/qB1
kGzAvxeqg4YA0QYNYHTHED4lPMFrK4VfV91Emo27gVN9NX3Ada6abgC28knCEqfq
UD/S2UpAcM92Qv4h7P2Zan3QPGkbxjovkIpXvzdEbIpJsru/iDfH4Lpf6qs9+7kX
dt/9IOnZHefjtoyGfJ/NzjFFYWdujPSbWcbINXSTbDKOa91Tyr75LMeitz1dWjNJ
bj3dv/IzXZpM+A6XS5mEUOy3N3ODehXhhC79yyfkHh1WgOAkC5FXVEhhpiL/W+5P
D3+cpcQ+iE6HXSeRxRAA7QgeyHn0kvfFC3lr7FL7CSJMTZ2wom7BJeSaDghBtzi2
Rt4LWGxEgz1hY6PE9V9IemlCyU7k3W7SbuI+XbyA4UG81TQ5mEjKrSJsKV+74T64
b2/dXFMlUaBRNEXQRo1i8hwDb6cEIdF4WUyg2tC1LPnuMDjEKnnldLRMI3Nqi6/O
FFY42tNjYi8B61N4OeF5NWxm5z9hMkJhVZZjvszGpbjC11WY+mUcAbS1CzUvdFmG
06OQGg6UmoEbMxqjPXPig14gGJZo1PwrvARvmQ+lW45S8GtDGny5mKfqPNGeQEl6
QiW3+NRe0D7VuSrvNmrkxGlZS8Za5qB0ghyoGCNIWb14G1yecnfwIhsW0a6uqgW0
ux1RWHEB+UN0g5QFySjkHx3y+5Ps1RkUJ2eQUDurAEtG9+ZVtTumpk1QxE43YYY/
WTR9NX4r9HlRbchWFeaTaXuadM5iLXpRHVYwi14fbch6CVMk8LeQQrW/DQei8B7F
NMTmJNJ58OfDv9cfRSjWTKtWkNv0+w6lABM+4oEd6xGPm/6Wbk7iDMmbvNy0dwWB
0gV+i28U/W7wau8/IAOtkwUmgD09na5t/TP2QC4fGxwadOnJ+BakXqLWbqkEzhel
r6BuE0VZZSJVUbh4ZywuHZBWerOfp/RPL219pFX8yJRNrwOdlfmbMMPbm8FClQlz
YzARZHC/PupISolZW9qmUUVqikAjwAKWcOWewQusm+YUdovnZ6EjY9+6hL9bbjco
xOiOyGWmreOK6GVkW+wA+60HDTGKgDquhLFpIoRTGYmMNOZYXyiY4qqH6zn8oncd
eZhZJzOQbnoePFQianIowoJ1mo1jXBubF5pinsJiwdkIeA/a785x3AjwryJsmbbL
uHdqz3BnqtKdi5DqrkuyXacbM8JAB73YZU675m8/pC1PuilBkXlcPUIc/7TRBsAY
0ODIfxZcX8K92AJisY0u0+f8O1sDeCNv30wAiEeJsStuGduwfuvW/fRslWvR7WY+
wUEpRdnd/vPvXmZiISFt7yb3Pl8DVVqUcKpqVLJKbMwreZA6U9ymUu498eMX/zaT
6SYlPaUzdePPWyYRG6kHScRCs+w4UV1o9Yef6iIey4eP57fD7OEbqEv/dzp+/Ywu
p6FUUsnCBm2ipU8OuFy7L6w5V2c8ZoMP7yZ/Q6WhxdRwkygKzNFFVnNXj9r4N76O
fOEwqTDb95mU6TOxPckcPUDWRURps02uT2d+TF3FPEgXRfnZKleXn0Xx8vxKGU8v
V5jnKCY2gU/mOG87Ijwvo0kSztKU+RYy1kdokjpcSJ7FphS1aJDTAiCD9ZEqS566
fOSNUu3W95X5YNS4CabjB36hHKIUwAUGuHQ8/MNEIqdM5AEkusM4iSPYi6s52636
OfLOtqQLQf0/oXuZwwryjiWRVjx0ezJGjLluRcwe9sVnsilJmOkv6puKTAJzT+jl
2sHDQpjG3jrWV7I0b6nYMX7Lus2dC+OPhG7Z9epbyqVCyVND8tbei57L8Rzh3q0/
ux/d+oXkW5lxfmqe87zhpFAVg4JRtFMn7swRcHv7111LSWIX1SmxhQQ3XKbpjjmf
PZdOlz63KTbRInr+B8AbxXGIzioWOJ2192KXdvAlf1eJEBY/MRYubykLlYCA4CeE
uuPZ+RMg/HHwhbGh28NHHwj8mCzL17GKHw7VYGJ6KosBKmnOos/Y/Vy90hLWHlJ+
7G2+4J/KV3806J1SlZFcathasL3s7cglrj7RGX4+HJNDhfNBRfFVVnhTGSvUUpd6
9OZMkIvpUzpcQEpbGahZL1f7yWLQ639rR6D3T2XehFWhffCwAPu6L/UdlyRqzo2Q
UlTMxqOa87tBfi59etVsRrK1Ch9tpIeC4E0fd44XOu2m8QF5bMVuoA3hZyx7HCqD
AMCXXdKfEBolfaqypiyUlMkrkhHdsaevZgXAYwb64G7b/MbrhEspDYrfGrwoArjR
u92ChDYRCwty3Unwwl+J0dXL5AV0TJEkF9Oz19m+ABx/xfEdc7420NMEMBkgHbsp
7AQKtR3qIoyq18vVBy2SRPd/WZDzG7lcYdn9oJNOz2jb7F93FXLgYUDPfOznUh61
vQc5/RCSH9cFJweHQteWR5xnYDSVsAoSb0yJ1e9JVBWOCH6DDP7YHsCzQthQsHr8
RQNMwA9+Qq1Bj6OPgsmbGzdufCS4BTvdMO7uancqAfaC+Yi/k8wUyRkskLk4Iwz2
lOGkk1hr5ze99lqtIECfh3vlpw1ILlw4zz94WILyiSAD4TmjmiGw24vD+7FtBMB5
5eIOgoxppHIff7BHYlazd1Zpv4ifIV0JCRKP0Mk2IewBOveAzp4Wlg/BuUbu5wKN
moshQwhROECFdEbHGcdSsZ2v/UQVY4RdTu1Yg9IaHY9snHp3F3lr+rkS0s/8rF3A
N3hRqsaxxOd0q63+332VXvnAxWmAriTgsIzDoEEVmKdPY0z5NlaaY1W8ep5v0IjC
Zc/cbQCEmqFkW/GzTjmS3jw89QvQlsXYVpBu2GkVYmu2HWheiUrUikOObTld50L8
Q5nCmKu5GPY4FoSlLrjtxDo3jXS2fkM3gQboU++ziZnd+9g+NyriZrXgvzNUKe3C
0iKnOFyp6Lw5QlIwYhxgEh1p0RAjbpeBuDs5k17zbDx9t7U8BeDSm1dwKS0kEeTI
t+WtJO5yMnXXLSzbsuWbLz8KZhHOemFSuAqkA3Sjb5TmWfuho5cc/Z3Jvf6iGpOl
NFNi1TIEDKuQv5EEh6y1oqGpJOp5fpXPgF2ZyenXUSdsG+BJEUXmd/NEKhvqi0GD
9M6AQojpVGi3S8wWXBm20UQy6uDNgH0zHR98KUAEb4QiFQ3tbEFFGtBqxNFxVm9W
SLGZYT8B+xwQEeB2f8JzSn+ovpazy0cz6P8IVlppBa8TNOJbCTON3/CoNKrwJbal
i8yS88fKzwtixDCdOZpHfoXKLjLcO4ZlnD0qM4hsTsiSbnkV29l8umDDiRkhXHu8
VmOXG2Z7y4Ensv4pDyPCfXxeKXhpJHihBwcZCNo2dZNI0BtB9d2dCKgMA5jIm/xj
IHfSvUwoXpZEBlmX0wpKR4oLkzj/RMc5dUUV4LvCAerxWLR85s8G2pluzeF3ZLnr
GiVTdnE83UJVvqJxFtkjX4nqciyBQN/QhPMF8listl/P51CtxDx624nQ/FEhvLXj
gBCGmJki21L11NqzSOng1DOfVcCUSWx0GM36Wwm5VxEpqriFiJTXyk8OVFPhndAE
+2VdSt0+92mVAql1unIfaPCC8hEjVB1IT4dkT18K14MfNxUgSf8IQqMC2F4m/LgG
styVzq28o8DYSu4+F3JZC61iX1EOnGF22Q4NnrzT3MMJjwNlaebb3xHhJiq4mTGZ
v+x91JrNOXpJrA40UlBMfiFNJ1/NbXUKgbehBA2eZS5g6bMkI3SOMOCHa0YCFvaQ
vQleoOcYQv/O45g5RtDIw10WMwmUTqQ+LBY1WIeu3UpRWuLcxrAmFQtqlW9duJGb
ZXucb/lwT3BeTYWp+9Watsw6RkVM4CFHQ8L7GNdhI0XrRti4kQw4W1xKCP5JGw0T
syxvVWAmNQbq4+a0z920hIQm+a1Os7q7P7dSWfF5fRD++o+gBxC2Yr5BPbBaCoV4
GAuBH5sfOU3FU495OYGpj3fta26V1gQNW9+xIE+Jabz0evaL5EcE4RSDJ9vE8wL/
ZBz8+Ntnm6j3E1fdBG8NmCY04P+/ZhsOfKNRypZLh4y8v3cj0YEFsgqVmd9oGDA8
fiLW4Dn27w7R6fK56SauAKhU5D4VQ5n/OaQSobnh+ospjYPIMTR6ryE2cp2ljrPI
Jn4gqLLKPGegGc0Wp2IifaU/Y6z4oPSdzFY0OG0uChSXjHV9uHnr1EIY1l8bvvx8
12LVwZkbO1oqVzpuHNm4yStxYUduOCsHFnz/Fzxdzst6+JFgVo0UbNe0/FYTbgdx
jqnTIXwlmfa4FTscPSgX0kEVdMzB4T6N2LUa2QVr8fodLG2bTXgklouos6KcztA0
byo9lM9izudII/jgzKoKLEnTL/kcKJwIpeB2jUD0Zd/3NBSoxIXoSsJLn4hy1T6I
KjV40hc9m+4NwHG+gfdHuNOFPTvTN3et10AriTNm6v8p33IBZZvrT4mmrlPJ8fRM
RcU52swh8eqJz2q09PzcUK/65s6RUKxIbhaQv5xp86Mw0I9P8zdk48exJE4RLlwN
bWGk1JAMklahoVFa+nMqVz0ohNF5A4mtwv6utXE6qeg/xlonOhovODSqI9At1Bab
DsJlugQZr5lmrjSA+uKR4iJakyDPsLA/Cq4NPQZP6zfiy+r3/9S9o3qeaRRzZ/Ky
1Pkbcc5Nd3hETPqb8uU7SUa3QXM0lRe/SyryZ+htTfJTsrhCVDbGBDAG0Sf96QTs
myhD9eSCy9f1v2VyUPdGb2XPM+ZYnvXm/mSYuNU77fh+vcQHCVOBMiA8IYTi30TZ
YVoQrSgOY7Tq2/T+9Q7Cd2Fgn+nUxPDpwBPTbL5uxwGpbAwBpGqNRwHNXYgqBkj0
HBdkAt9W72xIutRH5xiF6uBKAZA3l7WMmTNw1ekQXcH1i0+PrmnPFExxJkyTcXw9
4NPxZ3X8FBJeorS1gVMSW5+NcKd8SLZkyPy8WMyDF+/lFZQOrTkBT1uk6QAozKM+
15BCRlSzHj5J+5KoC+YiRegTthTrhH3juKWWXmN/56BcWw/Jpz3WqY2KBmXXTRz2
bmejFEK4QK29771bto7QZbcOL7pKj/xseIFXlQbMEyKfMChrh2no8VnTBYSO4uks
7bs9EdA6eJPOwXAexf/5KlzqN7VEA0D8sxGL+lZpPgZO2b1UdtyxcmDZy+krClNA
TnYv0mX3T+qjQeRCgfMzQrFGXt1C/h0OimnVQvKaYEoAQFoFEaqxBSWAFqHYB44f
/FRp8HZYVJtKKrbcwkO6KkGouxboYpXRblsnTWZsI0x8XnKGWD85uP2+7rAjEFv5
Vp7M+ouX44fT0PZJrprr5VoTap5ZasBcJanATbaGzmA5inR4f1nzn9Kw4/yPLVn4
fYtM/1yCZw8fpOaxIUFcJ3n5TnmFnhyqv9NFGzSBnNpvM/flonf2imtX2TjokLJI
xIdyoh1BU9HhEhEuhI/v486FjGyVdADsJbt81+SGa2Gh3XFKMFwwK+gZLGMa0iN1
WNS4PlkEF7pk5niv3IzgUxy9X4SOk35/BKUeqmPqPQWoRdhIdDbizGh+X7TWFkO6
JCpUBtwxNmnAnvzgcK4JGsor24raurKjY74P8HgoRBwopHz4oDkU1yWkwDpXwTeK
43H1xIZ0qrHHhleTbFO30chaMkUovEk6xLI4srcRVTTXjeKus394wCmKs84P+AN+
e2OXIZC9tiuzFIqiWiy/Pqr4NGmr64klFsp2ELEq8diGSEpbjXy7u6yX4yZh0lwn
OfUesGgtpQOgqx0fN7BooZYurrtnbELaHAmPn+EWNDcfK/S4tyQpgRToFBXPypAG
ma97hhcvdm7uLpuEHBLtGMokLef46HanWNH1MDM4zyR0wkyhbjXehuiS8cnpzUwS
ns1I4sah4ZgUHP1BB3qqdB60c2MhxOUs3WWAruS2YiD0znP5PLTSol3LTHDYpj8L
Pz29oAAMLwEqDLY/oD+P9CmHpcpS9eP1U2R2Z3rBB3UzNXiFwRFdERdICOyE7SNq
PGSDQBpYXLM/oFCmFvmQeicK7Nl/e3F3S/IAV297j2ZzdQo8K1l2jcWq5t0FTSO5
vyMEZlr2xzdSt2b69ZIDAzu6ErhVEpxos6LyJ1R2kahXwBl1cmp7WXzsFDiR8Vqf
i3Iv29B0i0yWv26AfRZnZXcCu3H4I+L3g8YQCKAr1Mu9Hdv6VuIN4DqKIlGvW0VC
VKioO9Za24fz70ONmJbLuf4G2nxValYSpmZFPuVwLM2sgTneWPvOjP/jMYw0nV22
14Gdy802v5HO3gEjpLwbGbkyRYuS+RZVUu0ZJPQWVPzVCxsqbQzfHMUx2R+WR0wq
VGpX7bJ8qZxlKLPYC9nyj2SXX+fgd5HwgFsu1OVOMk/01QuhU4ubBImroba9wynJ
CCnDmIGIlPZv6n1PGodpYAFykWn86t0ZoKVkcVHqg3cuPy22D/s52F1qkfGluEns
3CURcOGTVkueSdj46w9Etb3fQQh1JLKcfSGtjR1Q6Tp0KgOpqOywcUoSbvc0p+qI
l/oP/wjystPlAK2FsaROztaVA3E4X8Xo7A2iWM6zV4XUZ974g96ChlVv+IYOycoF
MoIAl9qrfJGbmW7nb8kXFqDt//dDWY0n2TEeSVoYyL+z+J1W/+lHICWbuvoG6CZq
C2ykguJ263zk9BBmXEP18HGPjl4LsOAYlz+PzxFTjeDh+iL1nt409uBlWqCNwPAm
gy3yqhpqTqrvAlvDhSbRctCA+mgGU2f1YeMdvbbxzuivthFi+CVHDW8NZ9xouGJy
qd3wS2+ZV6RsRuBqfHKYjuPiuKH80pD48Py1yVM937mTdVTaf4AioWAHIGOkK6+f
39PazV9609ielD6CamYf+sD8cjlPt8pIkZVkfDAuoKmbSE2aCWkyKLoG7farzLYU
eQscpXY1sREh2lU6L7UiOprxSaQN0eGJ6Np3Je4OFZvEWD6TiwWCYfRT4vy5eHea
7K0Icj+HDKK8i6ZJMB9sBZ0mllIglj8zlrg0vNjwgMZ17LTFGUQeFlMNw006FQLb
h3DLfyvaPO1Qg9GaQOPPBKVdNivuorkfa1gd5Dvhn8hdNEKMTI+8+KWitEeTjb60
bGtTKZd4Jpx8CEsb/iXCpyo2BGrM4gn0gfMutpgKfFHHnGHWm+TzRGIcAXCl1Aie
GjiVWeeNL8W9lPL0igK3Jcom+Ns4rLrbmx5UG84nwJ8xpEPg4BR7MSMgPBmzQ+Dx
QzZrZQUvqEvdScISHHasXGp1BP3SXvBxBS01v9MFUwfWiUdtbP7wM83/z9yNht94
SrnzEw+Q5JkCGBYrzHHbxeJEf5/JyrF+x2KGiMFGVOv+qWuUX7Nix0VXoAoPu42d
Qh9XdpD6rOlFU04q+4oFrAUxRZp43LxDSDT14y+7GlB+raGZsfAibG7AyU+MPvuk
gZZC4jXpf23naHOL2Trk1UAuCPV/Y9MsH9RGljN4jKUS8WFchSv+KiSCCTySA3RX
rasStKkfWQ3csaxjKgjtykeaqfjv7aqT6myzHLR0yl2L4r84fIFHVA2jY+LZ6DoC
zfetzYqzSngWGZRA9MXDpniKgipqIubpEH+ZLmI72eVplgOVWlUBz3ay2ENKxMum
SDplUwOo/1fWlhIXaFjMZPQX6/m1rcCb0CSe9h7YG/wdQaEyoYMaZ+W1d3+lQd+Z
ZNhoo+WxK7o3JVZbjmwD6jAg5V/akDX50C8H1D063t9589RedtPYaW0G0p5hsOKK
k4UPM0l9lVqzmT4QKQpuEs5Z6S/QKIs8JS3ZkLnY5IM6gvXV/tnjRMB+dWnOjeLQ
TArrj3iCBEPMLVl4tiUn8AHU0CvH/158mXo9lPjyGUxn/CnIigX6GAhGSvLlqADu
mAybJ8+ZQwrVh6O6bZZOVhPLew2gjRF9DABF3k8pm5dZrFBMu/Gz9aP7GSxtV/ML
cNEN41MmvUTWN4p+1SURVkNeoJqHUxbd8brrcxG/iXV72Lmkb2SNA9lQcDKhF9eA
ysvrLGOAfNQrc6skLUQj9bfzUvbzNeGxIEZ1NB+0N7TXBCxjm82mdOm7vPFk+Bwj
kNY8trnLMiJ90Z/0PUmJ369aMCctiMj9PZY4/wf3K6srPA85Rpdwj+YKxVkYH07p
Jb0gABOw9+q7BUU42ShmbkwSvkAwiYNDd8iaAQCfhBGGAn2bamO6yjXqVK3XaBQe
YMCzif74Xi2bqKKzXrwcIuDsdErg243j9VWnf9ESMp3HYr/yhOf1cT86X+kqv72f
fcJ/e0ANAakx8gyvNHJUKomIfG/aS/lO5iFhBXgG+9OZlWMnLEnz5IxQrHZ3M6Id
t1Ho+YDYDnx3siG/80pK7m9pbj/KziCcaUeRXWeGW0Ki/3MDjYab97yMXHSYrN1U
nEFN7ZyZzaU7aMV2mLXsgz0f18jevmy7gMxk/s9H9vLMgDhvYew2bN0h9ar5RRMc
m/hsBotPGxLMAGDvNhq3JUt1tiswd5XA5qM8We9mg+lt8zp0Fsca7mMvX9p5qbQU
OpHu1byfxlZlZVN95920meM9lN6cnxjHiaqdDM1sk8R8z/XGJXBZ2/qehMNxlPjM
UMNt6RwCAl5SZM3hmSatcoG/byQ1XXlPpO5U/0QybcvhyQsEb3eHnrbIYHTbib8C
guqps5EMf0FDpbkX34xrwoQKGrDZESFclF4nafy8fUbrTkEKZIeip+EUK1bkANya
qGecNWZYPwew8NajafvSQ+yiCV1ybOI67RzZ36ESbzjCRlKSkk9Hh3RrW2AafCyO
xquLw6ksJw/7c5TI65HlRAwmGcFq6XfCBVlYwBBhPfCIj9a/5FzYJP6NbYZRZOvh
6ARimVt2MwkUmz8uA8UKzS8cVfgC34WiXjL1GGFQhSHUz8SS5e+gb0YiozDSx0AW
Y5SSKjB9aIvvWx8ZObBksHK7+QuiJY7PbgHjb3B8sg52NRaRKl6SuwR6I/ltrVMp
qCAq5YjKi/MP2jO97OTYui36+7qyULD4q5tmLfZCGA/toLVhkLyTVn4rj/1CGGF6
84MyuzEIfvT+kvqlTSh/CiSRthRHtX7FvRsr39/GWN3CMOdvOme636osJk3UElcM
ljqDigT5GQ0IuDPhrNI0eAvIHVtCTZqDRMa2/7QPxN3D4eN3ia//3fhARdsiI+RN
BwSjRzEAeuEJtWeahqI50Lug7S/LGlhOyq07o8r+gqZgBnRGe64qqj9pfX+PsWlJ
gHWOtq4nTRmf70u/H+xDZUeJ0yd76xH34v2otFAaVTDt/V8GjiRAQco8izgcv6Cv
oIHz1+VbRUFBaMZPhJ0qFyD91HT+OLPDPkijpY8dEc+mLlgyYm5uRGr2e4dZLzKy
21m3czJYnQP2FcymND7qRtyVqrGzejMGK5feIFYx0Cue0X/TzJISrXgmhf2dT4Vg
fqCai+MxXVztT7EthVu7/C+z3cJmqeaDnswhrGonqn2SevqwwOMUHaeNptBqYSo8
SoCjYVPjR5IHw0SCbq4J0AUzC4lBq7WAVkKo1+xI4P4uTYLwJLFRbugoUtlN0qK4
/qHusHd1eGtr1Vasl4brEhv8ZgpYU0bOEFo4J6Yk1sxtb30jlOkqD7Btac9nWOCh
NwOcBYUsFdeZsa28KOeDcgaIETxUxZgsAcPA36jXyvbtkcWUNRYC5/KrttKJ0jQN
FERYENPo7rkkhpqn57sWM3Tbm2ViMeAB2ONX+4WeERt9NMCUC+tWLoo0l+0gPckY
kNVogfnEnGUTH3F2yLwWiW4iYlrRmVE8XIoxhFWBD8cO8/qfsVeUonJUuA6VqoLt
Dzw4HQoOkoZ+pSAUXAIxC9wkXEWaaVPu+LeuCZLVYM4DQQqVYpnqD0Y48pjsFTmZ
c07gWobHnCjn0CTUewybF8IcwsfFoWBvvTmicDLrGbQyHcjQxijNCowdVOZaL2cJ
SGPrz9HqhO9kh1nZCgi8SWZNDQDLsfoxMRmBPBgaJvEbsgK7Vc5dK/CSAgg7yja6
kCiA+mK/ByFzUwN4uXN1/BpM0mviE9mhuHldpPMCxZWQMpZlb2ttJx2tXfcgkkuG
NTloeNNaoj0ATIW9EN6V0uNmEi2gva14ZXIm9Rqsv0eRQg3Ftq/ucgUDBiJnu6Yq
OuNRXVAEhomnEchaxYoOAyPO2nLh/Q+qPeKJ88DxBi8EdCggBzrEMQhWWeqi37QT
qKYSUh+rljcA0YTUo5Ps9/+gRL21i7SpF1jy0vKnucla/qwRrMgXqsNArHzolaZC
5OAhvm74YkOVu6eCJyAwGOWWDFI29ae06xBUsqHOIcErDH876XgKRl2lvjl2iGOF
LL9bRqVFke4Dbx9fZHsTVWhZjyslRsW6ska2tR3ednQuIYxvVajnDgPMWNfOH5FM
TqkVlnPNy9suj3L0w5F6TJF9REzXbAX5BeAw/lg0SNXwlEFb3dRBggqj4BciaRiW
T1eFXEBU9uZ8CTpr9YikQItdwEGhP3yR1yOOCNbjW2kjmmS88aAt6mMcbjD2rERc
fW5UtecSJEbJHl5DI5XXeWi/6rsm14SWzR6YlP2TSgsR2C//ebx204Jnzy+wNxQu
4t3xXWt/dxlGeiQIwsejpSwhsgmJDscWXKn9VpLhOMXZjZRrvTW3F6KAgR5wMnZ7
CR7DqNf+XJGLmwADcu4p0utof4OfO5BuQefs3TS3DVk7Q04s3KwKLjnyhMVPXvGw
PjvejzJ055Elc/UV+eOceAl7PzJbLIIXho6qkZozud2SSCwdAUg7iJjwCd/wIMsu
lNlff4SF/QvTlhOec+8T/2nIg7PPpFiqmijW0W9xCkG93WhbeeBJuXqlh4Exh0Ni
WFxHlPxrluW/EPV7XybflxkD3lK4vhkyNiTYu7RT4pEo8qdwVcMV1QbAyMihDqZw
b6+f0Xu1Ke/59nt3u8GbR2jOH4535qfbUK+ng3gBpyTbRzZ5wrKpEJtLtzprdx58
RkiWmhFZCelRTtLVjAPpZP5XT758H9ApkXLg0x9LnV9/0qRQnQHyWm5+WsqsQjFp
88CKnLOgYuOYPoCpxACpnBMn8VcIL03FZWCT8zD6JbLCO5K5iLwl10CGwUymA4qM
G3tDaEvMvCaCgP8/cZgWkfdOgJpJZhsy3ZN5zqtnhbSucZuqwORNrYQL819dJkpm
uV2KZcvGBXy1x5VF/c9VpmdAn7EfSJy46la62MMZSXfbSS3YRrLZc6a/kodafhBd
YHr+eQllEl3d6AutAzwqaPm9NApbFD8r5rsAXiJAhBiNRU7BcaBCz++5MJeHZn24
lZ2C0et4evheWRhJw1mknDuaEYS82K97HriaAbEwTxM/Mc8SErH/L3liR2vkXual
A2Lg0p4OTsbj4PuW0G3L4HCrmi98nMalM8OBfZzjsmrzuTbjUS4YgwKD2MvpM1Pp
3/mZX70hB+3FxdX6VZWcXnTB+ByeT7GLGFOXIZzpgBD5Dzd0H9k4Nkv2yjj1/M1A
2eAWsjsRFfqML7mdyiImlAAjKROr9miZZUg9awiUl85FJ2MDazYnUwtzi5Gf4Z/D
r8BLgfcHkV76NB1d+Kc/ihfdJ3WNqLC7tPILE8Dgs4g/1psGx/dPdACx1F7l1aOj
4+DP1PP+1x4T9Y3Czv05J4kPmuwwIg2y9qxCzsAmE67YGHN2Yfw1CmJPGd5b0rmh
umzc7jiTxGKDoah1ObTLk19K5fCkGi4CCGR04ZwXvG9ajgoqvS+Vr6+eDLMkT0qW
5vjG2z4lr6OH8e7VKmsnpqT2di5Psg4P6B94U73ltRchgC11zt2bikJw+1jWzHSE
+1nkKCSJtoI4/nLChwBTUnUFS5N8pQZkoshm8f6CLcLdsS6qWvF1bLpHjaHAcqt6
9S/6KG9bswvSfy4nhDuTQGjWzSFXaa3xYRRdv/+FPlrQLmTFhgqe7dr3AwJYtkFr
NUwu398eVTAi0MW93+Bgf1XANMo+UFRjW3K9q1RCz+cH7ewhjVwOmgLAsg2QAVAU
DDtK8Z7WZrfU6lDM13aK2sa+zCS4oi2lb5RZ8d3fHkoBPC+fXfdOz9bITwITRreP
VKPyDq7X9L+/48stCTYWiXJmApEnxljRQlVYxGKUx3EReTLBWOw94wJCcSkVBmPO
CHWjkMQPliYlCAddu9BFfCaXqq9WZMsjZupXA6TyrGapbxVTyjI6Va6Og63LvCbu
h0EVWkVdtyooqeRfoPhIBEoRd0G4Nqo9LXGo8zrjxoqGpweOKtY+QLXhILEcjdSD
DGbwkolcfK+s0Y752MSQQTvU4ZK7UZGkpBN3WkaNNXOYlz6QArkgtgTdurVi7ojh
osDz8w5ehASXQBnm7/C5nu95AAidstRk308860n3JfDat60DnzoGL4/DNKddEjWy
Ptw2SKANcdVVgqSRqKdwlfGo9XFkIXtfdrLqC9+9UdUw7WI4aChL1x/Fy5ENGJgo
WZaXeL+gT0s8T+AIy41rt+tP25L/FGZXlijbZwtEqPmaDjEhRPW5zijCKER1Pfg2
Q7fG0HLwqXUpiXsEzpwu4gSHKFyfoRn9YBHBscRTnas/6DDHEqFZ0+IJlaZ/Ht+D
u9dNqS7zDcd67NuGJPuYRXMBqPqW8Ws/5Em/ZYUqVhWcPoZk63pG/QeagJ60ZfOi
i2SyxVF2N2gQ1lIkOw1rWXDqcF0AWPsQpugcQP3YcQuH3J+4thyfSO6WnVooGNpL
c4f6EBYW6nEpUpg1hVPaOySpvlG8+eWQnAOhnaMJeW4ICIhZEOlxYU2mgjsw3omP
SGS31vcO6B4i6jlSCYuZVltg3sRkgkbOdKo4tox+V7rlD4+09ck+nrlPC0ftPgDl
o6l9vbLFwyUEyYpRZeyeUcnoojxdiqB/KmBsrtYr573kysdYkn9AVXgeex+gEh3V
ty7EJ+W3N7s/tqYV2M6woljmJGm8k72WLOoefyCfPYYXd9nwkqCoWzG5NhfEGdaH
0Q7o1/63Btreh7NMnyv9ZrfZm9wwo0rsbFhz/u1Id3hDDFgZ+ZnrGC8YQ7t731CU
uClsbzM3XqL+ePc5De9mkP8Z62b5aI5z+NWGky/Hh2oTOOP3bk/J2Gvae1FYdlv+
Y/RGXK1zrqEFvyVuJQV4fOAYMfO4ciGtq6E9acQ+QfOBDBSe23KBVCsaAQiqzPAi
tFGbrA5rbyokR4hlPwZZ7jNYfeKMR4p7iEi6FvPmxm+iyenR3xyzWHiKnw6YVO9M
f99rvYxLhSUktjiEfZuSbIhChkkR/qmSh3jzn8tzv3S+GkudwC+/DbAjsNCmg7Fu
yRSolKvBYE+as+Ocblm7asYatJ3RfVWoVr/ahOzjXnnWbg5J6NshuCk21gGI4lxk
yez8ua5RS2iMR1dmi3Xk55Z3apIxftAFMl6uPNgEsvIrGWbTjnoFH8JdJpYSffiU
LQk5gLocOcTd5D3cbmFyL9dckY/kk9ymoA9r7dl0BAPx9jjNvZrIsWFJG/O4gXFj
kHuaIHYYfO+vtlv11GAj0PcyDVFQzXHjLATL2R3XkGP/YD7RrMkaf6d763OEf2+2
h6Zgn4aDTNrS8EwHppsibT+KeZCjv9hV6A8dyASh8tjcFAoYhaRwWj3XgFNUprvF
XYVGAcVzx8HlZwgn/GZvekpIUAgqi+ETDYsRNbdian4CLHVdFOlRcwus99eFChUm
TcxTy/CUqtEpUub6dFls2KRzMs0N6dzet55WgkJizTjnQoq1es0D2LrQ6xNHg2g2
+k52gDYQL9QCwzy0CXpErMU4mYovWtTCUjQKmyMo+HPrcPFbMS0Cpynl8yYhiE/k
n3bPH49pkd5Khomm07vNLtYdfhpg40gESPjP1D5z7SnbHR3ih0FyY8KYHOPLLtpY
UZ2InQPvGi+6IhlsWGrYRKiMvdHjUV7lBlKr4nYUtmO8q6TgbFJ2kfQymCZ7gpND
vObFoffOmzPQg+0RBepaZPSjueNPf8MWdx+RKn5FXYMgajeysD4Ums+O30efIrjv
xuZYw9ldrRPK/f0oE7AlFgdEwDwtYDHZhJ1RZ0r2taKh/P313o9L0GPCAq8k+Z2m
vi+busCrj+EOSMEOd5xKzbOtpl8WkYduCRyto5O1WpDKFTwZVJdAU81wV49OcHIy
A/7P0/pLOK6TsMd1Vfdg8UFGfEXx8NdoVA55H3SfHlBVZFmjfdRaCP7kb454EKnh
RWGEgZIR9rzJIJP4a5axHK9FwqJGNRN1o5oMZlte3ttU/HGs9AIApZb539zpj04q
8kiiTs+f0xcG5AcQPXKLVR6Ay47UXZAPemlpCUnvbamhrjBZx0Sz6kENwHviaGzs
3gY/Ye1N8X6bC9+q2qm3dgg1S0TlWXp/tYUiuxE8oHAh6MFbxs1ugOVfCrJ8epyX
zR1VI14DiqG+TuXvKCOLik5CrfxMkcmLPiNyzcOUc4PkQbjE0b9+0kHQf/nru0ua
XbS2YQmABh3OXbBSv9JCagDHasqrfHZQDxQB9zSDMfzLho5sTgEOHLMd29NFo7Oc
iFa3t6qJawMCqidfFRR26nKvcaQ9W3ZfIRm/yh4em3ezUMDJcy8GzvUBOCmuNoOP
DfkDLgO6T58gEOSPP9w8g+vjVgwsYKkzn1JUnSRVHr73unubiK8fvI62cnLzLsGE
Lf7QmxXnyuziQLpyG9PP7mnQQR4VjFYct4ftuMmyRNzPLpdRiA2udA3B4RodTGSM
HXMaRt0uWJI/6KhUqdeOAiy6xkg+2dHCyTk31z/77QJTpiN2AOv8QsbiEye/D+RF
YT4XAsmenS82n09Fxedeo6/iU/ZyEWG96mwvMhPmvYTKD1eazuvpJsCqHcSizqyU
4AfZ163JunK6533SsUqfxcwqKEoP3L1v56qzAJCrpv6ToA6WOAkLvwIMtLZdYf8p
63lx+rpKsmKIF2/id8IiJzi/NpWPjk+0nOX0JXA/uA8ttJ3q1mY0mxUW3wsq4/Rf
XEAZb8zUT/x7bOmj1+tdGNcokow/gcUorCTTFv20c6EZbe9umTHYgNH+5WodI1p1
TfgSoElMb1WudYsppr8YFKWkdhFxOYZ9oAgLQmxiXWF6EH7qfPiQgN9oIsSTMYbR
2YzZBNFcfxrUYrltJXAxikAXF1wNyuCM9NQWpZ2ZYC5MV3M8Nbwq9Uyk6Q8/ZfeK
vu2rOmiyKTq6CrUJ90I/7TQXvREv6QokzEkno5y2acwoP638OPLrTQAkVl7h3byp
ascaNVGdQiQoQJ/owSsbWolD8hGRRd0M35nGfOcz18KgXqCCyAmQB5iijDlPRRUY
8u+2P14S+zTmvyaF3x9hrA7awWqVeVn5OyomATNkcNUxLejDmsWUtanfVUJ/Bjju
W7cW+5gSnjt+jdSuqQfcgh9U3M1+WFJySUA0AgZ/CtE2W5kllRUdXzU/HHVaa473
0FIMk1PkdQBIMvb1ZJZCfVEZazcoG1tMgBgIFLxasmRPXe/kOPUD4jyj+PPxfM8f
8UOlayl4e/z2T77IdL1yeEZyFNc5B//K0Ah+3kPfN+2K5EHNHKF0bziW/EWN/+YE
xicESn6D2xzG4WPolrTIG1DMxHTt+zPG0JKIbc7bKm6B7PmiLyw9bYqBHAwVp+Td
DKc5gt47bTNxDsf8twODPQTH0SiuudmzI1rblIKbN0Iz9uSlgOqznVJ7iv/SHgZP
zoygAIvetQQEC1v4SRKjAvwGVTHlB79Ra9FUsPZF6/H+A37tSrUBqtROBXf4DKVN
OxrYj/1sIBCL+ROXlMSprKUqFNtzhvw6fX42gFXtuIJUgGSmWJedHx0hZy+pRNtz
ZlPK4TISiSHJnfM1KoHXI6lgbnQdLZKWUMVwZKuKZuFdzsmsDgw4/W7MZR2s8J0W
p6ZhEVZyaBrQmHV7KPfMzKTLfMTD3FvHv7wFlMZXp1WShUqnUneKdprSPYPEVtqJ
h0X2dGc6ZjKHInFjDjZ5byDpxJ5MG9TmsZcxGa44+B1xRJCcVwdvYgLyitJUhyc0
Y5/SLfyCdycrC008jkzGT4lcLThYvypNWJPoRP0Dkpq3w+YsxGaInt90Gskfr5Pj
q7Xh90Pk/lSuA+Ii15mqO4FIFDUtlg/kvf4UW6EoRdTOnJ2m1d8y7lp2ASIjxjE1
VqbDNxcGfO+zbspKX75JH5yxLMZKNX2vkFxMSXLvUhiXiGAyttVCSqYPh3u+URQU
1uzQbxWL0/hfbYQtQIkzkQ3/bOXhXhcbzyYifDQTJP5OzzlBOSK7g6gzkoIn8VDz
mBj1eblsM3KTHSKPoNOIJLopBtalEv6GzRHkoUsRdTDFgFhlYAhwpwz/iEAZiY80
cda6oh4u+WdOH6bQ2CLRvdDpfXGF/For6+Z7Q5oAjldgP3IZ34aeWGiR4rita9KU
aICVlXROjigQuKXixWIASbw9ECddCnIlmEPYT6/weQN389j2km6Z+chqu+ew5mZv
19dJFvpSBF0/tzKYjJzcQVASJD6naVybiYyHh2hOa2Jtr98GdvqaWIE8hcU1Kr7D
gI47L0f3Y9xLrym2HVxsdp9pt7OBQUhOXJ9PtMgKbOX0nsyKxA9ZcySsi4qZZ4Mj
6tHDyW5WK7Fj9RsNnZxCW5j+ke0AR6S68zoBapEYpTswh7v0x+BU2+Xox+Wvt8H/
SNNqxrx3tzK4aNT/yBTztOZJhVWco4AVT+MIRh2bmjU2KhaQc0xM7tDMyRDCqZB9
L/uF4kNCHKJdC24cEUGA5QCehA+Ur4tCg9IdSn5vB7ORDSdQrdhila4Zyphkgn/C
mOL0LZ8idX2Djj/h+L/MwMZx89occnfT+GZ9yxKGai5cM9UkZq66kgxMAlC0fjW5
ilk+fz0xFyx8HjM+zWR9Uw==
`protect END_PROTECTED
