`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npu79oC8nqQU6mghNE6JGXsizVRT0fSmzK+QsyE9GNjJBJYbeCWjA3Wq77+uR7nF
/nuWc4itpqRUnsK9rqW8RsKigdW2nMhOOEFCNRbSZecA6PwZ5JytxchU21KfyQAk
KmTYQ6uEfQWRvKmPPtYjXTK0QBy61NSyydwvSM6Mp5PWxAWONXMM5x1sFu4/8Z1b
2sVIoTJrbpYnSvkcEHhDTy6iHRgIYtw0oTJqSxIV7uVNZWmOxFg8j2saUX8mz66P
0h1wtwilWniNAukUXdnXDf3V4xswGMsjOJQaSDfmt9C1nS+GXG5McvYJ3MtllTEv
5ThgsBlA1OnAtX5V3Nxxm4Zw942gx+x4Xg2fDXvuR8NbrVzzz7WDM/vjE2IkACjk
7EGgSByE6qPgmTwD0XShg0a0kiCzGMuxxTwJRrrYLA9J4icvyLsQzAOV2W1qKNGH
pf6L2RUhmgYL3VB1UPtXet0/obS5+Q1tv3mEWKgJLpDpDlV5fS+Mqkw4KmBb2wVN
3PCas3zxWLm4bRMVvn5f21Fa2vR8p1WYwBla2fLxcGubnmNYnO9LLzELv0oqFy3+
LJD29eqZTuix5Li6R4LgGguutRyOlR7AtPr5/gifpeqmC8yji7jlhwAhWjbYg9KF
8X8T9RhBaun4dgM+7IbhrgX7EVy7e36JGFgw+Jl71E5MQxc/qjyuZ3LSqHHd+HCU
KkfZDPa3Y1YLzWUlYdD/wjwBReft1vJlU4H/kDKUQEnr3JhJhZS0qLZHTm97fyg8
xrnqZVbi9+dXyLlul803wpDRPYXCisy5mVyLM6IxbFiblOzMR6idkD+M24IGwmbk
MXZ3sOxSW2sH8UU8F7Sus0SMPOhqJjB97V6hVDzcH4NSonTtjECZlri93Ran9RkO
9qNrRJcp+Z/bKCUf0azwHtiNSCl7eJk6cFfc/PBnVp9AU4hcuVjreCWVrodzdGgL
HPM3ZpU8pMTFJzGTyXwtC3wVj3WhHfc2ySLe41mXophQhOtksR4wy6PYZAgf8MWW
JoBHY/tEUHBPsQrBsyawzFUIwTC0w/pw31+kGG/flu7ALD5w3VgB8k5iQ/PbRQSu
l+zMgIFU6bVGioSY0Zd1A1qTLwUxBMvliX+lAuDzvZL5n/CvK2ETPntq1OdqAkmZ
aizb0FL2loZnlMPoNimQx6ZN2whKT1XrTs2FX15WatulgI7GZF6Dk4Xw41XS9AO5
lAqkpYzNMbBeBfcef2nAzK7uoUzilHkPjTWVkSHU3P0wY/z+5LB40EcVez0R93sD
9pkb94I5xkbHACHxxJGaS/rTji8lVPaZbMl/B7zN3Du5ph9n2gNQO0Ed8hOwuCzu
boFtR3YNyHj7tuczLln3nQpGAW8P4ma4kxwHvnaCgSJ/gejzF7SIar1qrOwHkXYn
xaG1g+fJRyhTC3O8rWsb6zElaOpseGteEUZM/4RueerU4TKt1gyYFoIwvAZaVcwP
SRmbS1YLIZsffovdh0TPaG7e3GzGQnCBwY908lSmjsx+H09ZysiT/OgNz2wAugoI
UO+doarf3ipUBWcjxZr8PvIkkXpQ8qJvfK7Ty8xPGkW2th2UimfrPtEHdrf3maX0
k3aFX24KHaF812gcZMA7O/WwrCOvrlJuvMqW2JXCVYRgHBoKhjwv+jGr2tkYCWdH
52uCRHJXCDkyPecLmtUNfZEus9hdVo7KyYJjxh2vUWSfWv4eCNoqu6Ye92XpyPNc
RIvV3Mjywj8Df2qDnE0VSXN5YlX/K2+n2tCv/8lPRVF3U6QqfvgRftT6NrNQuW4Y
T4M12NkanrCV6ZICmLnDwLFlmU2tue/Qk5zU2FAzoDIyUVPfeZh65zj/dxH/jdcl
pj3oI7/hb6I0PHJGv+YT0TDep1ErvLdAQQffx2qHyiyRP+c1wOAAx9LKCkONAYC7
0dn5K0RSyqQiDNWOzTmVe4LFIlzRfvam07mQ/zsVtcmqEXVZ3MLN+Szg/9m82EeT
GYNzBTAQPRcDqr10I9hCbrl4cQKdo8WucxDZU9nzUV/SNrucoLIuNeSOQl0q3qSQ
Fz5OcRrYso/1Kc5mOCDDw1cC7tA6cdzeqv9sXlJTePNvfgRR1r/YmMInhIE9/szT
tT2tPWDrp+7PgijIdEcCQhyXRFBo9ITimyET7GG5hrRe191G+CFD8c7ze1783o6b
q0mWF8QctQ+NeWB30lJi/qvX4mFtPhJbgnzFGQzQp1mtGrtLfUKQsnMkgBdJGVZ6
1zUG34qCCKcqz6CyKF9nKKWaQCnMtC5/YhnqsExt1U7EeJvVvTsTzSbrj1Ppcmvn
bJyEItMDS1SPamKMo5cRAyiEp4k8Krlo62iC8h6clBo1T9vJkbbSKuBSoyQdbtef
YcWWt3551ypujvaReVzZXLYc0aSQit+6jnEMFgEIZBiYgY73XrD76AR7a+FmlVK4
7Ues+HvMMO4nX6ccigcqoOrVW1OrziJVbCT+sdz0adYUqMcXuze338ar1ssqQScH
53T+fOcCPC1mWBJZlv9No1YWFn8y+qvNk1BGPz0CxF+fY001YT7Dd6iYWSVgOeZ4
RC4cwULpwjQmx94VVJFxfOiqHViQFxFI5mXfvWq+HAY9zIErObl+IUSujvqvlnvV
G4tdB+oQcQgXA/ZxMlsXIeieHo5D1bF+u/xVNvw027uoXuQY1JUeKso6dE20IxpY
jYIOJ0HY/+/h3WFrJueQyGvPj1l7zxckdB1wqI9d90d6vDxLfPSlUuXeZSYsjUoU
Zh7/7HBq01wVgPaNK39D2Wdx9In/4SEjX5o/6llOA8c8HQOBOehech0Nkx+u0n8s
wx/4GL8UptSd4MOS9ClSad6/m+0FFIfk4fYHTc3A/76W51OBtJiEzjn/ILTfteN9
YiPLRKgMF4JX4sm5AFJbcjR37TGVvwewGhKsqWmniWwXLNxnv2eFT43jVj2d/wiE
BjuR8aoj4YV+DVMsPf0mz5ckpOACRmbHC+eI41LwJqvDM2exGzWqaxgv+AKsqHN4
SdirnvnKZoIOItzYfe5W0ZXme34ta5XBHe7iYtqyY3yzx1d5TBsQ4c2sNugsMIC1
igVXlh1sj7PXWoqKuG7QOXOoqKMrPntykPC27UW1pubXNn8SKzCbnibSv/VNgi9H
RIOvnTwbb979JoK8bGjHzASZNZBnXsKQRpdeEdYeot8Zh1mI/i59NwqlzZoduPoL
i+rOPHBMXf991+dNvJm7nUMNOpb0FFsMaEKUFxQqDyRAkgxscAlpzEeQA82XuIvg
9dGBJUUqT2lDwuZiFkiCvosJDxhzeGmPku/OJNZR+/plIuZznqnd0Spb9ljsyqoY
Pbv2k931dq+MnGQAIcS8TR3L8uZwMZ0cJt55G2wo+s8ATIYDvfmpDCIQONQt/i6a
tyMalYk+tPTBaO6kduDBOu23eMxzyYp7DkaXoxGYPpxXwKAuP3yWANvQaR9Ulard
ez3fO/1abSHc6doaP3pb/6BLytV4o+/btTNLr2XIAhrs7mF4I/q0XumBlZmaNq5G
Cj2ZIA+MxPv5WBI08YNP6mM2yVPpwv4Z1jaVRaFEJNoua7NxX/uSP6xMbjTQwohW
y8KEnH/UQ7mn5HpaM34r8kmK5e+BKQIG+bR/dufCyJ84L7f8mic7QLZsSoqAgcwj
20Q3XqfAU8iKyHKArwT+hHgu9i7XgCidTZHhUBkiM+I3xePvHdF6slBQNr9s9dWh
8Nd7rt4HWP5TdDX3S0ga/WIYHy8GlvqHEJ1rlz+UYuNuAjONEiJECErVx6e5myEP
/NVNORUL4of0wnDm43v8SBslrYEnWOgbbjq2jrd0VlLpG2aJmu+zvMrgPkVl8Ok7
dKXhKo1WUI49GxJ0yUCa+SC6/M2XYghjhuUVdRIq5a03E4oxIUuex9tdsvzS8lsT
wFfa6JuhFrySglzZy7Po/6kCaGweaQZC/xAgLzr34SqcPQAdspGadpXs5bWUG3DR
9SBBURHg1RPU0Fbd+MmlB+zPAuapa128HHwY9P949ligzu9kTewMnEL9v3DMrbHR
Eza/SdDnuqu41rfo4b/PEtX62O+drtfRlrMyyJASzc0hDaXU85WknvRK6JsxArF0
uJzRG/NwobsNNG1xtddnk1Mc2h7z/9lp4aiajUrhwvTAaP0oRSkWIjOUW06FpJCb
D1zk295fAApu3rTr7Hn9v8szBYDWmouZogDdmFZpzgY8J2VkIdOk0fGI6pUS6x9Y
udeMxKsR66gjwk02ORPAB2peHrPR+4n8FwuisBcN7Ieyx5/OiCSh4lSm0Yxqb2Vu
K9w7FMX7mc4TA7KY/nan6lZh4DCISg+UAwauNBck6bcM3lgBtzAS4gnVGlL9WsaP
c2npAxPpAXq85DT4XWmSXTS7a7woCzzFHmi8T5LRHwp2u345Td0ZWZSZSF9t0JSZ
off7Ybc8zCJw+B1YVirYUnsY1D6dte5bMpTqHXsx8eE70cCE0dHZ3RBkpryYbZOa
AC9wLHNxIunMdInfJn4VKL3zbDh8ruVOiiwLPeVSlyKCHX5XNtQHw/1MqNOXUkZT
mI+tzkQcLkfuZdl8mifD3YkAdfSm1CxD/J/xLHYXN3De7zsHQPIcKWQ+vZcHwpPy
vgHLoReMMNYmixnhsnFusQ==
`protect END_PROTECTED
