`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81amCTtl3sdGlHmzBg5AH1e29qaNBmRTChZiP0yWzlGcKK6tbpkiOrlLOJ+Pjogy
kpgabFVLLwJx+sX03R9vx1+mDCH4M1SVlOy5cnEoO58eGlP8YqmCFCW0JJikp0xm
RoGjzW+GV4VSh6BZWwccE0kvVTHdLH9ODiRwUwo8kkX9xIZDKv/eKDjQBeVbRC4/
HxnFx34x9DsYo1wlFZ0jNE9EwOPPhFLc0sSkxEHd/ihRFKoDN2SrT75JVVb/DdQD
RSD3t3qkXZH3vAWL92bF2u3Z7WGk5HlKDymtjwEYkVSaIzdqB2zeYyeKh8PN++O5
qHDcDuYXKV51fsM2TtO4wIiDlUB0YCji5MzrDFickqGmt/dpUuO8xN9lgbBobkoO
3ZwmMg0m4uMMX/V4XgbEk9j2D2goiXIN5LQOI1f21DeiXw9KHzqr59MuEkA6Y7F7
QA5t9MUuG6kVmOhmdz3Cp6Jera98szQTfiUG0b16tQA=
`protect END_PROTECTED
