`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXbnDsEbIYbJfvLrFbvuutOhup2Vnzj6aS/wFMfqWnLcyglZEBy0EnH7FduVZrpX
Kh6knySHxPN/DKgZWXvXEo9V2nyVatqtKuVN4qJ/wORtAVVxLMGgCYa/xr85fFxH
6/Qlq/6B26NRMkhSXujeCVd8X0XCVlAB6euRBOF6YaCyWv2ARrde9+4bumT3T2eB
l9DT9K7bLOTY/r8SU1TWUkd52mtW6WPJ/OgxVPDOkdEMwE1etoxlAz84pQWPVu6X
XnDglqI86vF/DgnDwW61lojBe7mDGwu5ZCRwDUSo9N0yMZ8nOAPFdw0nwNv9Hfei
b+CHNzmEcpfaQviJ2X0mOIQXRiZvFU/WJVCoZfc+Ar0GgneqX/zoHlr1gvoxp8CU
1cHJ0tO58qJo4T7inGO76fbGcvPVxK6gElIPEt8ZNXkX4lSLy3Whr/OA2nWy/b4n
h/lpwSqPURAm3Oft2+j0zHB0AgkmfnlMEhFyrgQSAZhw6fvhAkZjFETA8hclPWcb
OaBERF5tvMkEqj2CAmp4o5m8Anxi0FBwe5d/6jq1AlXhV1op8YL7Eu7/ZW+g5/MP
LxQaitEPrF1XCA01v5NZmv31khuoiIgT/W6AUh33B9O7yz10eZFrdaatWX+naHK4
67/QXjPzSWtz7v7Z4TygSUe/agVJf13sBmjsXIOmOmcbomAHTM7bOHhWYTzqZ5XG
dsVbfr9jUT5wqaFRqo+kPNowfHGIdYEKNTWwyW6NNfjqpxQfRFxqrUb/azvImORJ
KOZnsYi/1IwbtcwWhCDFReLJwFvOlYMUqsm+/Pty4Qo6D2hQLZ6sJ+S1fuLLqkQC
FpAzzwCFFbo6xizY1C9wKctPXnn647gOBW93x1DCDLvhcFQlczy+m1ZMbRWq+I3Y
JWHSu+e9dCPiR1vI6ic8TH3QoI6RjlkBaCGIYp1bG3dpicz+PQP1Eln43QYyBdD7
igUM/eXDdQH+t8FzIitO59qBmBvJnM38+YaNAJuEtK4SU3Y2/iytByX0VQg1PRgo
6pTBByZtoc+rJZZb1XzcDyMDawUSn55ouptkj1APrrha+/g+3UBadDubJZrgkjZ5
nCrJIzVDnBMLBYuZR2qRIeFbM06+Pl7w3WruuVEfw4U+Kyvlxt4q98p6QGJyY6kz
lJhVb8h253hjlFpUx10WT5kVwnsfUUHukDk7eb13mfHNVgPqlqcuJ/XltCwabGzb
`protect END_PROTECTED
