`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uD1220/Zo5eae+LTsLkgT+NpBLGDC/gFk61n6D9QyZfkXx44dvM3FZ5T0vtsBafO
CAnNfvdmpeId7+Tpoae98LlHs/us/BU3GB/YCs8Eq+UtfTdA3CLsLTndl98u4yA0
UWNC25vgG5PrLUFXqLQjIsPFFdtN7SBCfszg7qAujVYPjOSrT42gHMQA0sL7ZY1R
3S4NiGnd7rdtNJSIyImJzb5ssIQV97GuRMpHDntAgKLCxOgNNA1x+UdZcHZuv/79
10xJc/GdpPxP5ZlkAh3qyt0OcEoIcSm/Pl1OKjj5qdzcgOe1n16Rc5RoO9IGxNh/
NHNxG3WFLoxhhXDMK7+ic6xGbaPafScO4oxSaDcvrO+8kSQBoAytZh7Qj3DxckPw
H0d0DxwNvKjrUUU8tvV81Boxs9nhyg7Hmvtyai6qq2ACQPVJ2xoN2sjvXVnH6YsE
kECVMl3/09PIQAOkPuulIG+oCK8wsAEIE1+FOXanIa1Sr2YRpZ6qG+jKKzWYY3NE
wg72NRSKAbVvejwkb7E5lVH4+e7ddnxCP3AgSL5wTVoZ3S8HOYKKvjokUUJvd7Zm
AvlDNzjGVQyN0vpjmpfi27CJ/+gA1Hi1ZqixSlqW3dYPuAJp+s/31JDjwnCzD3Xx
/9WXCaHci+5BoghaWXlu8c45hjU4cJE34ZD+doUaH5gGjMGjGV7n2VAiV+uU63/I
d3S6iSKZ2FRbM7mAXxp0FUpyls8VcIX8IqJZD9PjMvNd4uU4rUYiEJhSap0wWJPd
oQLVknKz/dr+HvLjbNn3L7k9MVIco0oIU3F0zQMBetk1v+21x6Sb+70gt259pmTN
nKwYRK9fNmCT2Io97cI8FAPWtrRenxrQ3X2cML7JBpqqTbRRe2Z3QPd25IW0KSMx
85RFx5xaSrAzCfuFzPADgg45qW0Jk+0IMcfE1VdcNJ04cjJ5IaBMlXT4oMRrbfW6
bMk1szOsfuvYJLPU3Mr/cDj+h/NG6xzDvsAUBOG1Gy6r4YGrgg8+1Fv4uItWuYNQ
ZApSam6rU+vxEY+uSUBrEJTiS+LY8QZuJ1a5vjJSNat94JcLVfU1QEtDBwUUJ0ew
r0PafbV8gs5uQM4qDYpkV6y9R+5sZZJYNeBckIUxmtZeIRydDRnjeHAoz2WoduKk
9BIyfXY1r+FHXVz7Ik6Lw3+DBLNrMd4RQaga6HObiv3cd0VeSgCezhimhtgLMHXA
Z/zZKH7lCRDn2rTLRN2fRyPeq6VLLojsQXn8I1tkfQLZmJ3jbnX7vxLqlgyynF9E
XSRiyJUPtISaKO8aBad1kxkmAQUBESmBF9xyn6SxK0DwuTh+uMkolkj+/JhIgSeZ
ZZoh/2NNfqgJ3/fXbxq+ydXRNT4qp3vD+0lhgTzQd3rKtPJULiKdJEBBq6CCUxP9
km9fzcldsSosEfGRDH7yQQ0yqLwLrR/qeckGpXHjD3ApQlZdMWZdU72bkx4BViVk
wZwjWVwXAwNYuRIcc5jVnAiztEYSM9Scwpl0UlNXKqCpr8JiXYvz5E1pnPEdRsVD
0ZboH8CsIks3Vm8c8CU51qmSJb1f5I8qCmWDA52jexagHYQd9YAca9JNj8YFQXcl
oTvWbqBiOnMVxkSEvpPR7wnVA1XVbNh5BhBS/G1GEHalttA24c34rEpTNH+PFXsl
NxUtx/UGGLtMb4bze54IxkEibzNH8noCLVKWipqYCJzO8hNT6A43JBUvhvTNR0Bc
E+F3nZDJ0sCaZCt1LjoQTKhbq6HaIkD19d2MS2v53SyYWFI3ZmB0ZzJXHK2x2np1
E6NCOVEHfZBfqbasPeiu4ZN9/WPDStEeFoqg7lMlels07SlLF/E+cFnjEMHoVT51
ItRGbwduM2vxayeFDg70atcTq+vK2vRCnN6QhmU4aVJFlbXhLv3eMSeDEhnp0o9Y
eE74eS2DJ0fXGNlUfjS6fsI0h+2CrLft8eicMwOJSgsNkM/W9ybO+RuiaRJR/Uxd
NkfTk5YtgYFydRF7fKYHHfuLGXIEbjZa77J80XQHoFGFey80kwRYCxat+KzKXP8H
me1dvI24wx0DdQilvWxnf7XNTvcINHzzlgtfKbiKcrsGIcTZC6JlpB0AH0TQtNo8
t1SdXfN24FMa4J0vefzdT1P/+ZWZ+M+wlXt7sFim6WTXPbicAle60OpQslgKocgT
zraNa0IDbFEBeVwZISlH8KnietboXInRSo2UqHVYnkMHPHw06dmC6ZjvlzUPOXDF
ulRRciQcaHiPEMX2XpPMmQx7igZ/IkL92LCX+ESZUBoilfD9AuwY3gOaaozO+Oq5
6VI1Bex3cJnrxGZl4tqO/mnRdRLnBgIQHDxdTz4bQSB2WYRgdlqq8zsemoDcp8ut
B9sHQmE7MmixLa+DklTFWs1IBaK0ye29368iK9hz2RhMYTS1YwVIIf+VnHCqfxfg
Q+l5HmFb/fu4IB+sxDzZb899wHJ5V33JWw+80b1dT96MD9J/2Ww2ro8/NJHIppqC
iLq5wpzrxM42uhspdhQk/r4njOtoA+T1USnxd/wIhhs4LyIvK8XMtpberwqlUXnF
125xpWwywcBX8AW9g5i4B90muxQYhdE9uCiBPt0TTuPWhboJe3km9qbUQl9nfWjv
jDaX6y3A8aW+1KKPsJ8Epmk4N5SBWgFSCzv3E6y3uRlxCoKlFGVC9p7dHB05/lcu
OSPgqvf/0ASbx2btdxD2zg0ggxJ/mUk1Lhb33DrgcAjdb9hC4Uvla7J+n+5FN8wT
bjGncQPzFeR8KfkAP2atYMs78Cn5PP7A2XTihZ3udcgkRELl2tJuhieGDHXf9aAg
twGYHn9xYuoTBlD3EzDmixS44vzuf27NtxQoKd9MBAnZFtoyludALeN4tlyB0OCA
HpZ9CACPpW3IzxunEUUvbT+6hMT4AGF4RTWUe7ZKJL7uPp1tiYCOyYwHd9dS6/pK
MSwToHRQNqcjwc+QXJnaPOVzyPKs96IQ4cO30FcvJmk57bD4FLhdmhJ2q09/P8dg
alK5dsCSRB84rF8Ew1WTHwTbZjtHiaOx8AoXx7xXcfECbZPRj07dR4lx+805VoQb
GuOriEdtc0C8H1hQMPAK0YllQfHvfsoFJ12gxO3lFWYJuui4Mr1GSIukau+LBjKK
X6p31SNTB9sZM2MnDu6SGNbgsJJ6I0SSmrpWjU23JRxKEqPUf1Ac/VhYcG9RijC9
85fASB4T+hCEv1DAzTY81VyN+g8kcnpaNZosqz3JjC0DUTYOuvjjaL1C4UNrf5sj
dkZsKzT860IQMsdzf1DtkJ0Cex1LSpPrHzNXUOL7eUgTsTJtU3sASO9uI6jVySmy
ogG9cGKbfmcCZrnrPSlbt0scfKwH0c/X/tYbMCKNII8NI/aPzIu3SJ926Mt0kUaK
9dsVZhWhkA0PCCu6C6J8PH5wmFKrrHajzkjoUPgaXWgMNT29OOksQkBAoSRa79w+
eKYusC6i+vr0cISvIXgSn4ierA56EGSn7snPMj0uXyyIwmVWHUpYK0fXlIdWL2Vy
w6jaJmm/oc7qHC2Zox5ipqncLzntfe285jZgD5XBStOxbmUOZ/4s2K0k/sKGxg/Q
bSmalH6q4XK3W3ucq/czXrV/lP+6IE4kTn+xidYjuy6j/cxSVaqsUq03RF8FWzpl
iI+TPeDxkz5ybXo32ev4ZrW2odyKVzwmhMpDF72sQPjMm0BStdm3DQzHAsOgAtiM
F2jaKeHGtQM05wNTofAD0XTqUsPaPZd1JMz4AGeRXVw5gte/LC+caA2EXJ0aegRG
j4JB8TcSbOq+hVJGbD07msJLB02rNTZbne0OG/efmZgob3ZbFWuefcJp8j6dFLMO
SYUqhffDLPySIgdDrTJm6UVN18rNhDCThUCLq6Td5itJTuGurMDhwVQMgsD9n2gf
BPwb0g+PFAK66n90o4MfgBPfwuE7dokr2I6Twq0z3VRnHQURZFNjqjfIJeWf0kTB
+SCpMQHMac7RhmHQ0Zp7zdYvG/zbMp5J6AMpzT16bwUAT3Wiy95cxyXBKoYEE6dx
fMkRpeNn8roY3h0/nIRjP0IVxOcGBZO2TubjEt00fVQ=
`protect END_PROTECTED
