`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuzMOvaLjtxfaljqQqit9c1ReXTH36Xk18Wv62n9arpGKtKyjg8MUT42TM+kXuPM
t1/zsyDw2WXB1eH6k5F/m8m7/z0VgOP/5l+pFeQwjzqXpOMyqi0Vei+iXHq5s3oH
kTnM6tv7WFgd7IbjCQzL/7d5Tam89DaYtv+t2sDaLuq1JHnpWx+6JLHhgpQcz1it
sCoUw3ukXcp7Fvcgch08BVNZJTfSyicCAc0w6gPGgPu711LTeIUr5VqDn3i1oEYk
05I7z0iNYRaV91DZvyyZgwdC4HwF/rHOtYI1vWu8zGphYFTA4Xlq9knii6wPcU0v
ONLI+0r+eMaoSqhi6iOtFjLjUXHZFn/Zd1k+1y5vC8uTJo00tmPzc1GbIcDqHnUX
cjL/+ror7vc9ZAp85cWWG2zi0ngOB24VU6icaIpWx8g1+sZYp2q9ejaau0h1yX7z
zEstRCsdjYiSjzZ93A87uIm3y4kwMKU/g4wBuLpU6lo/KBr5PCHj3MX1SpJZKwIT
BZrpObSkJQQ0VE/WnhxzeUtnNP0C6mg9DwyIbrLlLlwu4IKnPj2Uxk8o7KiatJY1
UJ5Qe3G/OLj0rS8EhV1bHMi7GVzuutBwW+kwvUkfzVOQUdPPAy1geAKVc07N1Jab
BFjjaL8u3Qw/+O4YonqcjbWPRV6eUtudnBKJquArPo/WclLGX16Ekyj+KTrahzpr
EKis4K6tJMKwropYp8m6ZXDaW1KaffvSAMNo/Wt8cMtaPFnvakQsI69Vu3h2EHHI
azh2wxGWB5FfraX3/zAgxAytDCzs6c+BsgLNyhSfhDRAdNlrz6JZ3oxJL/RuENNo
vF6Piy6fZi0VRxPoH3vD6vojsntF1887/DGqJmpf1El3zC3jQjYDnLLEWEZDUEAm
d3/FSX4mJ8eFFmLQfBkwgpRC9mZZXdpG6TT3NmCC7wJpLPEZzo7nJEhJO/6mHtBH
W5Sb4AKvGRhdTzwIp+2v7RNxDyKUOoXxHVf2k2CxgCbPHTkjmiyD285+xPGOK1ow
lpKzhQGBFpDIul1x6AZn7iH73z4fuaZrDbnwrNGqfTaANjE4cHuhZS5rRz8fMAFO
vbonuwACo6Ee94zCKvV8FYzZYE59v07L0agni0yPIhVdriV1W03M+nddp/v/yj14
449tnHxIfoG0mapSF6tIaEwUWT1t8hannCN9Kce+8uMALodtn5a8Ld7V+GsEYPeP
NMk1rsc+cmzbsQlCbS9PCEq3TmbUDre+n4JK0HGFu9A=
`protect END_PROTECTED
