`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IF4mDtqErdsns9lcqqUYAE2cPNvxplzVge8DKEPlhnPwvs3n6mJGo6nqNPXgszjH
X1NHw2uCSzy8XXoP2nmI1FGXlEgrda0fbPKzIXd2v2NacVZZn8JlFH5GDcD5Atz8
mewhr2DeXfCwvGBwDz3hdQ7cq+i/ih/hgl63bJiyk8MrY/w5AhLsADrMixeZAFgl
ejeGErq1EgrOt14lQ0ZE8/9AnZNoFueyxvoOgbmJlquSvpn2+BliEbunhJVwroCM
5rJXU+sgLYxqZsrfcCq7EgTg4IQBo/G8GrDRoTaLwFQkkRgcd/A7bijngkTPJbnp
BKf1qIh5eRs4jD1Cq+ziVU5n22U0AtYw+VKeo4bk6fYBxs4aZSg+V21euIjj1gNB
FDxWYQ2Qm4YyhFY4jvt2qc3ZatomF6vDvpl1G5VBEk3a3yIaopYJ9vndz6xvyx3b
u2ST9wCFuiblAcHYSl/7P/tLBUeU71m++33F9108zlDeAEU3Bs0RuHlCe/NSOyAg
+JOCQfLK8t6fBB6aB8PGESoH/KIjExnlInXRqPR0GrQ+IAiTMoluyYBVqhD/JHoi
S8/7auOOXXSq83hyVWK65EzcxuGVbFLs7R+PF+ysu+Dsf6RvMktL58urOv0xGwPl
gCZmxyo6jG25qbllkCqkPkNryVzD0L8yWLPsk007RB6j1yIiISvtcVGaYqyPq5+9
vZpctkRYhfYoIrWTXcjS0+fqX+HEo+EFD0snCjqsaWSVmNobaXQd73S4su0a42ab
WfWTcJP9/aS2lQJeToVVBps6erOm5MBMASHGeJxL9QaK2I3jj9gXWPl40dZkFSBp
PuDfEaOJH797O+cQyhO48iFeetVcvyn9Bv8sCMDCiykC+XdUk9JKVvkLe3uWNRbt
HlvPHXP36REA5ve+iIMcy7312GwcFq7E2zT6hPJOJM0vw01yZ4L1F+nDpianK+bJ
gM7aNvJgE8T1Rj19JFiUum6J9auCKAKjHqJgezYIdtySFrAMX6Ahr2ulzv4aQUXh
O1lJvgdIbzwkwM2eJMgnNtxba2sMpqiG3q+xbyDqZLBwMkVraPD04f8coihKOeOV
xP0tSftTEyzBEzTSd6Rjq9xnHZuSOcIT+nJzgewQveChJRuhoo3JJEzzYQy5C20V
lcPxI/huw3jehOIgYDoUvOULCVP6a0j7kFJwQ6GVKzuiiT0jGMIA8cdJEFvxFqwm
vmkptfkkD2MIc3FsNdmeVaaUL/xOpHKpNGY7uSZrlwXhPUVVZ6wNvYGCZJ4Pemw3
3OAcIrT2ZXqSJz38ENxuPYdQvCvt6hhd8In9ygwYKAyJY7jIJiM7A+4TxxZ0UMjB
FoBo+siwnmH0OjOagd/ZGm9qEaATvJFZXmFmAxwNbcq3Sonhq4JZJZnn6uywNtzV
5s86tgHdwXs+8SbcXPBH4sXo/VIby0nXtXYnimhNBrvgU19fNqztj6qsaehtbe+i
wBeJPaG9rod3gSXbKA69iZY6j0RX7Kgk2zArpd3hUvX9ZOizG9KP0PM9pAx4Eue+
LXfpx0T/7VBUKzrHLb8K0bd8u+xNYbpYIwQBHtZSX0AKJzCDuDVzqmXfpDR5nEif
qXgr2MI/qpQcBpukDMeTe/5bIpr5D0IM8iI8ECiQKPxEvVGlmrPlIRMcLHAEZMwT
ef5mKb8pkvBULAGHYjLsaxbCc8YQ7kUh3nSH5ed2byqXncu6mOkVRtElWW0aKVWX
wCCBNVhVgorqHWinNJZcI5ODmHF28MI4Yt7DVC1Q1Jf1tA8b8gs8nrRuyz61RFOp
qxWA/6R+4yv9JSSZ+FdxPZiB2WQO/WNG5Ws1yohLjs08CudzL0B8iUA9WlL/jf07
VG6YjJwUW8vfAY+/j0CfMMfw6CrU+i9J6Tu05YUeUH1WOu/9oYFLLvUKOPv1+zxo
NOM/LpBAuo86jenb5q6BUx3xFlu02YRi0ouu1lToCKaLVf2K2Rfb1WkLGlprMYEC
iSls0lIu6UDiyQQ8/J+mWcB3Zt4Ze22xajoL0CaRbQVtNRfwYDOQ0JnyDVEcHxNX
x8TK5u9AXQIGrIvDnM+wjUSjnvtvpper0uBgX8Z87bfDWrMpXGhMUa2lZKjcKezL
7F5ffoKQmdU6FKN6jkOUJud5drFWrnkLWu8mrhzG1uX2nl1961DxqBBj/6UGiNXl
VTyxMpqLVOO+TT7ejhOIP4lV3tvFsRCY/y2pZEsA9fcxa9X2i5ggj5yWKFcGgwun
wUyrZjNQRZzlUGTYcfbBgbfw2SMdi6rFWPcEkyvTdBfqpdO+rWF2IHZw42S6/Mhd
TOxBJF3PvG0O7mNwqdRsl1DlM/npl528dxpahDPc/kyhOS+2dztWyk9A0w6c/2fB
ivutRkPuGTG7ScLdH/9+HL6ftokRyphm3sE+h6T+n8cbnUdjx+Z+EoEIGYQcrEh7
YysOXlS8gREslqkQSzaQmroDc1Q6rE2fHQguX/YYcGHAL94p0a8ymCSVMMc8dEC4
SurtSFwjbNUmw6Guj5H4VNzZsN8vqFH4h2npV40PeVWki0nUlK7+v4v8FVnvLDM2
XgXWd/XMFCPIGMAXHbkLBw==
`protect END_PROTECTED
