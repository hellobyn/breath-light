`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hg4fTIFN9V2Mzcbn5pHwlTL6bsyOIRYkiBgGtYRBlHIb9YUY8A0chB+K5+9Xlsau
+SWQBnTgI4g3s9fEQnpztl15/qXyIHfx5iBBc8L5vvzC/Vlp+q5B2AofecBBPOHD
k6r0FjwFl5RdYc/Mgc0pl5wp/3Ia+y6undDJF5CBolX6L5DScXCP2VXHNLK/USr0
V7Fx7zX0HJH4budz9xLDd8GsF7m5CHdKoLrP/ey65bdZaQMqD0/11pOc6mc/Cxmb
a0eV4g712ltCGAeRDLgXt/3Q1qBhdC+QUBgqKQyivmnxDEqkkIkk584Hlmdoars1
5WlFIN35pkdtLbj2JvB6Q65MNzN3rFoetrEiFBecRtufgqUjtjaXXOn+QjIO2Cpb
xhcQ2MsfNKpffwuWrCSywMoC1g/f+6Yk6bZF4KrM6bUNSsabT/AfZKIw6zdIpuK1
AlmAZON+LJEa6OGB2ea6ADHBdGHrds3/EXON4VeE0751SwC4YGrKFhnQ/B8DZqE9
6ftM5mIeCgpa34o4ROm+vfe25F/YP0DBftPG58sONMOjCDqyKmLzwzzPGbEp6hTu
3UL20TGYhfSe7hs99OuvXwM+M5UrBtXJ24aiLvnEydJyDVywXvf+DeTsx4x/OjlM
LTvjzJzyUlQVojBYcmbo7uN0gTCVUzumaMcsN7fRmXtr81E6waGUuT6eVl0FjlhD
CIuYD/7zjCzL2tNscKj1+4gteLDxGgFUi7JRoKaBS0Wf2nORpIDKNcG5DKe41kof
aumhRqxIbNJIxUjj1qVePAuZoBGjVpczEsZkXFn1BSlKfltAOFaqT/jlw4Ov66o+
ZjE0p9D/ADUOWCd/+i7Iij3up6jVNqMXda8hITJ8EhemzXacOeOj7gRZqzFsUbRk
QU72kM+uWuIsWl1ewzA7eGXvnP8BfEpyd2nHL9Ft+d6G18fxUYVmlS5WZODE79rx
Pb5SqbE7uhpxplBLkqJFIm5mqf2bO68vzY1fPKdCCrDz/uJvP3ywwhJO7oC4CHNC
ijuTBF1kdv4xarol5Bsk6eSNeQoi+jXJJc9jrgHYDOF0lh+jKolWHq+HKBtgM9Nd
GO/aKBE9K0tyMemvZ5QLdfj2o3TNuwHguY3HGXboa0rKP/y9gPq1TWFCnkIVEuFs
bQdGEI9EsZy6C/NZ+FwG13VMs/WDacELm7ShsVGlu+EZgjX2MuNuDrKFh+Mk7lG7
a0r4j5fQ7xtAe9lfwFuNsULCAocTfDCq6IVdmY8zwHJBE2lmLhKo1jZZQxZZFVh5
JGSLHsH0ZhS6yblM1lEp7Sm0+78JTa6ENaBZo64yBUJRPXiVo2df4tyR2wOUG/UL
oGfLYpoDgPAfHjKD/eyTEucsZeqr4yxtCLY1Uk1Eicv/C9QUenawbxrdNFccIGp1
nUBb67KTHAqTomcFZBv28I6Q2/yJEDSgdql8tyK7XAzmG0mWgEimTZTh6P68Wm8t
mA52p0Fjx8IZxrGPu40QK3X11jZ+B8NhoH08MFV6Yc6MtjwQ12WRbInlswzRBMuK
hJnK6XNk8rZwNHMb9vBK6gyvEBzPsQkYg9UKJIpaiYVSjw8cy9M2xN9M1FZI7Cwc
eQi4MHtJ8I0A1/98HhVHzUTbfTwpBdIn99Ul19HTZTbBHtk9JvijZm/aK5E5pTed
hQrUUKEx2PmPaNMrfspSjEorHN7K3eQtvBqM9zgA/0WBeCUQt8K66J36+sWzH8t1
gyXioOMHJYMUeSmWfCbyjNC5OSnU0e3kYQFF13fOcSDyv54ZkreO0ryyfdY2FX5t
8V0ObVGIQ0HsGLKG98BgUxgxpNgeBDwvi78UAP7wlKM/004a3/fPqAJtXL0AGLkt
XAY/XF3FCgXzyg92p9uwJvIvTiASaTRdJWljRYpP5MhhCHIQIhJqffbyDc7mBWZz
mGSLy4V3kM/TNF7L8VQUi+XvL42ps8Dl2a58UwafnNx2iDKW32RDbmWyOLZnwBey
sBolC3aB/nben5Xftqim1GXYt8z/mWGoM2XsFuhphNvcyFQChMtV6vw7TeGQkhjA
l3TrztPkTQFWzFVMlqdT3Nt0kNyTf6M1u6Hj3llFuOiu7eGHEoiaqbkWKNdMh5kv
`protect END_PROTECTED
