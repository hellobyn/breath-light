`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7LEeDK6O33TzW6FNQVVyFgHgxGjT39HByDM4YLXUmAZXhgytB7qjkY6Chl5Yy1T
3h6wk3S2vUM91L4HuSydnoD917u/Wlwj3u5U5l0uq44iB+OigZT3djEtxEybFL9Y
xdS9bZyodiLPd2uovZUmK20UveFNJtEV7LDWARYje/osHPgvq7Ue4QdQ9HIfMoqQ
rq4l81MxNA8sa+3/bUjZa/RYPDRZKlegeUrjSq0+MLqerDqL3PSjPc7INS/aCtbF
+dlbxmiy9K7DzsnLcNxy1RyDLMUY37H9IA8B9mw/24h0EGER2kx9JFikQ72sMD3/
jO25d/8S+bfXqP0apTD9xXy+ThHxWum7l/jbXo3d42NLTZ5bNtMfDiuBMejNIN8R
kunNE9lrbqv/XXl8ssFMBjudM7izN1gpO5xVsRabai7H9PPrbSMbBuYMOsSIoeYi
d6AlDgplAthiUQuzNNtFenNdY873mVdBZ7IqlH/TanFl3bcmVbWcRohGA86T8afI
+8YjRCVS4yHHCR03i2SAM7DOKsgJpsyxCb0XdAgQh7xLsK6QVVGKIeTQYGiKF0bb
wIh6YL9qKDGSZO0xweNQwOQjqR+DLh4FXgsdNIhFslApIexmxccCHTKTIOmKZVzl
QMZBnkmH37hAuTjiuJBsInzFPVJkfpUmzBbTiA7sEudqtRPmKhRiOJB+UDPixkGC
gDGGlokUn5LdB7OJ+twSATtKrLHkz/2VejXgR7/xI6J/IR8YHuz9Q2o9D5nAOQyl
7Bcf0JzgQ5PPgkdGy8sTeRkVxAbomf/cjQuKGRwLOSYCCmCS1d0a36qpeVLnkWwf
rvvio7hvKg74P0S2bMh6ImRL+KrhL/MHdCrr3Tg2VIg53JZVsSPcQ6I+xVn5F9DG
JoZtXK9JsSiSjm7MR6qc4msjXEWXQORLuamh5806rYFsuPxBe6Eg/KLrkVUZixFG
ECOko80Ykyw9A9aVvMFkn+uXPGp7O03rjB2AY1mO5UcgQ+LCtqGp2QcO2wDXu7gC
z8wCD/JkGfq5Q3dap45X8mybMQhhEUWOisEL7KbIRMaU+ZHmqYTQHULL+gX7hXty
JGqLZruRC+t73tA8PUilBXQWNg5si2dxLBBJX6oSBi2mvZImFzNAc6MhfpwNj0TG
TW5IKBkfQft0BM3gXEm6EIOVpTFIxbMR5qV+Wg83ZaBpIXDiMwH8ORzp1BvqhtoT
0OrhLnbK/QBFMNxh2kuzmLhR5WPHe4lLnd+v7gkEWEdxZaL821BayPI0DgsxWF4s
v1AosiVS0MOkTkwF0C2oxfyNPt8ckfjlMg8LZFtRGjy0ZRQRDbDsahdLQB14MvSz
slIWkIv0ACLMrLpZPxb3FU14OTXxd+tvQtcChJkdDu6LUNsSp9JwMA1JuqI1LYnd
0ZLkz8QEXNt3jpE9PMUJov9XUrtCx9Tu6yQO5XGWhVLoXImKidXYylqPX85OoQ70
hhOoz5vlhRSDg/8bDPUVA/+g57EEg7tdITMz7F+kqwggGdV33v/CzqUS0DoIpnUL
eZBwFOzDpjihSrf0MKHk94zc74gUy0dnC8B/IEPMSXbPSltcOINtfb4KX2guXSXT
rbEnQN8XLo/K5n68tPKr2DqG7DrFMEDHTBZUoEDuo35UNogRIHSZ+LXJ43lnSOhq
ft8OF76R8On66/Gg/umMn23onS3kE1M40zQMkHkB8K3N5Wp9jmQe8lEqiEr3z/hF
zacFGPgLSb+IswH3aJuRYXQNy0jpSMU2rKeH4EDjeoFbyZYZqDPgL+nwbSxkTdsX
cdsjQBnOexUJqkDklZzqDdiMF7itludMBT2TCUAbCqaL5IDcMHVdgcqoEJh42hf+
06czdBSD+H5HthAZ7yuBep9BLQfbUYu8qzx9LOS+CUWAxjpmwT9diNENxnz2S3BC
vDjFcc2p/qMcKweG64scRTdUC2vG8tJfDpNYO/zHqv9dWDJ4yCQ8oBudrX/PM6FF
OmN9AhgYDOlKmqGzdtyjv/wjdtXYBucxwIa+iuanTR8HU2Hann0USq/2KKkGDizE
udyaYSCTCsWEZJV+J2Y9zIhvj4ZyMswX4+By+atslcR7jXvajJQktN3NaW/KhCXq
c5/tdRa/ouWe8ezmr4dIArQX4sa23m7CFSLLA19IRRy7iom3XjEscEmdcpn2kAyV
AbWmNPigAJHaOEoQldy8maa8rURaij+YS1ylY1FrzEGPZnDW/PndDn7/YnuzjM8j
zGMUHs30kyBAoMCvdfs+r0qD4A4eAVJtW1pmlvvyhEpOsRFeLXLOiZrdJk2opA9U
fQEghWWSG4ln+yH9xyPbsRsUNaa7FW11k/45coM0m7yP2sXhkn9Y2At5G1oQKJ0n
SPeZa+fn7AV3/1eAC4nsWkxStSjNUMydIDniq1yutlNycg73u3uqWFcTZAEexV8Z
vfLiJCkUklSpY/SiMab/b957kqQa9H2nUcGwNMZETDT6YBdODBrLQZRap9j6RVC3
nyUKBrzY0Mj+fcRCa5grYKGexgiA8vweVI+/39SL8v8MYS9HzlS8O5QUBCafaUDH
Ejq7hTQcyibaGQpd5WDK5nBSfSN1I9inJGLL9BXaoLMuClsjg8cIRfgTFEsqhzF4
J3d3MqCenZ2wJL6oKEO+42n6kE7mXLma6kLD2bOAfcu1txRVEVedvs7IGOGBl/T/
zowqFTX9sL0ema/md/k1QuDIm1XWEJRW0NXLcMp+7uzycZ9tVNxQqpgRK/2/2ZiT
igosBjYQmI2qy6XXY+OklixTFsIIfaKyGp9cSK9V+BiB3/Wy2LgC89Ri/BSO+/Xo
5yUuOChBnlQBme2C3+rabReEMgOiEfxm88TvV2PEBCOgWZahd/Imoz2Wr5FSD4U6
8WOMHfnjPW7MWJhy6GzJlUELlMNbPlhgltYmWueKDnN+Ri2DTTwdWQElLNBM8CNS
xzP6LHjJUtSSGIW9ywCYe98iTUuS3bE38DfsLWgAoBR7DS/9Iz0ESn07mt4NTKsF
qFVXqYiUiGU+LP9y944TTww+8onncA7k3dz8ogEE0uhfoCkqcNysu9EyBzH02l+R
CQZvOn/IjgfyloytuIzc7PMsdAFi7/MxqFuRUplcjB1gswW8/a90x6W8gwbRFqXP
BwWBA19GcflRgYTDYJeWgdfZBznjo6VpFrth0oUJsl/ThQWk7WQBZ0SqeJXtShVr
oywe2fiEyzJmz/uS9OWeB03fv8JjZVwezIGtC4DFwU9eK2r2KC0qE4lpZByz8EQr
E/F5oeh2PRXIIV2cV5ICWltbqmRhnJuQ+4ubaK4fLAcIPmtQFMC4XPG7pF07I+pQ
cv1rsEBv/uyuhSQDaBpcCj1mlxs4ZKWKUic61PaS+gvcrQLe8IzLtLBCje6Nh2ce
YPo8ThEOvZz2yBRxoQktygQ7t1os0gxI0LngRliCudP4ZRRKbBohtjgdBrmWERmc
wQoJ/lON7uMCU3O0DBdUREyRYqLjSP//UTpocHsb0NSgNoSvLy7B4KpokWkdh/TO
SyOgK3wgjLt68on8jljwvuACLOOynUkMW03sKcl66x2yhZtg1G8Rxd8iXYuGT2AV
AMGz616q2Gie7vyO7ewG19R+JwPmLhfg+geJllp7DhD3/eGO00ujbkkpCqO22Q7D
i3re/I6l/7cYWRQz96XAI/X4YYZF6XnfXsWrYDYJQ5hg66RumUmzu6Cux2163SE+
HcOm0/H8xrRULo36cN54/VaEqnoYP7QiEU8EQp1bFc+Vwgr9TAoc11KuUgu5KvDR
Fxg3g7Ogs/WWqKAzhnT8jExdPkdWvmgFdBKbD5sYVMU9k05ASe3zBm32JLTN4TEs
zchLUoxE4kf+U3GTn3BrZiQoxT8id64FCufK2QRDyF6BsDOMcz15ch1oT1qazeua
pV3EAwNNT99djzORouruFneU4sccQQVwMJ7bstcpWo0XWqSmsgWbb1v8BFEIqDI2
K9zsXNai3Co+zKBlPrPrBiuKvkIG2AQ70RcPvMrvkT5ayM00bSRzSaK5XxuP0HDg
aedlW3UyECz62hN3kdxPuQmjPqRDr4NG+B1OBNGnsug2ncheVD+PKDt0yPC5ztYu
LTr4P7j4g1EJCx5klydN6I3Y115Ev2KtEzufx6uwtRlD/umFkNpRZTLQR0Vbz55e
8h32+FchpvsLRJf4BHl32RzLVIXKLj/dBs5Ds82IT4igAUfZ2IBdOHEPn4kYrii3
fQVY0wHN/BPe3jpJcsa4HzxfVdAy2uE5GSoxSqPOwbxSolsAALsNKQ+6njPHcc2E
E0Kpv9j5miMCSUitbQErX8UdwhKx4quvgYR6A6cU4eRyCt0nNoIO38Ni7h1Lall6
DfLIXVmwE6AlGNlMENqNLAHwBndV9UPM7LVugFesu0R3EuJm4+9p6zIjAXR2RAHA
xSzPmQWiRWaw4AVyjNy3pB0VYgEg73wYxCT3ZLKy+ppN16UHGgoy8U85BI2yBnw0
BM8UyisgRa09QGJ6XqMcysKnUN5o0gdjgc2VWIVzsjKrfnLMnYt/3LVeb60TzKjh
BpkfMtz7c6ELIYVpH0QI4uuUQh/k9b2HujGdUW4kAjAP5eyOBFdDTJr9vD/utWhp
fA2B4XkrVLTcFVMq0ayePr6xNR3sYcK4jn2JY+wLMmCONJMqruTFy1wPvvVBI+MQ
kxL537V/2AJJSpGU3bT6Yu9Is9oeNLCS2aypbo6ueUO6su1GvwGMHAxsjgRL1CcU
WA+7eBH5ngffmFcAJi8V1jBK473xo521pdnr+rqW8V9GDJJbCPr8885zssSDnPBn
aMWXEQ95vnAe6TdFXyKzSOzRZcXTiC9nfSSpyxbAzazYbrolCZOC1kA7s2FDOsMK
GCUb5Ix1Le9OyeZW917GEuQcR8NUCoFDz7KZP+LYJ2Iyeg9E/2jAtR4V58USE7hb
NPUI7Te0kPZ3UFPV1HrY+B9BzWxA3JU4x48rL0GYd9ipD2ivrCfYkuaqW7+ZfcTF
AHNBiCcPO35Ap6KC5qqXs6yXBDyILoHcTRk+4DslLsTlspLFGfq05gniHXDQQmyS
Uk22BSZqf9dGeBryRgjSigpynBZ/eWrTAg95x0tkgcQpBdoQOqaDh6WhmVcefVSZ
JMuIUMKmSlSe18FCshdNjZQbxeYOEslN6JaU1EWtCwBz3ffo0UKX+iLe6U2ffe1I
ZI+GTnq/eC6NLcw3oDQIiacCcw+a9Cxzgl4f81GRLk9np9oNM8Kgv37bQj387ro2
AMtSNUNLP3wOIXW6wPpGJNTSECHNUH5s+Jhxhb1Tohgs2vMwIvvd7LtGTMh7pub+
86M9LRnzY5hmGtAKlU/KHb0FFOq5e+4uWDNEz5laKKGJe3uWF9ATqmr1PdQEy8Ff
vPVmMsVeQDWhKpWbqtuc68lpL0c+c0npZTJ1Lpz7BaW64LjHgj0FS2UjytNt3dtW
KdkTzdYuVxQjIUxQgwbnznRD3BPhrtH0BVYQEsNSU5XgXAzdX5BIkQJg+2IQjeCG
Pr0A8EfQoaOKM7unyb+nN6MVSFUnSDPOrw4g6u9gcjKkDBR0zlQhG3skjycYy2pQ
xSGCY+n68W36KjDRgDJoJ5lcVlFrOmK1PSe++VrKHRg8K1Mr9AIykffowZGmrBhs
kQcUb+MVdTJNjCQoDcHBsgujxsZQ2g5+2MXEnJFoT6z9hROxAz2VuG8bqFR5jmtw
7Q2H75CkB0M7tGkj4uX+ffk+IXLnIqb3wKy2c3S/Ov/kKV9Et82rT0vzt9kduaRm
FNfuw7oDC0fiqucG+PRM0CJU+VMOj+QavcojRc95LofkhNUWM+3jlHkkO++g/SZB
DNBz5CSEN4aLxihGIa/mAGEtBYZ6IEOBRvCb13NP6NE0wZNFIODCOAhSTFWILjQZ
0pswvWSdKcC5m8JeeuVb9PmaeCLyNmOmg08Hr0rlN+flfo8yu15Y49A1FxjJeKQF
LdSTI9CJAjKFVjygpD6gjgOvoOezo6T+qv6T87iS1mlQ38X8c2keEb1lGNWKDmS1
/Bg9ek8ERqpKa+xSOAfuuL4aLEUu4MeKdUzee1BchifChdVpy92DrG4qi1iLqZqy
jw5XD4cCKNHos9x7/JlAvkfzuDj1WqIaSBI4TUOpqFqQIOOO9Ae/x6eMuIKxFUw7
F5jY8L0S1ABNFdrs8DbPDho1Z4A/6tYXDSaIzyWWwy8auwz7cq3aJOcBSRaQBce/
0s+fAnYUT1mml5hpaLVU+1IX7ie1aSoXGZNoXDexw5SAWBCqGYNJtc0t7i2ezJcI
e8MeZsAxzP+hYyE+0llVEjNaVpzeZcPu6FdPixpeKSCeMnHErBrIZZzDqii27BZr
R2+Qs9sjWLzwYQA8dD8xYdu3BUeHb1ms03RjVAJ3ZNyfQxxVhthVzHlHyXy0TAxO
4JVMZugZi744E3lCc7VQmEYZOOm9EiGxjDXn3w7Ql9mrAMHoDl192M3C4904aWzw
H9u6xNCYdIfNwAVOQ7x/2iFAEATM43Rg7xumN+PJbXENBwhloHcvk8yQJDOIG858
iCZItSVCg5owK0p6TWfxtw2CsKyoEry+Fky8B6J+k7U3LytXxD3xeJUt3J15kZ9r
6abuppiOHKa8csJrazMSr78o8ZLSb7rH6lsWWmEy/T/STe0ovk7NOF42iwNmNn4g
xnky1AHl3mOdwUq9/faJsGWatCnSo9uoqgw40jLvomtyextqQPnmCRdNYDKHUSU0
UE5Sbe65PwjuYf01iZr4pMQlhkh7C2HbiWe5tYSUOnYYqqoNOkTVFNcPiCyQXIYW
qYP6pMhKOTP4XxDfVl0KOOO6KfhIAZnpeVbGz/3ydOGBO1Cw5RyyevbyMlUsrGHV
SeRaY8JUXeiQWH+EX1I/GLG/PabeDCEGJV3Hc12SvLssYTIbvZ7cOH5kahhhoRmM
s7reI+XUwtdG0PhPZNqycFQSDv02vXnwGSsBo4uaT8lUrjrAydBrtmMzfugxR2b6
ifC6cht7sEPEArHSUd7+O7mQ8kRsi3w9p0uzECS0ivpsfiZRa1zZaukWcohqhLTH
C61jvGyJ/xRxxR42Q4C36IohUS5wcbyFWiYpuyxrAsN8+Y034laHEatbR1bfQ32J
ayNx+cXhqYsUBQ+wn2tc0ak4Re5dzJVHwMRkfq1pruIKkpLaBbvRwoQEBv3P1qW4
Bpau3QDmNmoJ4VA2E7hwRXk3HB7PQsr5r2NSyRmP+eg1TCVdLitgHhewsouGoTFd
9rJv0VEG2yaKy2M+ujbw0yKoCZ4206wpretQdvV1H0L2xPHLC6ijBwGf97nAVnHr
pCkLry2jtgosi1IVoa1TH+VpNm1ieDPFJckFJoh2SVjMcQkTpldlxTFpErOBLVaa
UfuVvEwdJTtQk2FXfq6VBdBEYsmX3MyNN9E5VuoiOncwxRysfh1nGhErfCth332V
2cNmfel5hos3vPo44zrwvyvWplH/UUAVbsd9YSY4NP0bEpML+Li198CSt/HoSlqO
DtQ0nJ2b7K6yecyDkhD67wbFna5x29i2wrvh+8H3z+I6B5UYdXgf9DgSV3DeeMlE
CMUNbas4amv5Gv1LZzxaQ3JN9OGVgjFjapJ8yxxbgZXmHGKrO0lEKLKsrvD4aJp0
IsMPP7eauCWVqMK1sJVJhqW32eYz9uUbJo/fXqkDBthgQpa4HBUZYquSRqs5E8Ia
0dHZ4Myr3yPwz5etyMYrTLvp2RAo2TljeaWZPykJ1N/D5jczoQtGozzQwosOC/NP
cIyCOk3vR6YT8Eld54o54PMPW3GOxGJamrwH/o+lgA6y6K/5YAH6FJ/mpS8iQbKx
rGY193i2FvkWSG6+9AOwL6ynSLowL5Gtg0RRTMSdd5UWquzE6ssFjRFF9zNEUGya
1r0TBo+qKjEKbnJopQhx9XX9xJ+DLW5lf70AxOqNwdWaLZ980XoBZvgdTEl28CwU
MVNA/fX0CKdmqBhu9XPtx5cZeh/yVurtj/zWZtvrd/xB27Dqey0sPBRmvBKrrh6R
Mxl2wGrb525uSM1Bu40lakRKsk1q9H4uGDrUXKAuwjpUWUGs5qTovrZ/xN69Yp/L
JEKBRdcL/6FepUUNFs2UpCWVrRoWQqEMYMMyUB6i4JRQxwAE18nxoodrzt7mWmM3
s/FwCVzRItE7bCFqp1p9rAyBwQd0jpHD88gesxJADqDIAn1/beSA+Nj3lFTLAlhM
eJ/IacTDm9ydZtuid9JndT70nZy1zo8/71aP9AYocTMco9tqNXqXj/fDghjZMSwv
0vLUw32kQlDcYnb1hD6LMEfZdQp97wdTa7znOB9a4BbLfxAwYxJC68ae9SB5ISt3
joWdbazXzixeQdaOoeacFMyTX4NITp8z71BlmCsDuDLQ551Og/d/iXmPPrkZJ7kw
3QrbdkpldxmlctCkzn7wQVYuoFJCQOIY9h/t7clPTaSLIYwkFEgWWZ8vTK17k7Mq
HCPkArL70OC8W1/EXRSNS5qj+KgLlXg+uZhmteB7I89+o+PQzL9XD7XWLuSfyH8j
MlZ5CTeKoEd4+yi1KgtENxwXpAR0WtrU6W+G3obc7eFnYlWXu+AKfNrYYfFHYr3E
u2JVg/EyKAldQvX48yUo7GUB+A9TkjUiSUh2VIjIJMOsI6o5x3qC/s4oJUReJdHy
FlBBJbTAL8BA81jo98Y1rORiWoVqr3c2tScXK71PP70a+UhuSiGJgUc9tQaR898k
FZxpRCWswSokkPOYa9nLisUcG9Bfmo1p1MTDjJ2yukifuYrok2+ZiEMLwbIt5C2w
DkFNzp2Ahd/OkQyrgxnN8jFmrbQklUln6mXOiNE9ntygOnYb58rcRz0EKwOn6xPb
T5p+8vBcAHwkO6JLpsEcQRvRqj3Q80zKfmPYN4OWVg7f4qKdselRBwvoubyZ3Dk/
yjsZL8UtTyKCHM88P2ZK4h26rD75+Vrywl8fSBz1+ENwiA1Z+JaVWd0utlfUTxEZ
ROdA72O4crQcMRLvpYzzr8td5BrjrzjUkkbmxy7bL48gRoiPuqky0hkZxuHzAQtp
vnQoFjOjaXjHrxvPtZsTJPJV+bmeTw4h4i3m56Udw/t6VSxnMBNjEpP2WyfL3SaG
DJ/y7TvDtGWD13HlIn3bgoBI1RPnyYbCz5C9brQ/fjtNLCkcCAmXuh0iN7t47jto
i7EnQzb5MFUBUu+4yom4yp8saGCV6LjUEVzKsFp4+oQzqW5wnYie9BNOtQ09WK9P
23Z0GVpWo0RaUjDRoqS1zAioVVwyZk/hf+l/LSJrQhrgbKM9LipM8GF64Yym1olT
tMWZi6foZM7Br6FtHUX2vcXHCDMDTmKFZhyMtJmlJ2W0j5WdXt/73lHD3JBimTSH
M+ye85JXDnC5H/NpAPFqmRTKdgxFNawvlshh1E8NDMwyWMDNb0IXgGmPk+WNql3a
ws8ZdaT30RbqjqfsjVeMPopqLz5UPIIgHgxbdz/TPKNXqGhmxg7koT6yFhh0N5kI
1ZdwgrOu9DMNSiAuJt4fBV770G6IwgFRajWzigAkfsDMtcrMG8LQrQH62R8zQ9Ln
+JY9hU38rwoQQBSr3WqgeW7X4gHnz0/4EEON7KcLGBCM0WPLNWO+s3QGXrwsY8PZ
Ab3kYcxVCBt/EQC6UcAotzMcPxm03sy8TzoxnVja2Q5kSJJCLGimDbkW7FV53bs/
wDq32b0SQVPVjgoMp0wqzpJe1LvWNTl0EjkLHXdXd10g70yx4VuyE9zK1hQgdlsW
h+4O/1gtenrzTeG68sjoRSfggjgvSKWrlVf2JzF4vwHiv86bq/Wz6Uw48Tscwvzo
6hm971kQr6wqHLioM5N3m39EMlFdVuH+yI5ltKLXM92Sq0Kt9fpfyID905A7MyTL
yXCJiENeLtOtvWtZETQZ1bGF/l5u2FasCBflOXfepLpw3uU5ZD+lRb43ByCwvz/l
BHj5Zex8dea8if4JVXFIkb9xVzqmzDc/SURl5bN0ECOm98LPjCUQIclkgsq/s5Oe
lcRQ8ReWssLdvKigtY8mi6xDDeYX9vbRgDdsMAGXXEQTHvNlaMIH5uavD9E6vaWd
EGHaoKwivqxY3gusRwrCiHn/COGx9hj0w7wZa1kaFgOex+vGEbpeFOqwtOGAHSs1
LczbjJdiU2rPeHeIc7cUN4qXcmGFe4JJctiwuWIqLXtMlayctTwL9iEBnU0ExOd0
BkkJF5TyYEw9MyFXUNduZAsMkChytcQmlCS04T+mbVLwnxWiM+a3pSbDBbHG3iJo
YCN7NHxUVczyu0fbnRiFYFtOaPWFyBrfwJh5e+4JG+Gc2b2QBB8aZT/ubEgdpCUg
qQRJdgEa/HiTgyaNPUEXqG6f0j3/adSGTk1Hv2w4r7XNPT3WXRraNTyNQ2jf85Zo
nzcDYR4zgwpVxBZbBY341i5DOu9K9sxVTO9jpxPjwK1QuMb+soaSJRlv/P0hAHEp
sJtv+LdQloKguTvgIsfFkqB4VrojLzB3pVlDYBkxLlnvER38mf+nCa91A8i1Yf9l
RbbzwMC0QQEd0NltQ3g36A==
`protect END_PROTECTED
