`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7VA96IuCvG0jT1BT0AxfNkbkYTx3l3MWPDlZuJ9s9C72DHuIQn5nflgHDZuU/VP
jsRKGU1pt7qgX+gGTtU5la9I4LomoWIrVKDSs3Hw40ox/0n/4Wjv0lmsiY29iYuF
Zvld/xnAOVV7A9xgXjLooXhmzB+i7w+IxucHbxlO0MFy1Jqa+kTHoWoBKHMjdwMa
3SWMPW3jHhq9fwLpYu9bbpKgchrerSVzMwP0DkinRBh2dBR79ZNYwPYpS7fqM77s
SyoFQdrFmpAdBnkYldJlKFAs45SvKF1o02eSd9hJTK+GKBG0MNe0evbicLWIJMus
eDi9KjwVXsJ0IbQHhbd7mMNmkRLFJ/yPCeK6Xyky2/ouYkYxBHwn4spDk/V4e7sR
K4dCBn1eDPsbcfZE7riqU+N4FPJfwkFlqVGi7lqwW7mYKWwceK8QQL0ugKywScjG
fNJHrJna5HuWYQCkni57yt6mhDcZ0pIGN76Miql9hF8=
`protect END_PROTECTED
