`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEpkg83DTF/jnmFzlDSsf7yvntShIKrkzn6g/TygqydadUNzv5+gXjqanW4Sw8tC
fCoIuASh8YADp4mOPAWA8IJTI1oDXW/X0BCHUhuoi1uoJXupHVc6BkT0GDleVOKG
eSigdgkEi3V3Jqd9gdsu8BFaoW7hXLmoBjJiJp0gnKSj2clDZG925Ezym57+qp6a
tmRLMvw4XAKO60vSlXc4lVPjRZV24D6Fk+iL6ASm3bG1Wu0CmjQXbMhqtqMeoCVT
4Gv7LKCTnmGl1nw7Q/UeUsWla6/JAbXH1Y9ssdyMonkpHKJinxvXZu/tTjeyXe9T
Ioj5NhfASpQ4slfzeP+s4EPos103b0vHPCVX5nhgMg2as+Hxkb+WwtbVHrQZuHj4
kEkFGRJrK6JstzG+qVRGw5xGHs8ZKb+w94s2bEs76MSxquZSXufK6j0D53dY7dEd
sR2+i1qAyM+SqH7tAAieA7fnj9RCoqCPnv6WQiGurdEGAaOAFGua11WTX9qQdAmP
IOHUzXR5GXD5DRthmtEgCT+nbwPpVGGChkRiA1BSj+AvO2bv9Zn9WwAqfILE8F1h
jNL8c8A8bYnRM3Rr3GmArqZdqwGe9oaOAm7DU8PVz+Wuy31El88AQBncks9KbyO3
GgHJpfqXamKTQWNrLYtS9iyxFGXPoHgccfsRG9xF6cxa0DaDuGf1p7eaKFWXREVy
cKa+G3MIr5qnSEwmvDBrXJRHwkJX9iIRMH+XZfX7h9M9vkvMxEf8LirsVYr0c/b6
bRsio7ZS/IknbN6e+n8VoRsXA2VJSBMYP2Qi31ylO11U9SFJ17aFhmhAinXvM5Zc
+JmqYdVBHlixCtaL56Sk1SWAmQ85C7b2ZDVwp4R7S7e13BgoFcr/6KdXGkrYpKsj
7RbSvlmxTwOVp9mU+pWTYYEGzsGQCjm9czM2ULY0xqPVkXhSvhHwsX7MW99+bG8W
uawDaAf5PmiaKGotJvmaqULZaz65sTogQCbDSI+nBK5gKmZjuNJ2dBDl9TOQaf0U
U+2XPJbtSftbNwHvJuVDkWLHpkxW/rW6MU3JJmP2fBCjLOYM1Mzng0TBE6UbY4GD
Vre2eh8IPAYCya0ZKNaT8Ikl3JVrkhCnWM2ZJoFxA45WrEor/E80YBfIjCcwGzYj
UzIQDEUo5E+4YWu0/RchzFrNnzL+fm2ssAU/wgmKfjkwQUc96NKKOrxMsRHxqp0E
TZKrl0c9TgizU6aqPv6qn3IDIMMD7CXIbJB8BfGXRds=
`protect END_PROTECTED
