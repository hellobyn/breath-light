`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3e3WljNSYzDPbz3ftYGd5u651Pqy5MO8VK43zlmexyd3+jWsC4HHQLrj3gktMhV
oGUD1yWqQ3/YqFLQLpJVqmKZD48Tfc7buyJdGU9Z95g8mdbNsxn+bpE3gQohT2yL
aiKovr5pwkwJVofsZJkj8FInQuF6P1trcMjjB9G7EgZaXMVFqO9IV73GgA3Pa0M3
Ot01WajyJDmvHq1/DQtzvz1lJx4dGHk1f0BO6IgHY+O5f6gq98zEdPTGVg8yU4WQ
ybVZdBOnsEwYnOsQ2lkxaemYS7hVlOgXBk9InqS085oieAY8YrqkSdqZOoiKSics
EJIqn8E0Egh+pYQH3apNT9svtYZkXn9Yt3HThrIdb0NV5cEXVWNX2mTvUdsHDhqH
VS5UM01zfGt8kHvSVqBpNGeo06IV6um7CaO4f2NMgJESmtexITTrpoBgTNwSSKjH
m1MsuG3U22HboEyVK90cim7+JTmbL0AGbVuY8UA7HQSb8XBtPFbiJmXgt/vT8R/Z
KAydPjiZuaa2vBeFN8XwHzi/1A5IgAtUDtcqftjxZOn/bc28g/lpQc0iGF1rlhdy
AaIXW9obopgeb6wDVdc/msGWqRZDOpjTPztVVw8szDAPToNDvg0pMA1xN591Pzil
OIwOkmx+/U7K0IAajeVtBCiMgWCEsNckVMkzovNiHhee95ecxOrU/gSZqPtZlbM2
QrQ0j4sUU64e/9fO7Ht8VM0JtoTURrxflSmw6TQgj6f0u0l5tolTwE/TwlFU7siH
b5mL/OK/rhxO35AxC4HpjlqGWn3lDeeouevnxssOEX/OMV/VkAwueib5DivHhBp/
5LTA39k5oOasZv51CJALkR2kIvX0pq9klxF2vwcjqdhdJ8pynzAS1cUgevUthmQ1
yDClY96BukQfzbo8VRgnaaba7knJFLNkybpkepfnzLMTlWAbc9FWuyAkBZpfb8Z8
9ZlwhvgjL1Bc0nL6uy9pMpDfZdmdzAnAkuC/Ydiwv3xjj8Pa0VWi3LvRhDhQpuF0
TuMtkiH+VL1eALDm9IYfze9BjQvYJJZgoX1TRvqsaNKPsxLZoKqVHyvV9DuNd65/
omDbFzu+7/3JlXErshcm3mt9Au8xsEPMOEC5PEre3TwMfOAwgNBmiG4M1IWQfwI4
TuDETjlOrDw1wFJSu/wYSBL32xlEfzKTdGoAQ4KrICI8QY2BamtSaZpjR1+kYCBW
Z0l2qMOmIKrI6UvaQXl6c2oecXSA70rCaHwnZ/prtucIL+o93mVoYUpwZXvvytJS
6bl/y6YAQ73H/GqIoHgeby2lN8BHC/nC3rQdHfjaitUDG0K9tIHH223OCcSLwZMy
PmSYQgbvHIwULEjjCFaWs9zqiiq3D+g7PMLn13X90BljWap1atRl5QNFVoDIT64A
9XRA9n2S3DpOTeNymYDbQtmPg/DLaoq3/chcSEkdplWn/cP05HwzQ4cKkFDRIBJJ
57RjRPxHpI/ejd6xmTNBiM1zdBpGOxH95sTqP1+4e3sj2/Qdrq0d+/QykPr74Jb+
cArupAft9HCliHM/Kf0XDxjGLfv0KEusZM7fP+30U6eWO+yxeMWqkDO9Pdu2aZYq
+jbngrs/wkI08h+5tNEtg7GFU6F5PDenpOgW97JplACXztdhFkDKfwxLeZ/vch1N
2ZcVzSZNHnQBo69QDuvqyaZOzLhqh6KzLhU+PCKSksJKsmcc6eYiPmL29+H/w+6m
oXO+g3L/+clJY9pa/zuFfc79ykJzymU4NWVmWGu4iY/krUjf7/dPYLcpXwLFCBMh
9rZWDJLg+eorBNotNdRhUopbdYbi3f+GiLnjURCLiUsi0iDpN1GQw/HYnggmD2Hd
JPMH5jMAgT2EL5m0n9hUYToGmAchaBC6N5aRAnQDAqMyZyhl6W8DJwjScamLmEpu
tPceYrZ8vZb+kSBEh7hZ427X0kzmPYJoQ26Nkl4/+CJMBMD0dr18WN6FNXaBzlE2
tZmjGyEwaUZrGXmwduCut24CZ5AiBryqn8p1Bi6H100u+s6IvIFiHIn8junOpq0F
PKN2OH+XEvz7icqm+DINlv7Ts49PbZAtF93qTheOc934wg/mNoFDDlOn+Lfm812O
vEhSFXMC4ZR7eItCQysIxfm5LCBJVUwlUJh/rRY24CJaT8bEDjjHjgOg9TUsANQW
bL0LVCBapw/lqSRpJwClCeCz5SvHA/hvrGa1A7MpiMdUnWS6uUHlW1aU0EK5zde4
gA/Te5QlQ/UFIY/KVK0fiH2GPpPHTTN/Lcx3a0sy2h2fv0+fbTXfd+2km8xRBPpE
8NJ4WyJa6Ez+Cg4ey+dYV9G30r3gNYhxugkddHmljvXwgUtkusqILlvxZrJCiW77
rvnmPqtdXEiUtsOOBmgUxB6KnPF85zJJ+jEM4qqzCwncCPrAXfeGLz1YnCSGa1In
6aS8zFDZbOc2MbaCriVIoOvOkR+u9tmABYBrAhrcDGaiHuBGFVBJC1lIsKRW88k1
DiUpsc0jRrsCum/GLNa8/SavoA3SBjprnMKpF2xChbwj6y89H4TZNccagxa2bpOf
5EtxAo0m2MBkoIy/DZuJkT+6rnq9zuBbF8ljrEMxbRxTko5OmNfZg4N1XaQwM856
oZM35dc3yRp1bRmZSe/ithqXrZRXzslmBXGubS79bfhnIJw6O6IIgQEJwRm6qfkG
ILW21XnJXRMhf3v6eJ/FiOuMQXlBRXYCA35NinXK4VVWMa5TKAoeDOrvfRmZwpUo
qaaldvat5ObZXRaA4Kx7IHghAe4DzeAaRv60SV/1HkL26PY+mNHeZAqTuRuLuPTG
fyU5FS2NPC4cy0rhECaUo5Vv0FF4IBF1/dtGczkyjDWTIV864xcV+v5SToT/rYDP
FFLeX0HA4yWBssnEox0fvAV3UBVnDInmnALzkfmPMYKNVKS59Zua4ecvKWz04Yx3
MoRQFeCqxRxq/KTIqTX8wIUJisrmLe0rBuvZ6w82h3HcLSJgCiGChGB/VU8swRVq
oYIxP7c1f3C0/WUIqOOgPWhsxS7fia3jpsUR8kh89X1hmchEHnEtXBX73Hu4I6ps
DbSMkFfr6jhLiIRabaZCX46UMdqYY8JqD/Yx7jToVakot3SoMmKJ1laL5LoJdhcZ
qVoVa2N9gj/0QsU1805k/60znI5ovQKowvZspuTm4eCaL69e9GzP6yE5gYDiB4GY
VhFQUUlxQRcvthN18++KDAK1BzoLTJN8Z21PR1J9yn56n9t3thYJSbM5r7rMQa1k
xzRnKICMt9mDJzh49bzg6tYB2FaCL21j1/S60u/LZfPAZ+ygfvtLvjB5rdOr1mm5
FKwacT69wGAIIhfQsHFU4h9ltG/0YjLyterHLLhKC/1o1XCNXgnuo5L1XhMp/9E7
/98zWsVhQg+R3bnCsA9WpjnH3c++v912k5jU/wDqeRo6p4IYACzbV2GLLNMcYxOh
+8310E7UgB5bIHyt5Qx1urwUQeECaYjYPWUAK7cR+qK+mT5P3J6J9xTlvACt49cX
rXzIVlxCfzruTWrNaOVFMsSKgptpQQBXdefABPUXuSRPvSnrmFuQu3XL5tsj1+sU
j3UcMFCMjHwwsrr7/OBKYkJQKhpctWWAYgdKWo2KrEsIgPYVYS1ybTgrGwYsrTVt
5pIZfxyafxoiZmiuNSMyh1BeCLbj+7wK7quACsI7/mfzwf43fRhRhUsaYH7l34AJ
uSSmj07KPBYcG2p2u6VSfoeI4SlERRcgH4fz5/bf+hzmvddbI2VuuIz/q+WvW19d
VO2d4D9DF5ikeEHFPIhxXeJjeWypSl1wSj7Rm9XDhrIDuErAkVjnQMOKcF0hkbbB
KzC4zkgJE8KYGSpTJFA7cfA/xvwWpyl0kmd4HSTIFadPow7STw2J5x8roe0s9e4c
KXr6mkrDUOgyMPLN4KEhew0I+ie/OxW2Z2QdsECKCQD3DGLDByYvgFESgWwL0xmP
ycLJoXJWyIBwFndT1rakRw7r8Nptw7fmaCSDSi9lc26n8upJXV3UQAPrRcNpYZfD
IJesywUz2w2p98jj1uyxm+VBqvqvjE8xC2eo+cao8zP+EGES3fQ5RKtOItBWA081
01SlyVKZxw6HCT6KyTWbiyWxs12O8dzQNoBU/NfPEg831fAbhrQsVEe5463UmNB3
GPRbhmzqFuDmtSn1biKZg7osWPhrKhIAyU9g5Wd+C29uQGQE0YOpunbDq3wuzwn3
UGI2cmW35N1JgQPg++8qRMzc3MgQwsNnbofY6V0Kcqy5uvoROe1OWUGmFncNK7zr
Obky8aAvuFz8vTgAMcLLGcrzgqJxJfaGH9OXi1/hfp6Q/WoZw/p8K0quWe+U71yU
bOx/Z62+OZf0UTgxExfq9jaCdjBNRwNlORM6tQptJ3G5fMAClPK8BV7NwRWxQmlu
ndNs7dYtITRPU/RQ/TXf5P1o8y0vxaT+eCESFvOx3VyMWPiKvnyzJna5EO1M2R4z
v2rGWRYPBthNY1rdh28Y3y9wmhzmqjlUing0DzUZbwEfH/AV9YQYD3EVYxSlHnMJ
T88exQ7tpDqATcCwagD9xDzC/+DEEaIxTc0AgmKth9N2C0m7tSatibRzbHuw3dSO
AX35Vnlr5la0/FAiU1fI9hckw1eaw3SBfndHIZXAysHImWAt8zxZ3H36brftXlJ7
uzwHXSkSMgZW7cWStmm2vfTMxYbTIYR1xlYonLXj8Ta88xxr3xKyfDOXwW6VscHN
KxOuP68AwY9LBuQd5gcUBTW0E5lVtjzQYxco+rMWydvra2BObZFJll/TCdzzRfad
ZjiTDrKpJFP6ORrtMr7ZVRvmuaysg8N+gCQAe97zwYH5ZKjugCwb2lZ2PQEIkVYy
xJfQVOP8twhmgeoK0PrP6fOaKIKep5d9eWTHBL9h/UjRTMXIR/mzJzTJzop0dELx
FimD94/O3Pf/1YnWMVA7LK0t/PxFNp2shv41IfWhLWwd9q/u2USE2CR+GP0T+7Sw
VF4Rs6e/5ooC2urp/SsEh6HZiQNQTc0b9T6XyxKf602AA2C2MdUHSD01DjifudHg
B5D2KcsKCtWCFSHzDStnV/FByf2oX5YamOl39+PvTkzUOMKmgh1G+lxGWKj9VEI3
espEAPCr1Khvjbw8Q4BVzhcguF42Dp81AuQxHctmT2W6T/x6G0SYuJUYnpKRvkdi
JfzytykLwazvgQfLIKf6bc0uAKNQ97M+uEimbE5TBn7CYndCN5Aya5kfIXzlB/NL
5NheAOzubmR/micqsb0bXn4vactMn6tKyTg7VIQj8Bp9WqhT5n/VPk5wKOHUeYwf
cyrUwfNyUS/f9ycvGwSMD1AZybPycFDP8/1QKFgww/b7A1ycC7ozsVdOZOPH4xz6
1YeAW7kzN/TUP+XJWJ4lRhYgGeW8X60GEQK4DOTK/4A2Gyp757Ry4nmik5j+l5a5
42vtXK3yiUjNU2X8uFOyTJwFS4YWz8hsigzHX6F55Tc2ezFxvfx7KiLVqCw9Fk9H
qCvo9dItk/YE3EzvOiL+k70FaNUe3QdsWYpQsfs/24HtiN2hjR20aHYPTn9qb6+I
G7JemlmaTIeUdvdkLwyN8IMGzumrT4HVKuc955babFE1IVDt+DWotMNZZfkv8Q+L
Wse1JYX0jt+JbL3wAKMC0X5L7vcp/7njFyBEXRrFT1jH9w8D8OAfmfIl6NO5Itc5
6nBPQJt+ZoOVKPTp9JmvFt9FlChsfiHq1t1+pzj1goRwAjc11M5TgLDlqWcd04bH
ccC2KLC3WBdo3SHR9WkDQBgHeHSWH+0dkqk8lMcbr/OAD77WaIzAXJmOnXWV13Lw
eI0qWx7q89TgYaBiI90DUpcfdCa7jWy6cLE+oelJYSNU3bd+kVKRZDgOdfECqRe6
+MrOVk9Su/ysPmZPfEDB3JcEM7bjn6oEF8kWs67h1Xbjynz6bI4uCX0ngc4Nv+MZ
xXy9T+NSyTtoAuOCssqalg5QKUmwL8xOkkQ5chi/fJxp2WVxgIOcQTy9MjbdR7o0
f1uBVr9VNPOtG5Ji+/Bl0TMYFAk0KXVyppg2dm8a0PAP9eYpkfZdvPkqChZI/Q8W
6sWSs2lkpPyp/sc1+mC+B2g5FVdUDiCdFubBEgHjRZ4ayhAtFhCyRY1N3GFj6jnf
QrNEpXvSVMPXluucY6aoVokATnL5QPAbUbbuJDEMjHEkJbrgRY5J51DOJMxs/AQh
fUPzUyBc+8x/sDd9x8/7JRyQrVdt30plkeEfH4j4eZwt4L22Uw6ehFYBjxJ3feD2
8W5BKukJQPGkpWguPIlVi2yEo9W0re8XkuidiKKwqSPvBShWOwIWTGK4nJMkx0Nn
9HnVLMHLzRNaVpZN3I+O2hOMqXqDRSOVXLS6zOtS6XO+6YUYulk0JG23vF75OXWE
DE1RtAzOhgTyGZC3xSGF7AZI9nYON6HfAJFf0/6RFk9GS4rOtpWNsTNIYJuOy1TN
E2eNeFd2ZsQtA+Lp/ypbnm1c+foIQ3q/cK96y2ovIW19NEJ7p/fwXh8MAIP4i3BS
Rk5+CBmgxgPCUg1mRSIcXtSepFCcAoyAQz1CBkxa0IklwamfAUiR3XUtGXIvGE5X
yoUwWnt0ThO6vWnFwRDGM1gcIdyUlfnyxFNuB4gDJFlgxXC7wlQUlB5wCaEFrffd
B7slPotjCCkUfWPkG43DKZJ/leezcJFn4HB7hOIyCZbLIH7+9Mv1kAOtLj1iYvdi
yZPy50Km1s4g5omk+/FGswEXFhWPU+32fC/wfVkebNm/SqAy2NxaGn5p/ZKdna94
afee8BskTHj6goWEhPkSDlM7XjYKI7obD5rSCbW5MrGdLhuzpbTrtQzuUpbvEMCQ
GvxDy7qL404EcXTshwZR2WJqzC5htpttjwMtFidDxUix4gCywUd/2z5zULvnCFbv
dbxOwCC7ixNtpdDgs+sTPq9MXT3OYMGBg43sVEl7S31i1KNQU/VUFbCMkvp9k9lz
EnKF/jmNZookVxZBwmqr+5+ywaYrtIygvxwPxTew/0ZwMU2yA5BiGoB9ktlELkI/
mSoYIqk4BermtvKfHT3mmFPXEH179iZ1o6qdRYfu5XezVPYIz2wsSjMe1UQH7fO+
9LlJIlU4gwtfOrfJ3Gi8S6HJmVQsyOZLn4rVh3dH+bEBe75i92qN9GULOD8fAbkX
YzYKzjt42foA+jI+0XsZMjjHeD0aZs+Q2OJ3ddwIXoBqR1EwYdGQdXLNz4XXSNQ2
9gCjjn3qykKqXE4Jsb2FHMeN82S4WkgA7qrnSldbsAghgL7j9jtFbufggIGNecdL
dOu+2i3AyBhXqg8vdgRULCpUkyIxRrJlUkz2j4bQSYMBPohEeCaKYuCM6mEtXRX2
CgmST0DrWnyfKffMJOBbFsVEClPlpbWLNTs6zCBOWfYgHgS27f4yP98cwNYQuYWO
Rmv0MPup5xBIrw+UNuGYwq+tQ9GadbHRm5WDd0Z78iRtdhYTIMHEoz+HUgedAjLp
dlabO3rnIvlk+R13I+CIaDwGb4e2YqpAsEd0BP70aRANkyq9Hjk+g2y5lJzvaYMq
qbmzedqtKCOircDINXS+zYYQctlPB04GkwGB76SkPLY8uHO24FupnOM1jlZ+y+C5
BonFptxWMT8UlRc2gzukE+mS3to0i4uR6eU4NJ9fOrUxU2MgD5Jz3PZcQuGdfjoS
VIyIgrBVM8GczjnMlYvmEvLMfYmCHyNTO89JqAgyq8OkmqLTC9nfTMz4ZYkvVsmP
jrIxz5Rt5X0FzmE2vgE7bkZcTBBT1Xg53I13AgRTvu7tQcWjnQAH7iRnP+eB/HHh
qQVqH3Nm/t2zbYXfGrcJrKYtiDRql45NW3WhIwPneCPLyfp42+PIMl2wO8L6SRFp
dvPW7PF7FRfjfk/OvEu/zmF9HHM/ATs94G3V7e+ykfofbZRKT8YUo2yUM4WyEeJq
GLdf2uJIt1SPy1jb7FPBSZBnSAsi8P9SUR9QzRHfPoRAVXHA50LlaizG79dZv6pz
KXzU0lRib2+IemJThWbI4PBWujSMn3cBtDDsj7Gxun4TV2iSNc7VPxIKO5Fm3QAw
dZCI5K4w7WuYajr8PTjhFRY6VkH6xwxgPFu/Cy2aZ/DGrHBsTSRXb8LZ5klQmrrp
zDvp1yx1FePWJ2+FTCKPsfGG6fzk7P/MyH/gEiiD3DJFF8U8cI7fGvSnyOH8DaUB
ADM7RZsJ/Yy2EnHWgMqeezTkMsccZ1WGtDuDRWaidf22j3Ojr5jAM6npThoab2WA
iaXKuTyUrH8K0M101OQ9e1zejFnLcaw6SidAHXB6xHMYTiBknECeYflFNh0HNk4r
QrCVUmFKp5aM7HLgHpAkD7/uB65Pi+RnQFYyahvjdl8pBnIFqPMmfZiLYi77A/RU
Nmgiz8YGuCidIfcF+rLnFegtcAfXKAFHQUaNLYCCoC+SHomtc6NJE30Y4zmaXRDs
xHARGEFrLLD2lF7hF1z7f1rbT+DqyxKPUXp8PgMfVjDoKRSmyiJwQ0FQCmD0wMqd
sd+u0nfdmcTKb9yDaNN8XdprufnFFqawRfWTUk61boHFE7fVFDEeFPc8vabCWNK2
OUyz+HxLNpnYaK2NPfq82FpxcW4Pp7GJoujt2S0wlLLcwAf9+qkAe+bLp1Rq6Yd5
IzB8o+hF9/gYJLM/QKzCkK+uc+LLQnJRQgOiWvCRnzvCtzuVaMkYtZhq7DVqHpdN
vr+iQpB0Ssa8eX279ESWD6/J1kdfdsaGbW3zm4g25AORz50rS/91VsdQZmTQc27I
IC0fZ4rVY4kYMhDoqjoVecIWijTKC+VmifGmb1jvckY4CC9P3I1/nyJbQdq9m+co
HcjTfidIQXJqCcPG1WAfVEokHZK0i3biVBvzB7Uf4dM65EgcG6zB0F1+4VD4iZ7A
std6cK/wNtWvr8q9PfrVFsXMtJzG9VjvCqnBoXnB74KzAXKdpumEbPsWTJIeA5gS
8Wl4fUmITNUNvSWO6amM31FhoUd6saw8YeTw021dPrZrGBXdTL8nFArppR8AeOVz
yRqPND68q29ESTwFYc0di2E3ons4iFQWQLOoeiD8VZ+cJHI60RQmb4XNCJ9yQ3g7
u9AOHcuErwxvJcWiOpMR3CJiD6ZYsArF9oJvTmnUT2UoqOVcHdpkTxBWu327imiO
fWlZ6P0/PeZ4QX8d6HmUStlXsEllOTUyhiJadjLqL2I0EFUxwd9AsDJMVWP9tjYd
Y0dDsGM/cZl8yiP53p5i2HEEqD+P3y0EJFY9nqNA4OAGUPkZEO0G+h9tOU1tU/bk
zw31IALlWQA3EaEfDd16VvZBJQ+ClMzqsCf5VbuOnxvlmwnPHV426Ktbr0nhjKgN
5n2EN6RIPeIF4OhRVUvkIOewBLdynBcSWaZs0Vu/Nq8cppOfITj8mLCbzgHU3wob
qqhJlIbAcmnpK1f6Xp4rNOK/voTvZq1rj7lDA5zzTPfX+Aqxmlk2uPSn2DnXilop
Af/O1KeXZz0bHGVLb8wCoOgUXPAtiaooasxq8uZUHQNgyqGm66qOMk9Pcb6m+bpr
F1x1U0xaRftHL1Bp3XpFpY1P1RgnlN71zHcpy7L/qLT/umMyTdbsd+jbQ62CycsA
LNi4515Ci+Mz3D0VHJv0aR948YCeDJR9uge99/YF28SDWasfrRuLdO8kfp8a2hmk
BUQk4Bmz21THVqoolCNrgFR4eWm/McihWJoMBPcS/MxT5jivEIl9zKtLfpgxqGOe
U1VQkEBrdxLApqcq5eA8dJ1Q8Rzjlqs7rIokZ7hxtOFzvGiOS5OAL+3a3E3/ydD5
BfgZPpI0DNRSdAS0RVRDj/VX57bmVGOyzPQ+eeMxyGathgk1ReFpqfwQHsy0YiCx
nwUgJD7sv3/bIMMZFOLVa2b9HEiz4ikB9x+Nbv+766iQMXaxW7HiJW9DqOOhaM+U
tNN67AwifvFFHmEygRKbr5fD4pHLuWUnAdPYpdQyyqcVr/T5L4wp8UgizC9kG6Sg
3ljws5/BsctbKkEaLFzTL0OzX+NPoZSMawcAXyB3WsMs1ciY90uMSKjOHXSRDjzR
/GpsA0MnmtWbcNpH4qfBskSlAT1s+lEoF7P5laKa0I1n9tBDYOhiF5GGvhBGBjja
DHqLalUVMxgUnf8EJg9uxeeCri4CDE9gVwemPOIajjvU6DAz2+iiJJsx2lRPsltv
AGSYfHdL6VTYtlKhQ08ZvZbfIf0jLfqA7X9appQVCvS6aeEEGMAo5H1I7kq2L1L1
gMdgY89Pr95aic4gXmPkHokgS3dubCqY/xo0wk43r/UUlKSsI9ds4J31dF5wXPbN
V35DmybLQw6KycnPBIbgwh4V2QF5c2ndvsvdTmkWWDLD5Q+0eCpsRTE1ZG8TX/+L
1JgKEnaz/vfzin6jVuXEj4fLkQzxTrAqzap1yxk7DsEwci1RrPirpKHyFQ02qmZ3
508MwByASyrUD9+w45MD/JDcrBGMP5/xNe0xOmodwT7q4fDSfCQi2bfgCqgigdqd
lUUEeMc2N11WqANdPWVpPA9Efu0pdjuUkBetHCQPm4UCXPbszrOmsATpJDlu3hTc
Q669KgZy9Xdx9UGQkIPPT0W00jPOqQqiRWK1V6y1vC5xFl9wN4R+Ilj6q/439cSY
5cXYLfmdvym3G11TGgOwTIqmYucf3K+/6I2IgsaN3F5KaJ7QrdUyFPZQOlamaIYK
PtDvVBkWeQUOk6aEhyLhIa31L7U4G3yNSsyoIzNqg1SdltORzQRMs1bnipwZBpXz
BevHu9GnADJ1SR5Avb/xWavnwC4rtJxJoPo+YOcVhA8kw1BB9KTsi1I3afIiSZpY
v9UFTGmrB/mJXRBmlx2ELNhUx9luJg1Q+BF9/263I2TsDzpe5X10Wc5WU22hzbJg
Vh+iqaCf/IchT/Hw7KM32Fpot8SDFZDTNWQMr9zPgZiKTy+DIcMIdBb+0Qx4kwFa
6d1R4Ki/FNYD76/y6yUarqpNW8VrqgUHrsSPYEaYbyf7AjgBxiaS1gXsBESRpgBo
p1mGAcODEH7io7PEvnMIQzNABqCxwF4MMORTDdEd38TLlaujH5YcaYirm/xzAXet
0a7FjV42RsoBSMeAYuAFNCvu18a/PGzSrRzN6WQdWNBxkG5DcGqzqvw1yQc8RE7u
BoZ9pa1YkmuY5G/miVYXinkIIliijOS4XNwz6Jq7f1lrl0nFXhS4L99mH8eZnn5u
WOG4Yu+iUTynjOJWQumx0mR/xOfuFLq9VA6lgc/F4S6fSZGnHi+VAOYUo1Pe9Pol
HE/jB/qEzrOOnXT0hZgKQPyfKtL/xuUm7GgtBVAuQskR/P9vW+oYtnxxs9hMjst9
lYXSpP+PtvoexhLmyCSardINR/uDtP0dJGmTKKQxaBOLzzz//li4wCmBOkx3tVjX
jLIJcDTpt3Lbgl/T5O6fhLKKJlEEPpJkU0HG5cTSIl9hstWiL1l1XfbHFef+K7B1
4XjD49ven2l23Mu/2+1mCs17lhYBOsM8Wi7HQJFNNkiof2UAbivhGHRcvwHr1Fk8
sAoCCOO3UiF2GOVPL1+U8YkEMoUM52H9LrxgugBXFwBnwhO1y+rG+QJMiPOaELNJ
yucBVu7Xfv5nVqiojngQ8KMrmAvn46AoEpbys/pWgTvFcGgoUSXsCvDWVdTyR9y4
BD/5KzXrwWbDe3K5u1sxjbfZ2x5tZRkQuLWvvqrP2d8Zq1iin/bkBES8dr4ZdrGN
OXnfyETPAkwQ517hpGVD+dhDx4LV+0NRbt46lShwQ+6LBYW4dcrcwTFdW6V5dzVe
FY8MCGvpbbEgDtnWXRkNXA2T/kfsNlqPviZt60aBRNPlF4ks+jPLAb1kmRsJDKRd
ANRNxkQCP4E4HzVdBcsoI+Gbl7Z4XvdscLRIBL23l1L7NaI6au48CKUfPe7lFGaS
1ZQGcfJ+Ze8CIW5KhnSxf2wVxx2Jl6LcPFRdgkXBW8D6jLNNOwRPYdSM9XDD5YTT
GO4x+0ZYrR9EeyMBbkM1UmnZE8FXv6m/gIaSzqGg2gb6vBneviofCaaMQBUwwRUJ
lF29lvjMkkud63qGKQp5xkSXFfGy+h3im4HWoOHyGqQNdcua2iJH4rXwb1WvdboE
RiJc73Qecr+YzmYG4r4gWiNsVTYBDEzwnMpz1u01YBR6/gQyg9opBhyzcV+DObow
fhYbvrUFJp9IhGz2tE/hob0ErJqyz3JJY/awjleEjjM9sictDLpXFZ2LpEzyITke
00ug5jn2AzFkvLHPOP8yTBwhPGtxmdaiXPpsPL7LSasynw5XAfzs9DuzdRcsZ70D
CWvAd+EwuppzCrr+WE3zHVWTYim0pHM3PiIaKHUVc5gsRHXWJ2x+UallLUuyUjvS
FDp8dwX2kC4l/d/h63YP2Ae5FGlJtbwM1wts2Pqw75Rnj5F9fYpEYxZuhiga2xeX
BF1bbMcGuag9YSOrYseEXVhhfRAlZ9X+CsjEFz3AshnJl42C0qe5OA924QD6Ahof
VxBCThh0ZlBEMWbZ9IpWJ7bjfYDwh/6+Vd/PQAzkeD+i8TrM37OXRRAvFcvFALV7
PdJBZdes/MhSGRtbxhBx2GIAvjIvq5XP8OAfytguDWubxpCH3+UzVpJMpOC/wOJA
0t4JQO0+tRGGC2fM3jSmATcWXwq0lYCyxVlNsDSMIagw78Xi4CnYGb4rRwl+X3x8
2m1FeAR2FEP3g+b+Lqn+afZOyT26MowKusbDy4fa2U9DsAKbYwjo/JgcpvqxRe85
vA1l+IbOab/B5afU04Irhkxn9LhlSfNHRWillkj4DjY/piHwos8K4YLyJDc7g0Tb
hOqVu72PacencfvnwCQsWexgDfI632+sk84ivKMO6TKxtNbC73o2loXadch6bNmH
1G7Ejh1e+CmlmrF1hjY4rHNk7PN/2bC42WiqK3YwtxRgzRUUVCVfLzvRQvv21CLu
I2fhpDg0T4ZjsShWjm1cxK/IO6ThdzApbcPRd8IIWIvkoMZGW1QVjrztXT29aP5G
VhnpFNIA9uD2KIviRDMLrmDE1ZKWF0jnnJgRlfNvxGFfHTQX6SUkMRCiVv5QzGS/
oG1qw/z8h/U26TssgCt3KPIKBJanNrDtKZJzbfDAqalxFlMAUsf8eZMOVcRBK7Hx
jQn8L+/McQyVA31m13ewmy89jGr4Dg/90BlJiJHawf1vNaaOuZGxoWbY8isX23zq
Z5fYmQXrPROHk+WA/J7r1NB14023LwY4FOFFcmoI9YTzA1zhuuR26cpwVgJ7akUD
MfLxVYAdUdJrZaVB6cODt5wdr6THFSJf5J+Fb8pCvhSqbwvUyQ+xspPEnTf431/H
kQfhnolQ2NHEE4d1S7wQ+wCBFc2bzFMhpsR6dqv3UH5/Y3oFEYeaXXxyXEP8Kykx
TYVcwIRvC4NH/JELTkWUuvcx/VWXCWxJtGzDdlEw+MdnaqkhPzqzOG7bKErcLQx9
nkHKJ3v6EwO9dd4gQY5PicVl7nGZLuN/bswdPJZUqug3Lwent+eT7Q8YLZdVGVr6
yLrCyg/XxoL5u7eFwB2rbiVA2m5f/gXgknSPJKg71yndjuztRqCpTWEQSpG+kOIP
WtzJ6vr73z6VYN3G2e4ObNhogNIyIABeNEyr6zHfXFQm6QbrP0+SQdWwgPzNmlDE
UU3CJuCpHzB8i/SPxmm0WuiuVOGssApw+qvT+Y8P56QTFAdIEFNHXgUKVhzTa0nc
sAkR+tXTLhmQkYmffE6ez+GgVmAvcv2CUJ7jy5+50DKNfd7TJjnSdnsf2MVTIoRt
Zfo/T3THjbed250Hjr8Z5FqStqqaRkgCdWyzoYV0m9v90X32k+LH57U1NrgKJY4R
xog6K1RFY1PszdySAp6pb54sCxI/Q/nN+Z03HLAedSnIARgMoFD59yW2YOS3Blqu
b31o3HpoQu65jn3pEYAOME5EyCwFjYwbRQ8nXfvYqtL9/ydf97BOK/AmTR8DGqVr
p6b4ZEB7XZtQbC2r7xiuD5r5An808lfYb0XZlYofQEaxQ8iezax0l7FE5nR4TQO0
J9Pf697TNXEDwIbFdCOmWpnvUwp9XOUBjeo2XEZDIrwDTxULd8m8W5OKtP4L14wa
05wWHRtzuQJzseyjhlyGZZ7nGUYaepA5aBW4C28zGwsKUTOXUNRN0gjUEJjLl4/y
yx8P2tGwu6P0dx5thNrYq0dfqYvJSIUCgw5vy+/cq0m/i2e6KkFqewoY7YECaLBn
MvXUQrAkvviH1BELlZyBG1I/2rPOa2JmaZ0HVty5j74Vh2CaYjaoylamrnhy8Nfk
zojd0esF3gfvGzLaNgWKWyGOf91NdrNeiPPLEEQ7may3fwi1X7OPHu8vYhuMYpna
dxColtw8q1owKFDH6ldtSBsl7eXacg+kZdttpb6Y7az5827Gpywc9TLWgFOMNLKG
Gz524+H8b+2Kn68Jp/5JwlfBkvfVt/tdMcpLbK+5EXcQFZ81N2WkRKUM1YySmvpr
E3iO2TDCxlcZ0nTBOcLc2nB8NMg5dcdQMvwJKbludenAetipwO6AdKWZK1iVUm89
dzcwcFtPqKnAKv8J67QGePIzJeuHmCsB2RqszuS3/Ie2l+C1qQwTbAXW9yJF171l
7/5wWvQYz8oX/PBYGQ3Iw5+NjllYfBiBTkHFikbICXnShPavor2KPqMXzX3CbpYS
PKTC+6gXGss7ROrPmrJc1iNiHf3J47FUwcw+tQ6hVXcxMRyA/a/Ns76rubJ4WGrG
ltUG8IbbdVJp8elDEpl6O7E4Y1w3u8iHyFmXOAI+Y2roCBLllm3PPtMKYHmlinx/
D+E0JssNwHWFcXKLcN+F6w==
`protect END_PROTECTED
