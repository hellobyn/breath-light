`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pn/cDITUob9Y0f3p95Yc+tkcsjCJHiEo42TdvuK14xAP15GZrvrpxM5OhLYsW3J4
MLYv3O1nHsK+/p1pEj2NOWW7ZFCov4bgoWdOTxkbr1kD6O7uLbzKVO7e3I5ta2Hm
Jx11XhZDvOYSLQQ14VBVxT42F1VfTM/jOckn4t5mUXSS5fIhqn3/tPtGxYJpFb/I
rYXIoOqco39HYQoucyt0jbQ385bnYZXuBszln/BEP15av4lNHP4SmKNlxc1VBBZA
IH3zGKdu8aaGkHY6c3O6lzT10WV9SzRy6w1eqJbup6ToyJ5wqI/Dn60/9ss19WMG
OjHKDFVhLYNU42MtiGL0rM4G5lqKutgy49UDRtSDhsdrJGwpFOt2hUwl7Xnf8oxA
KVxNNeHv479McpWa/jo05pn6RDo/dsOV9Jy9KcjXzl59C4+lzcuQUqcYsZ2raXfz
N46br0yDEfNp21LJwDQUSJeNRFcWa2cn9JcWpj0pXZPFJHDjNUe/toBYUQqATUk/
XlP/ZqBK/qf0xC+ilSbOBvt2Lpk+JyxMHSbci39OMedeJBw0W7Amo9Kq+rLZkyWK
xMS1+WcbMs1mSgGPZX7XnukpVvXnNv4whtNx6U92HvkvgS/dHeaD28K1fUzoetyj
dxLS3XDzicEN25v/bJM/aVw+fag+BAi+iqM/TlWWVAU93WXuvQEvhYYgheyQ3g9C
ngbJ+XpLSSG2qkyCsqgr1JFY/IQzHa7gD6oarbh+4XrlGHBVpZZJ38uh/WkzB8Op
g6xN5nB0aNZC0l1+qvVag0kp1CYoRlwRXQ208ivR63ERh9e319iIUXRzDv8Dzot7
DiiPBsDckfAuVoqg1wQqsv2ZiIX58kfnQc+n198RgrHl46TSRtSidcwFlHeticXq
a7Mhtj/pg88A5KbT7KraU7KfhF7kCvEHXqKXswLm2bDPZGwnybratubfuTQ7gqZ+
7aWZhZpdOydLs1VpZgbMx60ndPSG6Q9GZB9yX4HsV2m39m8HOTVhAQIMVeWPxJes
EuEOaVKkM9llDg9eikULD/uul5ARhuTBshUkTEFSNUHIXYSlmOElZJUqnAurjxi5
iPkmJ/uabrl4WHY40bSgqbQJ9GbrLTfYooh+OtrrRrtz5i3/K1eTyx6qmzR2fq4L
8vPN/aB/Adw3wGDmi/LGrd6lpjXf2LQHcxekcZtiWpIGoqogIwzEnAPgAvwA3HQh
He/pwlnd07dh9y5ss+wB26CYEiZ1w6OnWV8yJhrWYVHUViSsVGuR9T573s8oCiBL
TtzzIM7ILhij2ViRJDpyDqqNKid4pNPgMEiI0MLVBiiuH5RXvd55vMV/o3nyT1NB
x6k0VFlOgJ2gsNVinLQggrSFzlh0SgO1creS/jGkRAq1W+DwwL4ob8ptORmUw607
3n8Cj5dFQbf2i2gVPiJpHV2/zOuhXdrIJvNzCSkiVZDNXstYKXxkWPYbI2BVCD9l
20BD5p2LQogT2rfniqn5V7vkeXg6FnbeaTbJvrggpFKY0GlkfsmLEUuTmLcweul+
MumFFiJB2hoglNK3nLMlMzp2mxr3RxYVwkZfpjOyqsaYOMpV8SVQVuofNUs2OI7L
El89Zm9LgFN8IItVfgwLwKwBczZf/0ckciWB1yv5QNuxz7vUDOHrA+GTM1NU3+AB
onzeqfr01a0+WjTVoV6hdujTJFaj/EnsBZnZOmGwtkbEulqkPkFx8Y2lVRsS1yAz
BICGjT8F5x9vqeHM1GwpLielmXmt1LbDomBHz6W9IIrpuyCvVN975gUu8shnZ2TS
x+E71jDtnY4PZBMYwdqjZw+WIigp6b4tl0pHTcqR6gJzgnJV1CU73OFURx0tmGGp
OL26wGhu8phKscUh8RTa1kZQgBS8WZpCVsxmfViub4IobqoTvvFA1e4QhsVhfZ5i
yWZ1/1L/lwlzxd/tvsK2343JcATHh02SNXCorm69wU+Cd1xZS6JTMcnIvD6zdR9a
IOshRgMyqpEhdSaqf1NJcygi5TpvdjzgIuIgfY7uzQQVJ7QI2QMMJMQdB366x81L
3srWC+BcxGffWTN8MeCPKuo6vYHBqU8GmR1R+XyojNWFg1rWrf0xEBWbTLzioRq4
RznRH2HtRahnLgTvtzXGRy0gi5dAtoCraMkXJX+TetOiXLwjnH0kSWfgxjtnCXCQ
0cLkIlv3Upi/oLHQPlTpwp7n9qqXb3bZbS5jZkJP3Yk2qsHMNb0kUAM4Vd7GahWl
0XNP/Wm9xQbDTo5TCzDHtZ8uKW3Wugi6J6qcVoOp3k9JA5+/wNl2LsO4N7g4UdbL
XJyj0z/WTn2lMX9X+OyymBUYCY2xeRvj+eBaOR6GVdmaxfGntBz3luW/8OvYS6dy
ui93/mGTfJP2518E+8RMYTsyNei0tHzxelfCDjq/xiw7q3K+FySiGDbidiGorMdx
a183vGisOTWo3iYtGJp/UI6qTs+Sy8bCxw5zeK4oaMO3D0WrRvH0I9XZfgpPCsn9
Vu6BLRw7hAUVKWAKTv0MqaB7Db7Fo2+szVcLG2JWShS7ey45v6YxvD9MqFqAOyW/
dyTiO7RFyRWQD9O1B3wdmgItjV4teDpVo/0ArvrEDkfaMiRwYQMyDVDoHKRndOTq
ugQIiXoTgaLdcqw1fAXCHCTj5DiBc12U55jsnZuKzhH0Rhczyja6bBAPSjNuDcr4
JuIv+Qv3sBt35lPOcAjpMfvN8TWJ96ldTMRWWsKD8zoNEBoi3JoUi+o5u6ISKM9T
IOvVj2S9b5XZHdByXjrPTk+llZA6WDAzhwjuVUn6XrfTck0qhvVPswCQxbzOvGvA
wcnxzb/kRLR8p7vbSRQ+c4VA0l7fdMJ9fKSexSyvGP6J5pq1DOVPwGcmzq/OO+jK
UoHq4+XODCotMa/vxmT8INFXfw6XifA84R5bsM0oJ2DH+0xb1oDTU/+IDGW/ylix
xVwIhpqgxjElkgK+NwKUltQOg3qqBYzeu3Fig2MhAjme9j7GJ8yfLJijRJBhO9Jn
hCdS9Honm4yjBKzW/rKSRpr7DYA/iG1XmXRnCnWJpVCDCyE40QrO+0ZQ9ZrTL5ZP
GkB7IEPgupzkzgv2UJMHnV8woJBgm1DfPRDR0ebNaG8mqROfDvYj0QF1zy6UPxHr
isfmp3SHxvmTvbXpYb9uQ2+Se0n4Fu8wJDWcDwWKm2WOcQ+mDeJ2hyNpxRTU/c2D
d1z0sT3g9Qi0ChMdyLllHTXGQNlfrizASc8DDuyAQCPZLsIBneCFt/pmBRpSdLSa
0DakpDc9vIw9Bom/XqsnSw6Rah5ubsetngovb5TgK3ndEUy2WgnQKegtI+ee4YUO
oNKn4VdhluY+RR6qKOLYW8x4/IghT6+qyPi2jw20t92NbGO9JqMkosU6khPRPSmW
FvC3V4//LWsOEmtOwR1CYaPuVz4nSWy5c0tz3B7vvqS8ruuIk8m2jYXYwJb27f+L
qIGA/wgMt8m7/r5y+CuCTGnUaInLuWTU7TEPANgCbsRSg6JvgXrcjQqg+EviJm2M
GbzVvclKlbvMV7TybiUbpYGPz2uRPLyFAfjQ1DdDGMGV053MN3Avog6ezCKp0hXz
Mr2krG/j3KTVuvWTo21XzH/JKPXdU3b6oaEsRFyUL5t7I2KfArjpVGm0s1ueX7l5
RneRSOgYz0lQqteWzC7mwHRwKLEMGrXzKICSuik54TusbCxlbg9y9WjmhvKNjEX1
ydoxB/7EYjuVZxgANkJQayEaFC9CDsVaRHN+cMOONkPLKCaPFzZNTR9k0Hi8oT4R
+E8VLbOFm0jBMHN5Y913Z+Ofr5EmKpvrqLGs88PAQ7U1O++t/s/3foElgqRnrpRk
RMeHQdUqtWWWCFZyQ/nTUp3sEyFgjCUbFseLyL7MDiM1z+CfcJXrvW2TTtvNf2vr
1GhKwlC/6HBCfCt5K3sppZXsEmwzv4Zak+h4ek3iP/0xzgKL5EsADJFDDKohQnFB
sxGfOy2m+jcho121Ne55ZbvmBUkqrq9jOek4zCJLJynwsXqjzOricsH85aX+0zYk
+P6sI1+CtFhsAgnpB9/4XpXUvWuC6Rn+5lvZItX/7qxCXeVLI+cUjQ1kpapsH2Fn
7Nm87/732LHGgyLt5uA1dAdaAg/zk3fGoHnZiVjzMVdzxwXLCYb+514lNOpJ+st6
OQ10IvHsu2G71qbuKvzUgw9Rd/tqsW16A7plcbyrW31K7G0ij1bDYa0cXYNkzgNu
2N+DgvLhNsj8wsq4WbGh9u+UZOCQneHMk8GwVBy4v8HRhqg6e0d6rKUtrm9FCOwi
wMyePMBtC/feBx+OL/1AEudyUotYFrKWx9nEKMd9WxyXIAI3BLWEIZJt217W9MVe
L72o1fTn8u6wA34xM+7WePbXl6Mjo4oEWmbc4Pu0bvPguUnmiejCVHYQGLpQIKqf
pvGnTKXgKPT9tuKAl5mBWHrZWH90eDlnNzVLBwFoGfALCg1Rvqkk0YM55kd2KM1j
qYbWsPJv2RV9hf6p+b83OydUhQh3OaVKhO8hQvTSLB7tc3Vll1/2s/DMN7XmIr0x
XCSUmTluIke0+huIk3Xi5qzQQ2z6PceJ3KHvVDBOWB/D7dNA7oQyb8qPSZKsGYJd
wcg3UY5XygHyHlziRuYJbL7GJY3kw+2iyuFtXw/pUsLcge2qX5DkrDqc/owB97s2
70VEDZ+9sdIxAYAMQylkV5TutIOUj/sOhUcTR46Tj97aP9wrQ574+5vC6OwJx5io
54UG5yhaThOSIFRDKo8EpViKi6vcVwaoorcgUqcjn3NGUHUWyiY6jI8UvB05Le8+
nOzjaepfQMJtdx14r0QkRoXMIWIR43Dil2SyEx92Kiq7YUhq6A28RuezCH/5I45r
pZdBAetc5Io/NFoJvCdsZmKdq8XxA1ZezXkHmmeeUTbf8hRwbDfhZE5Vf5r73796
4LXYdfVfr0ZjSqC8jZIaQQYqGN/d5JC778B+W7eV3xS1RhCIo/2zPLn5JC94Bs0K
nvx4i8+VoQ+vneih23QZfjuwwUXdTQrAsSTpuxhC6/aS9o5P+eFn2FZwySiLUPzE
NI7v+TrG6b5l7nD36D/cJnuLTnsWz0nYZTlku2Kyrik2vYoHXh4qaY+eZ1ZZuB58
gMVnwjNPePddrjrlzXyHTDVziCmuOH84RxMrHxrI+WMW87IFvTSFfoaK1/a2hLs2
E9ZYBl6E1L5SXtEp9R+I4kE4tCFtzNsDqLZMFCgkSLsINNhs+K+fi7bT/BUt/dPS
Qh8vwfBisSIct7FtHx4v34sQrIbg6fvrmEbUHPd+aCN0fwfLqCD4JFUPEf0uWthO
CVVU+JsHf9FdS+JeRGCFW7zTLFdI+6zmmOJ9RuJjZkGwXecjWOPhIIouPNbK7AUk
8TMBpvI9LITSnSgAA4GatT6E2HhaYlhTapEzXN6j99+WHzzVnUlym57gA1g5uwEQ
cpBTQ1Q5KI37Pqo2cFWOGPFvbMF8eI5w7NKf+Qq5tPM4eYwnNIdfh+Arqkj+kemJ
SMgBtZTsPOyPaAh9dEE17dr290XL+Ucdc0vKrx8V3K6o9bqT/8japQZyzuDnQ2/6
pBu4ufpfHmK1H0hTn9WYHyUG/sqXekSlS6YP268K/uqwrPPU38NM/I0/mho/BKmu
AstbdMTJBWP28OmZa5+PwwlP4UfIL6m7SAtRQjmlS79RBLfDmad3v/NaWCwU8IUD
IR5xOFlr+7rwszfV4e4nHn2KTKFneHDNIUaZFOB8i7t78+MctQYuLvr5nPwqVH0l
BNUa7+mC2uGNeLntVemGeSjxQAQ82z0HJ2LAXBTss+u/kPXovW4br7jQbmMej+fF
9SDpu1EgNb2EZZKcCp9odJpMFFLTz+N8yQ9c9jkuKx33Qi4S52P+lDvQbjADjOWs
0kmMK95wyeYsPOongIBp6CghVnJwCPy1CZPwsGO3YnYVB5rNIOi4UjDoJrX3V8zg
tfxpgevzBHsrXocdi55wggZO1JuZVvFYAaoQCB37XJ2CZXGnZXwvniMWQXTXSXar
I32EHPOfij0i9LzJ3QYkle8cye1VvaDzZSAYNFM8oaT/ZFqfNIrS+3LpRy3plFEf
wNEZBvyzXtq0fvfgFTmT1DMvAxLP2iFtu4ngDyvuRz5+NYnekgiQhqM/BWcOzIGI
PuCxSfUvOuYRujZUQlQgK/mzl9ebzxNFdhmXhsqY7qwGa7RZML9RVE4Iecusc8Lj
0L/avSTDBA3P2JtdPlNRd/CEvuFmbzaCBQMnvzBGh98LhC0AA4xSiSqkaywWkuql
2X7A9Gn7vNGyv2mYk7Baqt1LhI187fEYdnz4SjlDAV5TUqAjEemYHpaIuarJe5AZ
V1sAHbTanvZwQdJAFhCgxTb3WHVLNn3Ei0tkG8qDuySojVmG6vyNpMah4VrTeL9W
AoRSYT+vRpffo/kOV4B+UHQ+1t8Rdoxx1wYxHi4Sy7q6iQMqJHa2Iz27HqKxThC/
23kmEVbqJgCFY8IofLVFbxMvSKwxzvPzN85VU2o7PFhrbRPNdPoXCPcuOanAGVJn
0D3hcvuPpLp7blsaBubmSDlQFjtN4V66RuoCgCPe0L9w22j57W17+50I3zT2+LKg
SJuxsiD16yMn2GmcLxvZhdEemtSEN6JRhm6iHsL63dCpdzZC55bmqnnlR4i7/4pb
B9mTI4tJcdiPaS8MzhhlaY1vAxbKYJahox28LaTls/MEsyTcY8pGNk7U6c3w4BAh
Hpo+dLOfeyUI68TMiSGrxkpsDzp+G6eHEiugzavd+/BC4FXkfb8LB4ulCa+XTsTE
al7oYm3vQTj1hFRUG1SGjFpZBXgkrJzZge7mUqkasXcKQI+e5cQL7SeM6WfLIiLf
VjNbqt8ie85n6HL1C6o2ZYkQ84Tc8R45QLGY6AqGgOuLBLn3/2ThtQJVpw249wX9
9WIvDZ/vgeg7tTFVjtRXtSX5/OcSZRjeij/4zURNBnSM/koNcBb0CxTXkhmjX3Iq
idgqUnXkBD+LHc2FI39dX/P+61w+/w2GfuKYOCgbmsulkZnarkCf2fr0Gb9yblvV
EJ4/fG1ztqacXIvq/TibIq97ahzSI3M3gopCD0AztXo4IVuuHyXnBOnJ0l+MuPUf
bTJ3aLnm8Zl0pTKWmKXhpgOpE5Ai9mUhIdNn5h5o0Wd/S22gRE46WpQD61wl9Xm1
UpdPhne9sUqztqNWBsfN9Omf20Bc3TSTyueLSOf1PdviV/lyt3jVgmIDev6RCjQo
ZI3OyplHN6BqgJ7BKC7YKUxsDw8ZMUzh9X5xJonytJoh41P+PzP/5pA6T+4CTMos
KSvdSPclC4d5+OP1VPP4IEA9YJ48bG0sUx0zol5WuFApvSAULnonqGlHw1ZDCECm
7km6U/NrYm46XPWM3PxPak8xBe/UWnY+MSV4NhmEZS3O18Ay4MkMJwxZI62clH0S
Q3W/HdQtEFQl5OPAiig/fSAYPWu+a1ejjLZWYy3PNM60bNXyQqzJxLXzIKkUu/u2
soU922c1qrfGy+bTItOZ1ebl28qTf5TMLI3fFA5hIrpV+X39RybREO0CHCmYJ6Nj
lwjZIVhD9wwACvGMTIRQColeVup42RfpBl2RozJs02h35bqPLRBn6XrCTsyF23QG
iMdkJ1nI/pso76T2i4TqsqSeAVZFlJOOgDDzZApwjnmxNGDvvZsnD8jIvt1USkBT
5DI6cQjeJoHEzchcEvS+XCAYRybYKzNOwCDwmSC4YFTxkODZv/P4Z5xp2Perw7MS
PA41xaAL3zTU7/HRilvxfBLTbskdnkDVQaCcDU4oOvlfLSe+HRmW5hKRcOBMhBz+
kNuAPXb142ayQOtiaJLTNsXMLRO4UKBZ/auLvd7ArN5SOvm3eZ3s+4dJD7KPa+Kg
7V37rTE2/pevtkL34IzgbITrD+ouJEVmttWKuSPqQWmS1ZvL9WvTWcL/ynTSzXpX
sQcCTwlGvHkOCC1rhEh9pAykM8sazp/8c8dnKg7JvekR468LXbPdKvj5+N03uCq/
IqLhvkJLhE/CzxPScdR1RE3BLEBPONH1nLrrUf72pGoml1OWbpRGL6ibIoaKsYo5
dB7zBjM9A/Pi6BMEDKO3JXPvPxNAgoW7cZ/v9naLSYsMgup7xMzMOnuDxuvz0dDo
s2HCs8bTifkhHNS2s/4Wrwg1IKJD9D2nHbWA7VTT8XTkksE5oilqQ6YvaVR72Qxz
Bvm9Ajs3E4fzdHIxEvXqqFaOj8Pjk9+ltJf7JtGnYENkSer68JN2Sid0r3n5DkjM
8s1J3/H50BbLNArSO0ee6ufsLbXL3VEQnGrF420IrZsUfT1/rlc3X8UqWoFD9LSH
JaI5xl46y7C9C7oz6b0dUwXlG1RaDxIKgrdoSpwhN7tINQ+mjFURLC6V0b0e1gfN
6TC9xLDTs+z7b/T07N+iCJAmkZiBC0dPpgsxjJvvuawAH8lnulC2gxjytf/soIGD
CNirBNgwAwh96xU/thSnGWDs/lGh9neCjN/8kA3IGZn51/ijBtIbLXoDSVc/0/rl
veMVH+POrVpoyVeOeUQvLuiWbswaItNd5mjGEyV9qxixIaYnC3OwqeIyK1zMWHll
IXHe6GsDRizGsWw2SJffvk5bpYukMKNmwyJHAu+OnGgislIS8v7DDUpCETXk9CBq
UDI3JTmP64RJJ4NakDfWu2QUWsdFt+fp8/ImrLRww0jQLM5FgX3KIerBSJMBbRa9
jEHlD7CH7a2YcqQjjYbBDEtzXnGH6c9wsGSlLi42Grb9MvMwgZw1VmwXzD5Kk9zg
thX9k1N/6wHixs2HY273SBl7k4aWQJoVtZb9CiQLF35yRFVeo35OjPLw5BGpCQ0o
HzGebWXX4bQgnliu1IhkmtKRQT+RZqhJ0VuW1S/PS2EaLrG4q5VAxAqO7f0xHjet
STggvBqcMYGqBpVzCHgZBsH2V+ruphr4oPjw9HfnBxplMQJ0p8bcRt6T0haur+xG
3t9PQAIu7Ac9aApFCzNO4aDUxqhVynK+RyMZeNR8cQsRGzgo5jPzAmLJn9hrcXbo
wb2ztV2rvfZvHyAneQgZ4Cc/rWVamJbyYZpWvd8NLBOk/RTgdPVCRiAmeZAWLl/E
UShixaac4aoEkbeqh+dmG+Xjz740o2w52FxQkcljqjMM7AGzzLnrOZ9Wce3uKefC
qxDT2x+3XQVR9W7lvRoihVS3STT070a/xRuizlB2YzkK5YnhPWU/NHQ8M9KulOQk
pOLSQtHufggt1JpfuocKA7/3KHayk03J+7+v3ajqTRb8nJlGBWgfmpkIo3JG/Xum
rDtK6BUqaDUIq0f0kyeuirviBUqTKTKg6TmpEHG3xNIvwwVQw+TngW+szWvrlUW4
cVRzD4ocW7UplXgubykmOb95PLOzXSQLjafZfgg4EXt0yXOFOz1Ab6aNFs6PpiYo
fzoagAUeTOYQA7hOSfYOnvBhoGXWfOOGYEFDngLY7xlPExKrD5W4KEc7uKD2JBve
xQ1IWL3E/cLV8I9xggcYHv9bkb6/kXYl9NgUqojyz5x4k6COYMEj1BuEDpBLr1wD
WgHUX8HNec1SYPZc1ESwULn7o07nKw3C4QGEd6S5ynrJWKC19F12lEvfdTJIX5Fa
F3v5yhkXN9QNRK5U8wPbVFRY7sYmetCCxYDaOpWIZT4cI2jYSHH/J60meZzN9eO9
kwHvECzhpM8jhG2U1FHykKYjdEKVeo7Zkqj/yCmWNWDg5o2Yq144t50YOQDvPSq+
ffbiHq3QzvCTHFZW8a8clwspdVDrso4JKMrhTCmwwS56kQx02WUWHGsjV3paNggK
nbjiKLqRQzQY0XWR5jBnafcVDQaS/xONu5XjtkeiEY0QrAm42eNbcEJf8kP3K7Fj
Hn5doq3YgljzVUCy86TTF5PkPC/eFEkssFAKFrelbEHmau0VIxy2ZXM5xDvXtqN6
v6JWE5sBUlLvWHGHaAynOJqPlOjxaQ/yRLShoTXuJAuglZsyQ7ciKzojaI2AURmS
acnJJDFpVvtmkNhkIYnYFNzIFnDsYrqAJa5G95xTCu0pRgTxk3raVQ6TkED11bbP
1Tq7shEWdafRy8h6xdbc3P1MJl3Q296bCrD03lqT8Fiikv9ruC3b9oWw4i+j0xP3
CUZt4f3LXsO3dt5W7LOtWecp9yG6dR72lBjdR6sl0mxrY3GFslyQ6qHYhQERmdPO
3ILdUwcHwVNCIjP90rBbCc7kYFmfRZiLtRAqJSnHlIROJ8yKhwYruPSGkrn925Ig
MT+g6Arc+q2/03Nalr4mQ/7ADiTU0S+71hAEeDDrbp45uwTywmXXgb9LHRTiBDF/
P9cUjx26nntSf0RbGKujsHs4YKarjkVtYIHSzT3Ltfz98ItxdqjDIC5JwOhf7JBA
Tgg+yIbUtjARAMtvYvLUKqh0bhEyFU65w0nQCaji2r0Rkt9D2Ck7idEPlAKdj1uF
24ksb49P4+obWsGbF5Kzpga8j0aKGn88xLtC9eXbBjXpummoMLXQ9NLFYIXSJH0R
LbyUGy4MDkz0BD32xQDa5qtdPtkKSKFfhPfR3NH+i4S4KA8uMvX2k3QXJYVnHBTT
w59TGHlWhwAe6KkS4WzWk99OFDz8YSEC3Rwa8b0OgmM/oRoUOHaERb3VoDQm5LUk
j460i3d78ukKQ4e5IjISHU1tQcNE470r0f1CJwZ4J2IksGfknpid9ejKw15i0pSP
HcqvWrW+dUX0ju/SNaNF9udk79vJKaAm9tVJJVIiFDW8STxiI/yvZ4Htr3zmyT7v
spOu44GBfM/nQgOLUAbvFuPA9L8kBtw1af1hiuvy3RThwuuOPWYz/ckTzLrfiueW
4lJpsNwPw2dbXjJ8c3RZhmF/S1IqV0z3O2V/0V1Za7mHki8uhIx+CxJNDRZDaVDz
PsInmzxup2x1ULDULhYQ3Wwqfa9tstW6Z63hU8muDVKMAtehtzq/33llIEkrRBzc
oDm+SwMW7jW0bSOhpE9k9z+Yg9MjJlw37OuNi13sHw1PwIidm1mURMX8H1YcMn9d
MbMb73XFvBfIj70z2PD/XFYxfmHNAxBaXMQDFC909CM0qSm1oCdjA2HDcsfiHM9e
ojj1IRcBBds6VuOZxoBb52FPn2cX5sKmrpCVFu36CknpxKMvFsZrQ0mKJYbDsD/6
Oc0czQuXbb1VCLnjTX+/n5Kqetcfe2Li5NwoeiqoaDblpesTDRJ4KaBZ9heMtQii
/V1m3SR20RWHi+ZUziikLPXTR4stjYQ9B8xKhwHPcoC8UsS64S70r33thoieprnD
JBLXcVUxd6vDcpX+vBTJF8LGAFUCP1+RRhcMVxQXHrlC/qdgi73DavD6rxF2bJr9
WJcgUorhrAhBMDG7Rf7c2k+aNvhevxa4q6E9Vk8qp+oXO5J+DihlEjVr1H5VhV4u
zx8jUcwfWDcuI6LLB0kaQ2I7qOteaC90BPt1uqbqUDw+QBfU1mfX7DhVA29ZCEV0
E9QNkvqCAYu7y7C3mOTJRON3smtQxm7X6nPusVZOAWsM4cKQtAGEs2Nc1q/2cMX5
B1SD3+AYSucvQiWwAVN1/7aGUrdx1f/SXMES1Q4szdPY3a83VQS7E/nFQwOpacLo
zPhOUig/FNgwjAjbaNxfR10OfPM74rfe4XOxH3D0Q7/6XDOOd1i4xj/0XAdf5iD6
RGBq1v1pqpDmpyV81hIscNo6HrMZC1pnonA4iytMfk2w4zRJN7Xz27N/xZkXUpij
hPQyYTVP68LWK5oCnO5MNhfQ2h2/J340paHB8poGauwAFDwbvHTG3IayDh9ieSun
FOA93Ty1Ia5odJUa6Tiq9qlCMDDyg6IfvuIcyT2EsgeuTAyI18keRoOmQjkYzPwY
IA/VbNuUjQiPwS9ESu4mqfv4TMI89eL8hTGqgqt2FwQouKTZCgm6L2ztVTW5mog3
hsvtYWgEVzSpKtPzsY13H9jvOf/A6OGU4C8lGeCRg4fxmyxNBjFBTWMPQg6rOEfg
wH96H56ZXNaT8KF/Z4wWAytOzRIOiMrQJYAdDct4MEbKgDIg1raLCmz83pRTOZ1D
PRaf6iDAWbmIBSN10LbpPGd0WksWt4k07ixEy85Nnh6BOV7ZeGBX3c0+WBHoe7mS
UXxeLKYacqXOgnc86EfwoKxiGokMxUvOG2OL81nG2N+0iMymqgwuhr0NAA/sSfT7
TD01JiZMufxO9zjlwNFjYb3b/foAbjQlhMUc1mWWZ6fkNV9MJImg9MYo6jgBeOUw
eHp3eDBoSS5RfraBGKZdhOSahLQ7X4chBAvp7qS1k9E7h8hjtm11IVecBr5TD/JW
rDxOX6v1UwQ/zez4sUBZdvxhhye2JpGCbOFy9Pw7NRfyjU3zEBh8D5Vc72xau7ZQ
gn5XQ5p50N+0IUoC/CKkSNhdHmw6mQupqm/clN3kQ9m32+XJAVMiLKDzH+wzm5xn
Wf8+RBHXF4zD/av1iIA57DZ3p1EZpAoUBE4aH/2OkamwGzy3y7FJvOAel3hjK9W3
8AaGoohEWb0hhpOu7BeqOccotz1ZreLgWsVXhEQrohYTS18iPyd8VS3udEwUlns5
5wg5TQF5+HHJntfOzrBf4cNuVZTUylhG/wZE6ORD9go2T053QOCHzzKNRcQM6evl
WqDYOab9WYJeu2V/063V/6ogylI8Tr8P00r/aNGIL2sdsFRxGqMDHHjrw5ny7ADD
rxWfdKfACFA/mbXY42gIWF39epBgW+4ryfJWztSIYch7G+uf05dAycXQyq1JfW4a
uzs5trP3CzC9eSeVLiKjCMqLRIYNApvKxQo6HzYIgXkHVvlnbQr5atN3ws4mn3kr
PwT/V8Ghj8jfu6uZESIXpapKEtHdvXSzIdBm2ZwQcDhguV8IfOnqZYLj43yQLkuH
TtSZb/2s/Vx5zjrZGJIimrKXTk2npz+hATsIzJHvrUU4nq2+tcOo7QBB5Llkmy5o
+iIuBnka+mxBaV0GSN9zffSl9ir7b9BKu2ILhcCO4QlBm6h9iSLMaSPdFKfFwge/
sIKuTayYRmeVtTqZ+vMSOnKbfxIOwX8/k/zkUlK5PZaPxajaVC6hHSV+JJdMRQEx
ijlOOS98RNVOxgkuBs1K89oWvwrD9otehZra5qQD7p55iukROI5lwrCSxbZVayf+
Uf+cQQ09VqHDz7sApGRhHKqLKKm59roX5IP6DdmyDn19rDzwZ8lHyE9xZKwszhpA
jGdyqjGpoz8oPFT+oxdCpHSAZddjeRk1ScPV/NxH1KpaqDcUDQWSgMCdjHmhf6Ui
4QlRgrJbguoRYz9ku8+h+4GR4xRZAoWVcUrz/NfJI9Y7jF+/B/vzAQ9fearvpeHZ
J5T/oIsjiF3GCPmIN+0ixEiBakfksC4YMHQZCGcbTL449rPwj12uigdxUMMLo3sx
Q5AIf26+DDjfifPhOt3pOhLko4g4DwDS87pHG3CZCrxajDWVfuiyy1dmGaZjKjSy
SFPcbD4I/HOVJx7ht5NYvEedQF36cqaCDa7FPg7nTG6cwzPp25rAPi1I97w0RerB
LaMLsev6gDedGpKUYuLkeAwHeijhW6vQ6fz2DCeRiXKnAfciVxLlQ/83cDXQVsJP
bTx/zydUlcFaq+EeFHo8YvxotmTBB+nZWseXXTKOwu1riUcTKnIYokDs1K2y0KW8
0mZa3cS7d/Ef8EM9Y03jVtEf7EaK3igs7/0utcNzevK/eOw2kNPr60RjgI+BRKUJ
WPd4mlkZeKCnfQJwmr7pcbmQRTUu5NgX5BX5U5gTNUell56OjPm6QX8e72GeNfYS
17fYp9zCUxDJnqN2P7c9BuLViZiU/hbARLlLfijdfHGMWVI3z7NGWsyXXxJPxt1d
0uzH4B8LQQPvcet/hnJSCT0zjr4Fsmpg+Gvi4sr+PIO/86Qmq8agHucPqjwKBHre
9+CStjgCMpNiFZ76zvy1wKbY2y776npM2IIX4lCHor1IWgOM3vVzKKvWcWVWZ5zW
CIARZrn/D3hXKHQ2wsQQ6eO5A+x7s7HgaJYz/x6H08axkPdnBF1V7i1F4Pxl4etP
GsULPgGPC3C8MHa0+G4bCBtMsAhvDSI3dpwABVfypbwiISOTbHskdPPUsHdKRPCW
HjjF4d+K9+duILm2rnbZLiYYESh0gCbJ/znqT3w1poZPg0pAlrcdVLIPPyHzffC0
Q6VpHx9oQFtNFXfhBpiD3Il0vRDmghfG9eJ/s4Zk9wGCESTjBWzoJMNNNfHIERnC
m5roatCOzyUL9YzAlUEKQRCYRg1Y8DpK9elNxUPYGdvn3BX2okhqTDdioMgueqIo
3nhwOyEiaqzrh8LmhZO2AtRAIxl0hePb6DBqB5Mo0mWGWitmgwwDBYpAlJDuKJn3
BcFwaBToIqHJQcRehXZUjcaSE769G0LRzWI505/Na4+xC5i3LsBLWAfrW9M9gZf0
jB6tJYMMGEvccnDsVbO6h3Qx0kE02f4FQ602xkUjatvO068mCJ0qZf3b25GgIulE
VljDFtr2JJDiMgDKWF8Tl4mBEZ4Fn7Xd4g2wZr2skqBrGQ423mchBorH8LTofbwK
GHANcVsY3NRzos9nVtwN8Vm/bTXiDbmR05YGMeBaoveVjM6P2rzCwhkYOUp4QU93
wU9TSFT2gARKb3UydBKcngpxiK7bVkGkV2KFjpYxdRCUQQsiamhmbK9mJzSWithA
xbhX8EJlHN7zYCvG1LJdEU4UWkFrYZDaLQny5EHts5duKzcwrtMEkZTpgkw0BN+c
4eDzV5XraEjV42USbzqa713rOusya3A3u6LCMLPwSFepmW8A9OqsImMogqnUrdMw
nHy1+qO/JkCm86QXTae2EyLdlSr0ekowF2xDLAz0RqoYexnc3V17fbUi5/I7ZP3d
V8UKHMi9CasodNr+wA/SVwIQvEosrqG6fBoPKi1QmA3iIEpWzsQ0/eQpxSrRRZcp
YKDQKB9vhG86TYs1g/UkApTj9i9N9fa5A/6nOOPExhb2h1uVqUQ7jExn8A7sq+R+
PZ9bRIPLkm6y9nlzlf+Yz/MT47t3EV5Wjva2PfueoPTFLXEWoBFNfawcAnPTwRyd
6DXYyBnwfRucgTmZtTuON/MBCYE97/J1xxx1xRViMKWUMLfaLb7SXYG+IXV0eTKU
EmG5HS0/QpkvrLAuFJFxTNd86vhJsTujoUZntQofz56BMqy+KTqJu0vB5MSVd9QI
xmwWVSDG0eNGMc5Txn4AqB42iA55g77msXmWOywk5yB7ZiqeF4UZht+Q913PkDul
vopoS0xCMjGRxVt4XwQ1q+KhlNHy8kg13C+8IauQA1RR+Q/lIVtPBQlWwhfktCqw
ioAMFmcCcQHJxj0mL+5dMbmZ+SeFznQaM8Gzv9jjcxXeV5fTjsH2CpAnAzw/IucM
3CC+67GbH5EtrOcFXlLGxNM9TBP12t8lvo7roovYsKTOHG1yNHHJCEdQwO3MsRYc
HRqg0Q24W/ZgbKR36ST/aQ==
`protect END_PROTECTED
