`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEHsbUvqVP9sUhTAsjN/BhbneapRbpF6pXV3G8piMioFqILtir11znkKD4CZiuB3
23mjBUKehiLFLEWCxi4fls54DqKoZibsgKLn5YfBPKz3t41B4cMM1kyVoFnOcFKH
1f29BAQt1voM/9ifO3kUdbcFXYMZ0d6E9ltw1aHZc1Tzz19TKKJsduRbb1DGoQBm
uV8dPNIV3w0a0m0tItxk7CFRcaOuajmIFzytmTYo4sQo9yQparHMOOXhh7IvJS6G
DIlIzkC41vO1l43atvjT0gjupd+13spzJefsXRPQKpjc9x1ghviiWxhEVJv87IUV
tgxk8DLf8ro+TP2B45yZzQc0UcDPCVPSLzD2NWikh5fgZxA1Th8eIAGE2C7vp4/k
uiuwM1I+zMM0CpeO/vAFLJGctcPqrd+0mbDykBgOIPwmESBh75g75uKDUXt+Pt1e
GepeE/EK4Bo3z85vK10ME2Et5X2uIWQwvlTUndeDdOecQ3X0lRmaud/EMgPTHCDc
pzx8VmVFCk3doU51UX7jiujtt2QPEuRy0ubzmqjB+iAmwsqpUKH55R5CRK49LV+0
6Isblvq5ZWqxRlBFIGHMCUo8Zesu5cGqQ8xn1EZ6qwtZvGJ1w64leuJ8jmMjwQCL
TMVp/qqmaIZvoTIHfFvfjf11AaaS3QZqeiHTgfiyrP8snYkFhR0dsd7FmpmR9+ln
`protect END_PROTECTED
