`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQS6Xn1NTqeop9U3Gg5aZjDmQjTQ2JxbBNlj3Tx1sQWRrziEEk48krHGrO/BniZx
tIjY606GPgsWhUNTLpL1SCA+PUbJGDCoIxdEgso5t8+pGWkWCQ07oUpSB+r3To7y
WnrHFaff3gflOSTJNtKguIMLawbmkihQp0Rf5Q22HCyOe29oppj9+3twxARib7lr
UQzMSY0MYAiuRwEB+VmfsgXI6cZicDGaaoV5lEtlK6wBIZQ0C8wE7PRuC6mUbb7e
GIo/hAErrnAhq/0kuRVQzHZg95gXf2JHvuTPRboM/SCuT0wr2teEEfLcOcIATMwq
d9w5oLEG6BlRIeDLyDHuQH30kR005OBggyc9Q7KeaxELHJVu6UmMJqrPn4csprsD
E0dlQrSu9CsY4vaIvshXb8MhDSfpeRZTvYn4ZGNICDtIZZwD4jgrpSX1kbIdYfSF
9BgGgXAp9+edq54GjExU96WbcrXKPWXvJMpheIhb2agPvwbT86Y0skoEQMcXXIXB
y7F3zs0v6A+ShXSycDv3YmzuWZ0DQmEmzVI4gzXloow=
`protect END_PROTECTED
