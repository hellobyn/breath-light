`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nL6cMIeWrUQAl6AjbaEHFQEwz+bIrA7CY+wyQEIBDpvCFYAYr6WrxC9iF3tq2lIR
e5LquoF7RcOOpQEVg40APEcf/BAT9B3ySUZ8wk1mHH5bOzfM0YbdGD//yoCzgr+Q
uqYO4ofQrGg3A4z99zR4196ARiTLk/nq8Keg/1OVeiA/CS6OXArzd9GNr5yLDguH
zx5bbWMLmfYbWP3IK9jnom1vbU18Op/RMBnBZUHm0m09kY/QRobvPzMR4o2R/uz+
UXFfi3e9LV0WtZpcqlrvCTt/RDYedVQfuNuCXBSCKe2245Qy35CBT9kezXusc7PX
Lst+IYzKAQ7/S4AgxNBU3DawXiQ9hA3ppnKWy2PqH3MH7J29IbkcsuYnhdZxUZ2P
cVnRU77OBYA6XGsd2XVRCKoPy0OtXRlqIx101P27qns7pc6znQVwj/REwTPKpd3U
6UG6BytkS3BsS9cn11TcBd6+/yXqkN/cUKTyT3lZqtqVmu4sKYkMoF67YafhA9if
7YaDwzDhEEKj83OICFtXHq7yLWkqsiiurK+evDiFEPEj/whKCKlkIE8EoLuAwA5P
tm89fGsvkqKeMkHAihU7U6M8C0snCQ38tVMBCXyhtkq8UQ7DeWdUCysB8qYqmRB6
qXiNCHX9mdGG/rGh8pcuCs33FX76Lja2apPyoDGBxspBrNaeCJTP/1/FN9zFbbc8
JJZ/JDMqenWzQOmLZK8perzhPn475MoOK1emd7+zc+xna/fLR2lAvOI8tkj6QBS4
jl2DO6HnDgA8BSnYXpN9lfKdX8Hgc0vnAggum48Zxf1+cxNk7ypz82SOhcYhbeXy
fEvoqpx0fpddghi5frpdpdtkNc82sCUar6p2gpLvY5bVaDAvt3yVI3jY34XbxCCU
m4kiapu4uvT56rOs+HDcUhP/u73R4HyDSFDeg+Gw1TDf0q79uC4kHi4LmZqaaUfU
`protect END_PROTECTED
