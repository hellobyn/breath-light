`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2e7eqA8njv71ase8xP9Tb9d/wbrCJS48Jbbzvs+hyAoUl449AQ7sqyH1iaZEVKy
E+QbzJ4q1aMGNRdF2io1YXhg6otB6UnCYuA1q/exanglUoPbmtIfa2ZKCvgwMtX4
Gn9vZsT2eyxJzwc/pK+Xsd+u+f38ClxEcDP2J+nOZo7AVsVKxxieaFhYs6ypq42F
QfJgWQ54LpV363crH39RE5kXZ20Ukf87R/fPEsJCOIPQmHddzzeYtWCo4aBr5nWp
vW34qLebRsMyYurDU7295MBoafdoA0LpKwJ4VBJlri9KulgOgkmT6EGU++V2xdqm
7LfCD8AW0vCNPacUDty9Q6q3ljde33Cl2hptQJI9pfz6g458UJNetgD2K35xQsmX
DjTQuQidjMmTe9l6zclbdybqKAI7W1/kTAu+g/CLP4YkgsvYEQYrWGOr3OKfcmy4
VVJwWfK9Gm3senvR40MN6+lCt98kphDbdm/QDdlIlMNHksSxq2dnbV40WfvaYjry
`protect END_PROTECTED
