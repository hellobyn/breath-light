`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWOX2lKSeVmg/QuAOWNIWcFNFxe+1AgMUEWXMfXqGJawQENEAkcYGrLKMA79VG3P
/NcrLiCc5kOMQrnaMk5ohs77H0MDVk9n+RxPMry4Tq4ooR3LBFdyjRUiQatCnIRn
DUaCmFAAUw+y63uHW/12f7ZwbnzeTpOFYZzqG5qgvMO3ADrQrdq8KFPH7pisUrZd
oynpa+E9Atrm35RYfImxjAkFdht2kTe2UaLKJrtED6tEX/4U6Go9ZxBB0jxPo+TI
N//Z5KxS9RR6nBWHukhlybekDxeT+32hQn8wqIxeBlDfDndGO0EmdEgPSwsyQn46
39eE/nOghAPgavf7L1l7C0oBXSE68RKTjtgAUnUfUnB8jZ8nIJu5Sz+31z8u5Evb
DuOk/wsz3agw6R4cIz5owqdsb6tTFV+hl14rPomPbVYykPzUEHIRLlQ9D8JKM5gB
XpIPd/4J7R5vKf1wCNguwcuuP5X4AstelVTjlXYNDYU5rN4ha8TfrVCAqo6htjTr
gYm9kkubROq/7xz8lS2w6T0dySt34G7FlPwGIX9FiT74tc2TTGMb2NUD/IKwRCaU
egM7hWpWULAoHiie3rna3keLF9gclR0rL6SKC9Sv/M3SXc8AyeHVtOLa68IKWgpH
pxkIhRTSOHWCbscZhQexjMuXjrQ0xFH7/XKG85ULjVbLfcMcolTXdxWL98fWeDGi
Ns5zwXUV8BqV73Pl04toCJ8t402UV0DYVTXqn2kRlnCdKDbBzdv5EyG854YIqAk9
ZYOTTBgLntgDspxpzAEitvV7ljJewbMTw5fuAdDF54xYAtoiRGtXTE49ME5izjyB
HQP4vi9Pl1dy1S/HYTrxuU3WA+h55/SgsywMHQhH9cuxOUdku+kuRHiVgGOo8a5I
QCqSHiL1x9Vu3PDOMPkNv/AwCpi8zx0fVOShXc2gVbI2dMwRksEtrDodIZmQKsuq
YAbAsOTD3IJCV/ZwlHN3fTsN6UzZ/ifKIrxBVe2uhLg1ZRbOOjeU+xKyxJt5MiGZ
ACeayvEx4ODCKti5XdiOmafSgk7hPmMzFxWqiTtG0PQWlTDf2wTGBnGG9liB1Zb7
bKc6gMxI9Ke7xJdydEod55YtSoVRJ4xwG1CxQtSmKPjtlhDlw5o3etsNcN6img35
XyWBS59kjK5eclJbAZHMsD3Sul2QpU6MlRUFK24yTbxoxXlmUn5WB3UcIqxxbdgT
Jm8OPjh3r8PMu+M1z5EGwcsA4qgLgyWUe1o2i9Ja/q75thG2FmFwVVcT81cX3HC5
2Nqou9UifT8NGIaqSIWCu5qBrh7mH2vYr9AMJnxtz1DlVt0vQKlAdC1tTWlqJwON
LbEJI43mgFYp36LYA7yrQYv3hMwNlWvdZF3ARRAKEJ6N6y27+rZ2dt8VOSu0vJdb
yJdbx7Qq8MQvFXIGKeBCvpTNqpvg0yIuavONaEArBym5kIjJgUp5A/s7CRx6pOR2
z3NPAa2zcdybbL/34eL8IPwlXYw3c/IdRG9s3i0h/WwUk3Qy4yG5FbqMiFPaeBje
/MrsZqp3embCDg9bzB39W6JqLm1M0IIzlcMX8QcG2RDdZIY5drrTo2O3IK3CFsif
9RQ8MusiJ58bY2k33tknIQrAgUtBgLPNlNfKOmBtpcd5VB1+ynI/HjTzcXbMKPCx
FStK5DtkEzCqdng5jI5V3nfULT3fcshAUtH9Nxo5k/riuFAJo16F/JLv5tn/IB+Z
ZqhsIzmKkD9TugP5fjS33GOmTSVWMX4jf+EU9xLvG5boGtwA6Qlb3MTSTn/Opk4t
Yu4GsGiWZxFIzTBXpKo5TW+7I7B6DPGyfS8hXHEW3nsqrZKjMhL6zKcnLbTCXzx9
vVkudPq+WSRkKIftQ1P5W26ad5ouhG4vfmEC7JuurzR3GEPxv64V8r4Y0FT9xZDo
AkGo9i19sBr8l/uP525O5OVGE9P83McN/BErK3trhCQ=
`protect END_PROTECTED
