`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCTvdSv1rp/Qh52v8kMFcwmNKQ+dYjx38kFhboV8s2R2SgAcxAg6ZpVmMfahRrPz
NxLkp4opdD5lkG9gcx3eTwmlxsWyP8ubFb+V15UeMDcPnwqC5RI54MXaJJlKupWt
M1pjRWOhc/+xo4n5L+u0J9WKd2TuCWYt+4h44gkkjNuToD0VzGbc7U/NJElpxvJt
FyfH63UGO33K6/PZDdVSOXjhJkiXWnRFFbhuokBPDkhrHBY3kSVGveQCeYVMIQlx
CD8BVPtB6kQgcJVDzN4rPqO3/8u1IdqumPosStma/bNpEXFPNMjyRqKxBM9XNHUE
1TCBqzLnQowO5lKBbLJXaR1araCj6Z/Qrg+ea6om3GN1yuGVW1fyGh3sNLmi1RyR
34ZpbN65WNw6oURlYsaAktZ91WUX8M/kwcUJbu9J2/Db8GlQZI2/U98i+PTc2+jg
Umi/17+qCvPIaUg+PauLQm7ZG8RyEx5+NoAhsUWvs87VAfoc22GGRdxth8WGDSUL
HF3Pe5D/dhHj1fg8Y04gzUu6q/qWvtIh/zhwgDg4IOJmyjJETNhrvMtYtBnpBopy
CJlxQmoWgB72yE0EwlSSOZk4cHPzzGhyX7VbZTMfb6GxHki5MAMuky+hlZKDybuF
zXr4KjshNNg9DMesUWyDD9cQZG7nMm1+vjAbnT1nWT08aUEuYfrct5fPV6F+TyaJ
ves/7JXWjqT5zIiXHlpGWCcncdmLAws7UHMh9a0ZRqsqmaWV+Z5dQbIqD1OM6s2J
tYNTYgAISfj2NIvRz2RTMS2aT8exeKytbdgbmPhmF5BHFy3MOx8SUnvCYViakeTv
Etvnt6YjxY60hVMkEZOFSKPzh0ykw4R47/exBLtO4htVpTIesQZkIx4f3fqSkUUu
DY2DCMmr1jJPFZuBSFbIWwu9YIb411be3OJRQiko1zEbKXVYG5AO89qLNoJWYjMh
WlgPTIjm+au7EaVQuihiccoPiHZDqbGhdqp3XzWhdpX8J5H5jG8l08WG1AEkyAjk
vCrm+xp8N6WyrUXrf9d4aQM+jNI9ZAUSwcMzKR6VG8J6f2Ym/H5zLIVsvTQIK5nX
6GHw+9SlA1Tipxn5aHflZKQSPCFLddxR2vY/rXLK5/jZbOtRnFkxPA4EPkLyKPCU
lhlEq3OpxR3zh6KfewBpiu93Tnh6JpQZrOucKDnvkMoxeHmul2OBSMHeAUytPDWD
5F8n4B6yLe0RUfpWiGbfqWVotmSqV3uCNgQ7PTV3ChWrh3UfFlw2DBKuKaIpPpfX
rZEM0zCzjzTQ7w6anR/eG3ADc++1w5+3usyB7QPB4fjJFB6/84XuGCo4R13gRBxu
+62VuynfKrZQfiOsMva9ZPkKau42YRu5uCSpPqapke5rrv/f737lLbKPo9bYlWzc
3/29g0nDxFZuMx60DoXis8X15iDbnOmoNHkGtVp1Lk1IxK1BuR0gvpzCQS3mMOCD
tFK/Jd07PyD4IxCvMQxFcWCR1hD5ej3VN3odmAiyGoAiTpA5Kn8335ClPvzB3jSH
+O+EUms38yKHAHoCSdQUVhF8nTpFAhqp1QMZ1yB4dw+kQZVKdgMz40rPUEL/sjUz
vbwg5GbkhBDvsiXKrRxoSVd63bMT9GxHAw91J5nlAf43YHmyDIsrPDCbTax3YRF2
EFtrCN8lT9tUINGetCegLRnnJ6U5AlhD8mU8vjPs4qKTkMK18GcHl+P1f5+eHJRF
qshGBTwH+gUkdZr279xuvkdwBWZ2RvL7F9Zq4iYi691NlDX011MAMQRXbu/kMenQ
uT5b2Yn4kO5HNcD+9JFEqrZjY8faOTOM1RZ8gHM1JNMMB1EkEed+mBuJsNkLrsEx
19DQfYa2UY1GcPbZ383cG81Ia1eZ4Q7IdbKdtR6MBybLn83Xwcd9bOQ22LqJ7z7P
HDFBnJIr9/sRGC3K/AKpc/ZRi6YffqnuZ+Wm9Dg+LfSWpQgDmdJHA+8jPsA4fJBC
ZfE35mcaoNHyeBtnrPLLaEK/frV5QorTsaV19egTdyfGWqoEyn33a/PfPqX+lmcU
LR+e8mLW9MUrgvJBapUl+brlFxIvYBNGXBFkB4QPbYhwVGEIE3Pelyadl2rOR3Wx
rGrQiB+Js9KPXya3X5wGN6ixf0UIdSkfWUcmfoEkYIyHYp/U/PpsDEn6fqo0IpFg
bQs9rP9a2ING/GORuMK4ax2Pq5cr6TKkAv0uJSHRfMDeOyyt9lWE+Npp94yyZz8a
67vYepi9jY+qC+UiBpgf/ajLRBRnL/mD18kUUEAoZZ8Ni+OgTZVyIJ7NeFKBbmAx
zMH4un1B3N3ixWvsE3IH9WVrP8siR9z1ZMWzAYkltgogATawHtrR9sLcVJjoqb6Y
IhhEi61X7TXZMXRA/uHz6oV8d+zfP3NoV7UFRKxWsxLJ/BNhmKDOkgONDSg62Lx2
gFwsnbfL0Xqv3hBXKMBbq2Ox5yw8Kn32Z5JyvDky/SoTpYWQfWBcwGAam2whPZtN
kSugOqUWnU5QzRChk4+SFIqvHoGRSClt453fPGuhPgc=
`protect END_PROTECTED
