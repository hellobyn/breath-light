`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fv9dAidTJN07fTugtt1dNEewDIE7JbzJFJj6G1GPUHQn+nWs9GICC8Y9p64jjh4D
aFy/n+27XrzYn55rm7l6hrVa24Z6YMrwIh+XLhr4gZDhSDKLO0cZ7hBbSZIO8QDE
rE8bTOefrF8cH0CzjYuCUHiAAtdqpQt4CH59qm8saaRo1dwbzMxfk8xS6014Ue9x
aGb7wDZ7Ydq5JPGWrJvAJysw3MBpY07a6kZeDtrhCxVuUHT+4WXWxvRXMczAZ3m1
msl1c+g0kDSvgQidC3mEafCZ5HloZTrVQ83z2OhgKVuATCpjx+oOg4c+eALTVIOw
XRgnvJXetIL+AnWDbwRWhayMkYVJ+rXiKmsDTxBYo6CV41vHcQXtjcmcOn4izZh+
JUme67kD3VkqUMWk+2o6A7lXhUoC0RRrqF41LpmDbNK5yRFM78LJiRNi3xCvrart
O/BiXrhjoQlXewHEq4WA48LoLtaLq1MRYjfx3O1CLfEWkk5O4lYwE5ldEn7UIjfS
1oFKj84wYZ76vOlmUQNE03CuB/29HiPjb7kUc4fz7CvPbjdJz3vtVn8qUl2koLDg
a6cXTkCo9SRIk+/SJzF7VuDDyzjxgdGd/1JvSaJjEHeQ3h7n9/yP4KeH90p45YC3
iSjGPmppCwdz5W6oveBwpmFVsiWy3bZWQmWi6NAn1HTlD467ZwTIO5X7LND/Yqy2
1M5GU+SMJW12UKSE/s8z9UfGeNrnxldI6P5zMln/lQx4MynC70X/BQzFMFXAEFvM
nSNfJCqFVUws3208vYCPKzKpDhre4oSWfj774w6mrRI=
`protect END_PROTECTED
