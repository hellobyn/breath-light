`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6txlffHxTXD1UY/s3XvYPoBRkWCXC4/i81ew4t9QxuT2WXTiKKj+J86f9/1DvJ6
KtOK/zuGQBaE6Rm/L2TPHE5NrzQ26ixw7PkH08giIGqJNHUE8o8ZvwmZ8VN46YBi
bPBxTmt8JVS2PmHS47enyo39GMdSNK1Wyevr9Ka2tS677rn6jpYhuLgDQTrbWO4c
3yD9ORjryjkDlVGFSLkw184pIEMZvmAJXHtlHM+xAsXLg25E/zsNtwWl3Qfo04Wt
GjYyqFQSALD/sJsO6ISQaNG7e8zIvA3aM5q+xmIQlMIFS6bQblC2OL/vPHB/b0SM
I3bNTFb2W66IVNGu2Zerfmn5kUy1MndXuVI0qGxVBBw7ymhX00amIFhiCvYupqmv
ssU7V8CDwCklQCdh7PIJhBS4PxyZX5H/ApXFfwAnUnEUgp3voMIngUZ+zxZor0Ug
46tgwoiBc9j19x4lmQeFxwrhz0wUT7QbOO6hgVo6ph0NN2y9aJP8vbC1Zuwk85Op
EJSI+dg4KEjEGCiWy9cRTNWLGee6cAKhehIz3iqEvIY+S/X7WigrLi3kbo5s3Jua
A+cfgY0J5saBv3gI2hXkx3I3jTenZQAU8ezMkFquaSREAqRdTBtkuWNYfd7D4+9w
g2cpTzT04iompwgBEQCtP9mSJmOlSYt/99ynZntCgJRmDqr7RGjAbrsID9EvQawW
OiH2R+WM46TclYmxIpjDBSTSiFsWnxUupnBqGCEel1Yr2WmG0QBkDRo5/4GBmv8f
nAoGlavctCTNaHxdUz6w6rs7WtG9Uj0ySzIOvA1K23T12FYUM0Tthkm0/pdbCT4L
hnuxxR04IRulX5NIXMpj7a3NnKnOUAGEGNyZaBH46kVv2wktsmRN1RGXi3PqF+w3
WILBJ5vWK5VUWH3ha7cRBHC+U30NMFfnSNDssKr2EGd+1fz2PP1xCS+ScYZ49tnU
GOJ62ZRBEvijPwWpNWvZdHjek2pKuktBHXg9a6/HgLXPGt91OwbQt8AzJeitmL3c
kKOdgVxOJHAJ4gNMZkPVBqMYBCJERHThjgMMc8aAKa/PhhxqWbaH0WQmEx8Tzwyj
k/ytC/9jSVPyQsW6kICCkYzkcOtzrpUq9SPIGMhnGOFkaEt9E1Z3bQr4w/qHOjci
Rbz1d2fomPiiPK32b9O/kgOzbQVekuiyGq7SHMdh6BR0DsiYEeerV4vGwKNCfHR3
nS54F2Kb3RK6tUGcPDxC4rgIngZ3S5tRaeoY2mjkMdnZt6uc1qym4x2vBPkuafrA
PuMcugnNe9623lQibhlR5/i9+rRYOrIrmsGKL1Kd7MIFJYOPLprhB8TR3fQ44R36
J5ZPfVbXfKmaL81m0cM6yyuwbqstCZ/31wDRUPAK/Q2LIz5I1qgorC26J41iyCfL
sFT3+luuT9zyYJnZL4SKQ5jqIzkhZrCLG/qaiOr3X/kpvXexm8Hx/vaArvgiNKHE
y0oF+zeQJFkw6LhdHb0++pwARDiGEoKCQnlk4xq/xhzqEOf+akfNvKpm9VvNp1TN
QyQNyjYeB9iQoUry5lBCGVksP+KaBNIK63gI6iOcn7rU9JsuSu/bs6KwBWosFY7M
MszAoSk9ce8hL5pVPVBdPtyn4fj23ym3+TBESadvou/tWPk7QphxbGtB/2IQ7MgA
9tHYNtD1nW0K+97s9D0P4vb3oz+SoSI6an7DLbX79+Z7DPt0Ub2b43gR6zc7s2bv
dUJAS7UjRa5qQ9kH4tmozOwH+2vgw0inv5GJuF6ULQRjcQG8z/JwOKEtguq1KYjV
XMNH0JuIS7wVea/HPVnyaBdveCDOC81N0L0rhdXN2OBwk/TAN7ncZPgTLCwclcdb
6kgldCUX7NAbTSe2Kw4NmS8iTY+2wRyzP31N9t3pPzI15KHvQjGfb5aUdOdsCgnF
55ybe0HCFH32bp1+QRDxqQ752xvdBPUNqz1rHENxjLElwq7Y4HaMnnPBfmG1X0FY
3cNLUygkv/GpwCkcp5TlK03EAP7cFSHRkBcID62nqL4nBlMcMg+t0WHg11sbT0WQ
BUayBJzNs6KrfpBqLrx68Z1pBkJyUh0k7hkW+kJaj0tqpjKOMLDF+jpVW0Sf+r1I
79eVJCw6/4cvySBizDgdaMqFxfJGBfVjnRyTY1WUhukcJqQdA01CtHUjXBPGoFVr
gKPIjDcV/ru+kjGJBle/RZpfgnkU1HGut8ghq0y4decu6FIOxH6XikadQfC5mILJ
P9Wf0PvmD+9IpNEahCeT0Sj1Za2cBj0RdsTsmw+96PrZ2I+S2XPxzK4k09k2PlOP
trBFXR1YCD6IyVZ4Jnr1+D9ynwgqh53eHirjmtyHOZD9NDr5OGJA0Tt/ZRxlT5/r
2UZ3jHTE5mYqHyKdZEIwugt2aRNCuwAQAumBdtmw6kS5tPysvD/iA2sZe6tkHXI4
Z1xQLj955eiFD85oqqmLBNpph5DcgeNMXYLTLBUV5yzvPRmV3mq3xBRdfBcfKJ4Y
12CHbA76Fk0TppzNkmxE+o7Q+yPqdpZ5U65y7pFybaGYE04utydmDBkQxiaosOh+
l4HJkoK9EGsmIeR2P9kYhqmKS15Wj/LAzcFButgdVc1GDMBEELfsFYg60gPSRuiF
D9oif+DLoIRGF2O4GkRrIzNSCloR+h/XARpKJ/2mknWGHGvBLlq7Cj5zU4i+0dtP
ETfPokoO6N27uljDnSopYI81dXSSZ0uOitwh9gSRGzvM0qxOFOPI5RkWEE43wHgt
XJCWKKceWfJz8uayhOHBSWy0TE2r3tayXq/cQ/ySx2b5PxVQNEvlMAhqWuALYTZD
p6jH4JlpQu6Nrith1dlRlbyGQeTNy3ZwAYbKlceKaH5rF0pkbbLtyV6wLMEdhTFw
eIyJh8y7ffDvfAzN/s+Wh5oyASxItirppMQyga0dA8SDrrOBvkb3ZvSST6n3gnhg
ncW0Kf+fCgNgG19eBFWCpwxho6GJhS7F4pCewzDPOb8P9R2XiTbbUKupQ88if4bf
svpjhY10a1o40us5/I2sQWIFHr42LPgWFULSiefdWOJXAmdtd4cpVq7nFCyDQGkx
h4trSk4TAMnAVpDPOgl6ismNMDWhYp/F1/bh42GSCBNfqCGdKdtCSi3gh2kcTQeg
ESvJh55hKhpx5lzSm0LWoL/wFXz/3wZAjZPB1SGjmQEfgJ5WK9o8wafLeD7V5NTm
cf2B1ow+1jQ13C0thfJxI8qczXMqTatEaKgxroGqtVQtzlLGPf+W1DouVq8OnL98
lC0oaVvwf+11kVRrG+lFRpIdvSgLqzZxGBM3FTzpaPoQ/myz9+eHArqjjzd0nOKB
7NSNCaWLTrFRGvQc99rgAhTRehQbLB+5rEtWzhnmqnKBrD5lqZbs9nZ7K8LPwP1m
hGRxDmy4e9lmuyft3xLo5KK0lG0x00HyFlCP0HSfjfXazITMQ+egnZKVhC9Ygklv
CSvEVr5vgWLXVIoT2ia3bT00OLzbVb6spqYdrpe9iRl8MxI9jDLkjVF1Cty0RAPu
AkCmPzN2c2zJAC9+mcHpRA1h5Ci/mA1ZOFcqVwyZ249tMTBuSA69OI5knLurtHVr
cwOlR8bywNig2R1n5V4wxaI+bulwS6rLYfsaRSpF1jegM3a68b5Cir43E177vG4q
xx3pK4yIlbPbfP3Myyf/KhmKkbohfafPmQ5JnnfzlHkOFAP+BxADMk7A4NNQUh+l
jxwKT3hsGYfsa4pZkKRi1T8dMNUiM21woTTNUKacdmOGIoxPqucOu4lQVBNS7X/n
n+5imKIJ7Elfz2atduoG8G/hA0RGxzcJjSwQeB8FpZs3jI6rmUADu//5bZdfOjgv
hKT3HwJWfnAPxoAi6j9nqxOGSstdQ1s/Ekpg76Is2gFhjlWUEYpgd4FznonFQPvL
KESEIm6KH/3L0bfh+mqXVyIOx4CCYcUG52mzlVExsPhGo3nNEhAUuqvGvKCwp5he
CU3TJIqSo0nDPHlKE7hJPvy56zm0iMCd4DnbAufH6iml0wc/lyrYpx1bYPF9MQut
BRGyxSCX15n5/s36D12klZ4qfNAjXAoJB194EVkzsDT6T2VqeyDQ7OhHk5+PEBNK
sJgdVJmFR3q0L7Xdh6jC2/XgUyMcxA3Nlo2S5onWegdgVQeIXfhg0WQzeq5md9dZ
gO+QDEHdT81Ak5rbwQjwCltvtbwgMImq2Y7Ny+XrwR7o+w/sYsV41NL5af3S+FeO
nCKI+luRpiy9bPEdHcvuOvvjHD4JBKPv6TkEKc3r9O6EJydIG1GFD6CQmou3Y8S/
Djnr58LMnD+ktDl2d90hkW+iVm3kDjS2PzX76Sa2yW1MPEONyZBlXFisOu3Hi3TA
pJRx0e3apfa8KEhqG5gPks86SusZe8/bRlXw9gORSmKdZZj3+JDvdIVJ9HtNwNnA
aOQ6NZSgvm9B9FPg5rGl1oxlifTMldrkVD8OJJDh4TK1MK1YB/QrNjrS4hlAmSBc
9yH0O8IryyXP2duw2G5vSSh8OGG1uKyY2bJ8yyh/AE5l8/Bj1JGm3Atpo4ExmY0S
gTQPyH/xJPanyO1qgVEOoWrqeaNIwqVYiAufwhYFOm+bnRY3UFhAvrWnOMJOV9MU
ux1zL2kKNEtuaT8teM9EYNE+kQmcBR6ZBinXa/i8p6ok+UYjcsObc4chwxdxrvGX
u+YQZEsuYWy+N2z1gcc7iurxnkwJIoTgXTQuKKT6q+wqj5NJ8WzEW9v9GRs4pAZa
lsGS+b0KNZgEqQzQ6x5ziTud1N49JptkEirmn7gxAeIAv/ldO9bn7+NiVDdXI1GV
FNWE6+S9YNmkE8Bod+o/Aw1eFZMJlLPl9ME9QqIGQMZAfmvVhLULBkR9aV1FnjaO
PT/kIsJlu8AS7KTpbxu9YazD/o/ijbfEM7ERscDT+C4/a39SCopywRaJkFFHkxQq
iXIAewZUig149SKRRvVbguuFam8BHBQg2rmVO5va+hLBhlRXoANtn9nwE0PNF/E6
x88X9DGMz4w6RoI66dGw9D0ofsUbqYYGtTxZne6xNuPb3GTkPf6VnYvqSHqhKJwv
VC6UWnQ/EzToiW30ykD3ICEYb+L5vxJ0qv5fmjtrKh1Pm4xH808uvDraWXGHzD5+
9IdArb95i2B5pVMhTZexyP7C/+ZQ8NdQcf//tu4Q1YkjAqOF5Mz4rSMFicCWVwgJ
Ul/xkvMyLtiSkH+qlhOGyztXK3cf8Ho3cGI5dH6atl/rzAAqvqd1e12dnSEF4tvm
UcU5s06ofu3xtBtXNDFc0AXHuPFV9tS7tMwUJIOlwjGqRiL+ZOu10+/BM39m39Nh
3eqg3qGEqNUIwBXkj5c8jMNDHWC40TZIrCc+rR5IwI3XNImSazuR6S1bTO7cDnUm
zEx6FdyViPkf7x77fK5/zABaWtrPV+zcEWPhB4fHwcmnyldwOMst+Wma71XkqbUH
gMBbKSzHPVyHJYGcFTRFXzZhpCIibxXIJpGA3t0U9GEOI8CIr1zKRbS95Uv2VBtq
O4Rk9AUxY2I7Jw1CHGgD6+6YzJjQiJOW84eN3l6/lB4KSFMw2Sp0cMBtBIesvCVy
ha7BIyEW3DuawjDzSdqAZkWpW+bhT13VJdf2nMbXYmT+dZAz85T5HUH4mGFFN1Vw
ywuKMJ096y9e4g8WxMkDmnOToyv4RlIvbB+Fjvkdn1ZcqIOtFhb7qsq9+IzHNNXf
suDV1O1Dl5ZMYma2c7VSL2Zr6uNgMzB5kJSwLzhX9SO+oxVFLBfN4JNdoYOMQJQk
Wy+NjMgxOLqv6afY99+PM57pICUb3pTeMrcfBnD84P9nQUiUI/l0eSxwCSLA+JEp
UcFdLlnVmkQp7noZ4ji2qjmhfjBc9Q+6JOVgUepJJFn2Do751P+LMyEMw8NsA/w5
o971dAyz7czex2Lbr8h9/M40SjCHQs6JQScRV5jbW182L3N6RdMIRFwqaI/lSyDw
nEu6A9XbqAoVNLKnGhZdUcTIB11ZCo/KC9mOJDtsCNlS87//KIw45k82IycZlwSc
CcEKZS875+Kpybz/IDBuj9FTwBcAJIum76kRFa1HXgsqFRIYCp0YijagWpHB/4hq
mjz/vRWmXveLWHmxXvYt56zoeFAZrNurI2ZBGKXLewCy/6g0m8zipJjQG/0+ZTLV
ZkuXivlE9IcT43DwWtoq7Wlj8zhdtcmrEcbA8gzRQK5qj2mQbeGuxC17xFcSmPGn
8JAHhFmAojLfNS9Rn41zU79LSvCbavC8YzRM74Lp6p2GI9hN3g0/y/d0BkS57DF6
d/9xKR0QnJNhC/dedh+N2jsmnkubE+DyEM+Jv+E0hkjtCboIF5QUPMjLBwZuLw3R
GAUNFWFppxqpA1YhELGM3/lH0v+i92RNTfkTEnIDcIcsx8OR3nHMDJR1e/fOzF24
luB1X7PGORfK2g+E6mN90IRWuEloqYgkKPE0fi20V66zvT4KsCHy/fKGlH+eNTBd
HD7tOm0uCxwx4HvPQu5Y1NlCDAyK9FpCtSnV8PODwrbVD5dZnmg+mtI3AyAprACL
VrCB901+7PTNN1iW0x+xD3GMxXRh96pS5271w2zhzGvVhv/SFSllUbDoDBMAmIlq
bdeRldBHYw0roK8E2Q/ObCJrxba7cXT1TLCCPGsjXQ1mBs+cWttF4f6Evb7BdGZo
KMVnPGUfRRSxJdj9i56L2TOh381zThAqjyihN446IUE7zk0t2Mo6XQBtraK0MnCm
sLcdNUTrSK3rNrHJ99WS5sVB7VSgL+l5wN9fnkgqCWN8ONrMNoy2fAsDlOn/rK/I
as4ZRBA+dViIny2zfVCpBGTkxkpUrxcVUH4C+hGau66yLk4/6hLHB30aGsqa2nlX
GwF2FclROj3zlXeSZyT8yKSlp3QL+MZPaT2jS4F5ZXlGIXf2pc4dFUm7ySmXp05K
I2cCKfjcS9zDjVk34lo55Crp04uQGIRkfLgfwhfP5LriPi4Uqp+jTMrw+5HA5BVH
qFpoNvHYPmfFJCzngwZ9/P4Ai7hDcZjS9rM4aD9mdcbTuDouOQCvaw6yprAeLZpc
QgEQ8+SPvcwCj/fmBb5xNDb/yNqAkA+I/jKK2VaF3oLymlcPA2/x449kVDZf+Zaj
9yIlgtjOEr9GOn0fQ+c+W8UYg6m2sfIiZaTr871gS5OS99ebcA28iCy0RD+Cf95F
a0H/WzAVANTfjrBI2Na+tmMBKvhp7MbRHaoCHywQ/0/ZK0hfIjCf2vfO8WhkDAfk
8hjw9DxbAPF7kkByyktxswC3aiAc4znZ/Ctujkx0v8tDv8p5iv0UYCVRq2yhC7I4
NGvIqY2K5ojjm3kblnxydOoVxejOwtZe8BszTE7sQF040xqpkL6TZDYVInAnda75
wdWEau0xYJLo4LjrTe8fq1jb5bFoz31zPJ7HZvs86mipX+aqR6qNg3hbRXMAPDJn
+oh2eQKLVXPUrEcTFCwMmLmPP1vfdx6mytw8vjekTzqwhMHFwutCsH1eED63btYz
7phrxGVyjtqTxxIH2V6ddG4E2u0ulocGMOfNlR1XzaA9WsARwXJ5KToQ1g9sODGL
F6o6twtpHJLLdsi+rbDm6zfvn6Qobv1YXbY6pl2tmDo/0O+Bdm1yUCTM5Dhz116z
clk2vixjqjJ9bW8CeCl8iHenOzLuqBJKSNMVbROekCPBxvVKGW6zlhpxUc3JOmf+
4eIKit88gRhZ6YJAzcVASJfdmVoGswaHeG3jrGAqYuy61RrAMqMXxhvs9JiLLB3W
iGeP/DVTcxQ1ZVxMQs1ctt9Z4dI7Xi8PcOAKIpDQjx0fK8J0Jgr2U2CCQexJ96Ur
0rW5Xn2UHbQQyrh5iaYA44RTQxvaspQYmXcyOrdEQE9zHga+rYYyYNoLrdCzLyK/
QKlWfEt3a8rma5btShWu3mJtZFJIDFRGNayX2+TS09HpvognUaQfjIDxQEEJBUPH
iK64ELx5n+1IMGhw6hllAbD3b/2n4de4TjE8S/CoioiY1zKWDIBnMtmC4YbbBoJU
f8QtYpTN7nixpeTP4FoqfXo0zcVfMaH4w/bEGkBfljNBIKHqA5hIe/QME4NQn5eX
W4PH7KCOr01+lUmi63Axk2l2acMkLwnkkzpD6XgSLifYN06U0A9I8+wrd47ig57A
`protect END_PROTECTED
