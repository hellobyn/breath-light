`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYdRE9mBc22+Hzwu5TGXRZF/jCT9zwa4LUPilh2lkxRFsqhQD367Xtuwpac8yZre
DSOf9WnEqKB0jnMYhUulqkeVqJO+5S+Nt2ogLbAjwr1B8b9bdcfOQlcs6HzG2hRo
5tmxBpBj901elgxmuZU1wLcgAya59Z6+ZVPdKaoGTkLXiILhLGjvSr9GLpS/r0mr
Z4E6jnq6P5NJxjN6wcbW0ijlq++cGhBAoPEQ080uZV6n7nynVNkEB4f/2BOLdRzo
9oNc9+WJ5kqzuQSbHlTR5n2DaaOBkzBkgpz9QIfysdmllQGQuEMBKOKmmQH34o87
Id3ka6/MoFqPQBkfoa3rs78uKL5iQjhcZUMt+M342i5NFsg7I6noSG6/p0moF2+0
5Oi5LYLQG+L4+lZSxrtrQYfci2CYDs5jvRc6k2iui8kqVNYtDgv2IGZhAlekFrWa
ytVhEwIO+xqrAxlgO0896TEmiFdfpMN6esKGG34DwpwBa+0Qkixdvmj2u/SYrgz4
adljJcm07cR3YYMNvJiZ1bOOx6pftoC4IhzthO8HngJuEa2Nog1CiOMdL+Ugigrr
WXyVfgx9J6nGOhulFBOBJlK8UentR9FuolqP/C0S8qLN6oWrAG4xt7vbFCF8GRh7
PsUxxVxR0Xi3AF/GytpbFsX6uxl+WCnw6elADkX/LB4=
`protect END_PROTECTED
