`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A+bOez/CYekJEtqcrhyFwQCZHrGU03i1pC4yTt1tGewOG1YEYrJej9uCVYl7hkn4
HbdybToYEf59iDhvfTdGX00DbqYOuxF0oBxN6p1CfNfJ33/0jBCJJn3EQUroGbOW
EFm5zQgNm4EYAD2LuYgJxqVB3EoIi4NHf30N7VQrU1JD1P+SSb/ViABFWMyPE1E6
SC9dYEajHvqIace4fIWcjiLnso9dzOMPZJ0hRt+jBPD31V+oxGk4u/nTeLj4smjR
4Y/lNEVSLggQfML2PIYkEvUehe8SVLu5Up6d1E6i1pFBBd9DsM6ase5i61KpBbzO
Q6nNfs81S9GntSC+PkprFsETWIBQmSQEywX08zpw96sEWfsY8HMEL0veARFMDHRm
v9ttyiLwh6Y+h0WxTDSxkzviVW+vvXfMw2BtqZj3keP8OMF8lfib3oRHK0d4Cwu+
kuwHwyx5/pTKtiFA6lzA/D209yckd3Onv7yVbOnAw4Csk0/eXAuqU5ziPTRCofil
l3k+TJD8fvvcX4g986gj2gBaryaiSdKJ1lYiQYlfkAtiS3lwl3eiW1zJ2/dovTgK
dw72FAfzZY9zJskiONKpTpcAwFJdq31bgkoQ/Ey9NA+hI9tRWk7v9Pl0LveTnL67
jt1V3KnpElfkiovk2ZYWu/dZNATkew4/JLXdXzG0usIrXvjhvJ3dVHqprUHF2sf3
svM4kn8bygE9W1HoZDGGy5i2KBY0YEpanX44d74MSCG4PpHUjNZ/o4ejhBKjDKkG
anBiIgj3FMqm/gWqyCZ/5sj8BweRgzFwfuZgr2KlCUdgEmLSknADtwvuLbGcbF7B
PhC/lZgGZGCiRi1b2enH4g4ORNKGpI2ZLCushuzDD/Fj8XWg3awNFYW58/N9+zx5
6eAh7baCuUT/5ED791BtvQfiV9WYb+fnn4YlC2JDsM/abZ/B0a4rYS12mpfVDvAS
AGwypuKooPnwnuaOGkHfiBg192zM/BLk0mTdIHrWj6hOt7lKZtvyAWlXJ4Ua3y2p
QgtuIEdRVYNn4BdFyeM63ves4vKxflnDNxNR6pqIjrmHT3NmxzA0dcJkOnMH0xF/
fdnVEQ/lndYZMryciZ19gNEnBDurqhkKhbjYZxZOF2rbiEn4kxcMNj6eZJjpyg92
FbDfa/yPmF16DjdouQ1rl5MwIuibY451V3dQymqFelnXnoVEW8rEonb721r+Oou4
9/xWItQdphtYp+bPvmzCk9LXKtRzQ5T3BwR7Bmj8lcL8YoYpdLYgiZegPUlIAkVU
yd17ceeHIWyUhB6055RA9KjchGemXnqaxYRU/ceJ91QHTwWbN2wy+w6HuhYS1kW3
jCRJpr3acfPzvBjSiQZQBqNurzxohwUGEo2Caqdbb8asETARwueiOvKLLz5B6dEX
ltUTCP9/4HauwG2uPiqQgACHZTcOzpbtM3WgM7g/qYJGvVp3KSlieVgT1ZMmjC0o
/Ny/0Oq6J1xldHmQagFbGCgDkcri3GktbJy4oUYYwrfPLsviOnmeyZFIn7O3Kl4P
lZAw3a4JlWajMY9cAvaacJyKIJIhTNJ60zwOb5t602BjsfHm6Ro1DdpSYfulf+kQ
`protect END_PROTECTED
