`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRcVGp5bMS/8Foxfb46uNvxAYGQQurh9rOu9G5lnhSdjJ8fh4a6esPveVAGzKHEM
Ou+plTLH3cIDy19LGAH21K6f/nzzkBKjfiO9nhuuvn6CU4WTwlGpqWIOaGdHJvEL
nRuhSbiqnECd/qujaXAKomHbQ4E+M1DbOdFuclydKmmXdSC/jFKZq9+iouuUEJC5
iSP6AK9qiF6++vEBZiwUYelM/01U3Itei8aVK0vgX3ZKBSb6LEnazshrM5x+YUmB
BrMUyVmneKsHguon3YiC+yJlMKkSm1V5+RMLgcEcdDxNqDXSa01frExQdByRV6kY
M3kiX+InFujfhWWCH2JnNIIAxllF3sxkz7b6DdVu+hTnNTeCxc7kFYwlZK8G/fGd
`protect END_PROTECTED
