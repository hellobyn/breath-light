`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUqBBUGHXkF0wtJ6oenEr7XtyuN7rVwbOBhG7PXtGWL6tBmSlvZmP/qynqeSX7Qp
s7lLP/lC1mb0NOo/hIVDcdxOqDrRRtnrxySxKPhCrGqj1LiPKun+HPPmBPigpkxa
sVZ5ufemm45zK/bBnqK74zfgSkNIFr4WzUrd4k2D2Tr8WRUeSd3Z3ifdfKgW4Jz/
NJ1U52hjHXJNnP2MrXhalnB6ogBwBb/MD04OFQwBLtwno9W8n7hymCeoOpnfwL2s
Jog60IbtOWpEV9l1cvm3efZbEWVs+cxntknk216y9q7oghULS5IALV/B1vImUkjW
ojPaRSFobuA4wwzcla+5uoJKgxNFNgj2uh81RrhwH+zwN8aQbhXg01RwpTeYAV24
4n4pV6EgVa7ivwL7PxyfgFRYH5dHI+YZJ3GB2qQnUem3blrbuuqPa+eDhvXRADvr
zN5UXGASnkNNWz/seyje89Sd0Tu3VyhV9NUpfTA29ptukMW25we3HSRC4acwZcbM
CeKE7lLyLfDDjwMdFWy4caxKf8exXJDiOXsmCO0ovOdhMgz94bsQ6sA3rxzfLl3p
KOr09Qml28omKhyD2XxuVGk3/9VV1e0Hf1L6efWhIN33FpDyf5cEHPBbiiZ1gklO
dJQccjTW4lZllT29sVyJxldP5myBv4ws/izfsnMALY0eIy8iTLFJJ7hNG8QWopYx
xfGnGHD+pC637KUDPdXlf6YgGYt01ESLQy2t2jAsibRUUdLz42LgtdN+a5iAEe+/
BieSjfuvdZaD0mXDE+ublDg5dCADbWEr221pzMfwOIEMfqQ0StztI0DYp6WZWCeD
9ERuvn//w4LKd0ilc6owOF0ztnLLcMZjVPKcIDOD3Bl/5HEosmcbiywUZPV2icxt
IJ8AQDH2+WU3eBtg5mdQRxW3lMqDMMjKqJKZNXdwVd1Tk7QL2UOVM5XwgzC8HGiK
p/wYbHbViZEdPTAg3d5XGF+Trv5q8ZyyXnq3E2YGZY55rrASZPgYuw+vOwSb/ApR
k9h4DPqNPnvTSk66kBLCPo7p+Vc2yLwCowjymdByCwi21IshatPnobbnMtnMk3GT
ZM3j3BCLdeRBdMuKGrSWiAt8r34qYjynEb6qL+19X0GKIaXYR9hgHGc1GoMZhTLe
2QRI7n7Hsqd2k9mUOcAqvLB3g/fg7ef6joAMkvnwkY13ida3dCESqtALxFovDuWX
Qkg7N4h5Zcn4p2DOf7/6ZTV6pNMmXwfJIB2AAAtHKJSbAXAOXVkLjn3pCyv2POIn
70geHJ+MV8ygFHOev7Zx+dwbpqGJ4qVJ5hNhSpLSMysnKWmP1kXSTp4qAkZqAb8e
LydLMARjE/SOyAjZczwEmEPpHkbtZRtcv2MaK0BrYtZDmpJSb0Zt8dEPEg6GKzJA
zVspZiY+MHcQqf1qzNjKBrMh471vfwTpWxrvmXkajjUK+VTxdRwWI1TE4oR23OO/
BRhgmIxUFTMPqydt6wiFEWcN+0vdxS8rxpwCJmnLKjg77u5h4lsDDjWCdI5zdEj+
vPay/wZRMx66nnh9nGFtLAfOQTwHtekxgxlpAo2c8V6Kg2dLumlBTDQnjFGKUZvS
MmSJcHelvdKHi53v5o1mTRAACJNauBj4iXBQgV/oXb6bhIUD4zt7xAFXdqv3UjfR
hBB4oqFYHDvJ66xUxsD4j7cn+PkykIArjNOPxuym2rz7dd8UAHiZkikbUST2W3Xz
bg+GSoALq/8GXUGEkyGuSFK09N6Wpo2e3+foFHWts4tbp2zhGk3iFno2UXZXp2X8
PXO3rQstK2k2saAFpqoHKchbjyMUyF5xn1xJjjA9F0XZKx3FselFuwjW0wbKA336
iVntOMq9g+EVw4cF5VszXrH8Ck3BZTYxhITckUg2h6824sJgHYHP6dR4HPUlb4+O
p/zpUyp0XgiaKgmJZEHrBT/B51M72MP6c/dFqPoq4DQDnC23gj50kxu/Yhb1GvQ2
ms7x4o/GjdEB89Q/iIi6iHT9ATyTGcTiFezf01x8z3I6gqbVhhHE0aPlMEqYI1y4
E7k5rhW3o1hl0FEm6IazEiP9hWgHV33EFFLm2LkSn94M+8zHA6L9adLdHB2YVCCZ
1PdSJmFomto9Vtaa1v+AL1qUdDU59MfqJi/At3n4K12Dohwil2jc9yZIzlvP94hw
/jG4NhHZ0NX8b31ma4z9GeT6lvcrR8jBLoerVloDCHZENDp+W1WkqtMw3vw12Obk
r6XH3QQrURnmnMjU1h3V3NDp/ho3+/dfehuaJWFxWwd8LtCd0OlAiA+ix+D2SYcA
JYBq+VyxqCswmzNtWAJk1dOpUoQY4povN4pjBAWadFnfg5HY4iEPoEnjCw+YHMhq
S8GNu9gj/l2eoZtTLqhJt7V4FryUtcSiKFdXVjE5funNWriMwDBQLU0/gD8Q1PD6
bjuHpT3c8J5yb2C7e57EiTVFaG3ySvtV2gBpnCHC7G89W2O5p8oOM8ky+WQUJhPJ
WADyBSjalpaekOQoXqBKzADi78mN0I2x/03GF+67FvhMzaFfle4aNstmNQgQ6WbT
nDm+84pN3v2QBW7ld148VyDqjqlR2yIYAo0khKOU3B9yBUMTJxDn/Fu6HzGANEec
g7rZWzze807COczGhxI+HFkcuY70SWyhc8DNxrLyXL7GQ27Qj6wAbn6VvQMpRUYe
bxt8ykZBO31RDdE08/Q6xqc169A3bFKkSYJ45QWt9aPmqvk6z5RpO4SK62TQGCvR
iXp/qgkVD5HpzUEUioO1KFfgT4KRdGJt6HWGowf4leHJldmonfj6rZ0QOImkUDYX
AlrU35/KzaYfkV9AGhTy4ombtqP1SvLy7PVgJXEaH00SUpYeFMHkQ3tC5Q80jGXA
geYzd/2pQnhF9B7WK90kq4sIFOhSUw/5+EyP2xD3fkLE/Ac1eNd2vLMtqCIaOppW
YXtLGBbfKmU/J8MpgKkBWvIlKZbf8837f1HNlBm7Z2lQ5x/q0MXoLC+MN+pVAvi4
Em9nfXduSOF00Z3+8J7nYtE7Bx6L/3A7Pnm4pNwineemtTmjAkWem3QwQ4+45Typ
jG/R8gBvaBmajDvcj8Tr0GuwmjQEBOn3o8Qra+ob1XKO6GG0sEYy6yX5YY7QLwqJ
k0XpKoov/mJgnzwCjNG2IkRq0NTCclC/sZ79EKQ38MPe+CzxmZ+Tyvn1WJC4w7jz
I3LlXl+Uj7tKJxImkFcOOF5Bq3Nf1gfavUGvoBQG9oCZzu9+A8eQ9xT2zs863DyA
Xc9f2sx6qU//rnDRkVFjg5kDFx2UZE6Mm0hloP3g7kLOiTuHS1b8EDYR+PfoObef
fORARsk5gBED+/lp6DpW9ehpdWZ2MyplgV3H3DVk8/Cxs/lzibUXFGyS3WUPmQKz
LFxHW4WNKf7ruBivHHZOX5w/Eduz+ghmx3X2l8U2zceEWXyxReLHAd2poay9iiBK
2XYBLFUFposB8hILAKzv5w7P4YaAXXOdCa/Vm+WFGAEVlt4Sw9LaM36p7rUiNRj+
KvHZQBVhspCr7vf8THKNhgnTrYlRfdSSdvZGrQ53nmuZgADdsos8KH3NqMjnBeyi
jwizIEFEX9RB8WRFjCZ9zVhF9tWOsSiIULX4ycSFcMG4UK1DRuNA2l58yJTEjVkF
Sza80D8ifdQBarp8ldJLQsBtzRk6xZZm2IbiRGWWe/sIBVMJrRGrjYTu88FC13LS
15+G3AIGUDX+MYmnbcwZ9NvLhX9t4hys9WzyFgcjBTIQRMHYrQvkMcBLNuIXezqi
AnctV7g9EHJw11Yg8v4sfq8V87W2TT8q9/feyPUZLEi2lCkNdZj/ko6q9edRlMm6
wXF+aQNQj0PVdRj2r3a9BD/uqZF3ytrKDLcncivWXXlw5kK72KbxzIGMaoO41UgR
qbjaQ3u4EwtrlZYldj1chqO/+Rh8LBTagmJLUhpDRAj/PGSuJKsHa+hWZaKfpaTE
8ye3aRtslhNjK81R9w8L//neU/Lm3ZwG3IlhIX/x+VGE7/iZCf3hI+XeN4/N/r5Q
MJUpDrM+qpjGAoH68BmQZFrM8ZVl7Xtl5T/7h9vfVkTMpxCrFcvUyrLzL6/45Pr9
dd3E/FSzcdviXJcZw/FYkU8CoJnvf1L3uR7zPxdQc0Qw1YFRor7WvUjfx+hqPSSQ
nhPFTktpGb+J7RKVtsNnVJR5U0B/Oy/eAo4yAt5P0ADT7URLYE8kTMhBR+YmuUzN
7rkrMy7gwvM+aNn0M82uGnF9Xa8oCV65TSch+gKreZzhiYkDcNER4/LFv7orhZkz
3wvdvErtuf9DtpBq3tW+9SvARymC//N6oHvJ3d+FBL9FupeUURHewSLy53jFxt12
oJ32+OeSIanb2K6jmkLtQ9qzUwBBapLhXcLpqvMcl3TOKyCx7vGlMdVpt/niiU2c
5NAPH72Lw9yGuY7ANK3B+ZeboPEXadDMHklEixfVnv2NIk/+dYHmoihMIuPUnPxu
+wlTaiqaKvW4oiQ4Do5iSgR9aUe19mlmjTX3MQT01PUM7CAqsa/6s5n5rwWVFOGv
axkI3d/a1rBMPDqpCOzRJjzfuCPm2PWZ1GREgk6gH4PGhC5Qnsjc/00hganWW1q7
T+xktGvjkiIUTbyRwVZeCMyrVLHdi0FrnIag+SlgqXlHMbhVw+jdYHtYlBtM+Ala
d/2uU0XmeoeWxajpTouGiZr/43963Wjvb1VvcI7cc1RQhOZ/DNFQX0Oduk7p7HFl
xWkCI/kMbyLIuG+a7ZUJd/oCqauT+IrECpxP71Bdtx9A1QUjw37YgA+J5VOY52xz
JkteMKPG0Vogm95eZUuRfrvbojgmZ1omtu5SC/8MZzN80ayVc5nv/RB+LTgdCK9Q
BjYpBRL4myGqMYTWbP4nNCpMxfVPDZ+SpUlh2NzMYFv3wVM6wqFVsbqZaYDU0aPD
Rf5kbnHJQL4rzk7aLxadiefyNZyaJHWcuNr3qv8xvmGlqsHbI6qj0QOuvNRFMUp6
dWUNo/ukR6G7YH+dBpGNqGKEFy0cQLL0D7l3pHxAuecWMB9JP7kjUrXbtKjGcMv+
fB2x3/MuzuGqiez7Jqbo4uxdeNLTrLcJzqr5XNaj1sk8TObANfd2w/vML/504Dye
m0OAnA06aX96kItq/o6FAXUQGEJ9+jA5gpfYDZu6Hd/EtrZVjsqC++39uWZiogXm
swiUAuLL+ItwUupRm4ew8nJ1Yq2thRSHPqktJNy/luRvDLfAa7kRBL6gGSCqVQgH
nSbWRCTq+SUC20hnVKdQ3/hfb6NlNn3reajjFAVo9W0a0z403zPILbj2rus2trYt
KxzZghJdx+iKQNtFLuShzsS4FNmcGjHEBYAtmIuJCj+41igV+GhdOAlzdE1cjBkX
F3rT67ABMAAX+gdwaaBRU9JAbGGVgO3r7NzgOxHOS4gjljgfpSDFkveNlN43/nQ6
D7Rk+SGRtOlFPb5liqW+uVNAgqANMqjff21eRUS9EtFvsqekO4d72t9pwhupEEA3
TaoCQyH4U8L2EKwBdV4lawrEXf6KZZdtG+BZvlJRtqq2T3hyKvnQEK83SW+ZQcap
uqSqgeiZ/b6hI1OnYi0XcA4PgA5CUQUaoOGMRTXE+ZfuJK0Sw95+P99/K2A8IKMF
/cG0ANEMHqV7HxVdS+3SxUkCFN3VOjB7/NCS2HtvZvVJi6fPVJAKJZcL+2F983i2
CTiVdI98qhVRG/RylVkEKoodc13nweud8Q7KP5Rjbyk48evrJjXLVpf+TiAeTlxf
ULNVWqpCYfIW3b9VCJJVOsuLfgfffXXT4VePNHM6ktYmKVs/K45a4FHyw/zu/o//
7Xnn4jB03vOuhSPSWHMaqrr39Bvp25W/G2KFqE2OmH8BRsVM2rqis1P0pP9GCtPf
DTTa1yLA0TfQyfMnrkaNrGQE78+QpDea7CrWEFztZiNakpueFY+uIbzAREJsohB1
1bt4NtaVmFl+kLdbRW4glbm8BF8M/UcpHNLbQoFgVB+ZolFC7FjigMjN6RY9nnuk
WFsMGcev60TKYxqj7IS4KOhRhy3VEwgkYmt5xeXolOQHf31PBUYb3EK7cBTjxjl9
Kf85bMbE2/IlukjbGrXXcfk0VJ0uw3GCjUW87wDnTMUEw1OmeII1KyWve1ERr50h
gyK4xJSEcnVl+vB1FmM+7YP7aOdghMvJIj/Zy37LEk5k9I4FldOKaoxwtxpi3yXs
rZ6d4+FPnddbLZMgtGU29/6aOahTZdde59G/CsJl2K5iqzVjw87UxZ/nLNaRzX0R
771dvcG3FBKpVIbp1yogI/+xvsMZWjIXVhjJsi3vxvR5X2JMOexkWngmuVbNlt41
ExAqEJ26Gb2A/vyCrGJ8g8ZSXW//YENZskEqrf+jplcUHeoPC2Bf61JuamdMSXwE
eP8OMDDkqt3Sj17uhCYY93vU1AzUb7V7uGPP/vNCOHPlBNcJwCRiqX52LvB18jRn
geRdfradggRiV5eta0B0kO2MJTjtbxH9dxcK1QHcSFBm6Cez/Yol5JUmqhrrAhUA
grZl8zN9XfjU82sm98qDlxodHGBn6hJICRnyKGe8jfnKQIFfWZWT8y5nCYFXvos4
vKveV+ELz0nv3QjTQpfdOoBCFXSFcz2ndgA4W/PxV3DiELvGL3LzbiTDGGigs2dr
wVifltZnNYmJ1CLB68OHcCcrLHZnfCI9fjRvOOy2X1HrnUxxTqlyhs8atBOU75ic
FEVJkTVOdbawoQvjC39okTG926ILyfO2zMfxcUh7evyRx5TINwctTH3LHgNqsE+X
sQKd//zTyGNDQ+5hgylrbmlOU5V/SHS4m7HJkUxaQARw+8AG2lf1t7Ob0BlQvW1U
0F6BFmk6knndIYYznta6GAYf1BBM0ZzvFFK+Nw/pIk1+kJ9vbgl4EiHmo8YcdwlX
PZoS9eFMnX1MrAGNE0OL5/uPqpIEupSlE2KNxRNqbqdWzTAu3EMwJjnZXUfI6o2f
dcYQjOiyRf4fz4eI4Xwsn4QR0hZDd+ex7ogrN7meibX0usHy122uWyEkXEvmo8Wr
hhnEWudsTXQrz7O+QchyyNgow3sMhZeQ1jathQ3BmI79G8UG97hNmQZkD2hRfo1T
QNpVHRXAMbfpz9lGGYDu1UbMaDHfde4SEWenhRXTY/Jh9WztUVsM4m/N/aVDFcBi
689OlMv5hDClq0p8oUezVHn9Oxl8gIXLnu1xTctyRZ1J6nIIxi3mL93/LvJS9GjH
4hMQsr6opSeWhgfclO/yNykAMC6JQsokndJzT9YASrYvuDiJnf5omz31SXGWDK/q
Wzvvt+PqLBEN5SwQju+uk2cynwe5aeRXyhXQycsODnz/Hp3yPtC+vr4UuKqLEqWi
6W5sQJyLzUFSM0ijfmcpnOf1Sf5AB3jErwW3w5p0NMOt7ZTJCjTR3kf1Atl1UhMn
eR+BzoC0WKrKKJH2qw6aWus5j/nghmTft4I8Lzm0SGNVJuz1KW7rUxYeNK0N7c8Z
OA1/iiJdNHZyl6EpeNjP9oOQidnhznGtM5skVQKYK7ET6hbinSVk1xr50T+P8C7k
KwZsHM3+AR3P3rqnVW5L6TMiqv/EezzuxsDuuE4JDiCXLfjIN4RafY6gOggeFz8i
y0DxYVVHdeh+OsTC5Q+DUcmCbeQvKIDGmjoNwc3C/aAOrreNlfgLnS4ZmBMRYSWo
FwzZQrNcMX0EiEqv62flpZ0lLIJLsPkDMAMPfkquodTDJvhHJGVGaFhCHyvVL78F
3S3ih7FFyZtgrYVUFbLMvGnbDAAA8HL9OG2lLYbwH3/xD7w6I0p6oT+BOfxIweSA
XPEpxJy+wKNnfmIAQQlcOIqyv2xoevZj6GpD5u+UHTO9jBW+FE3TWxFXIxHZTB6a
KfIhpN19jQmgVJN3yZp2PsujCqigA/6439TuNEM6g3Trjx6CeSIXu8BcrP6/hbi+
B7q5NiI+SONy8LfW3nILp5ZS1z8mLSmoB1VVdHh78WpVmrmdPqX2VeJ/lRKR4ZNp
vPZm2kEfpETnC3eRLKqZgRJhFIvksEFSAc8jonN8JJOBkVSdtVW2qx2+dVl1pLd/
fb2DIsYSHpPMuR1qsZLfACgo5Kk7rlioyUWtCt2RwYRYVzhK4ZDjMYkVup/H6hlv
PFVpDiczuHtKQhlMmkL8axFpXIWIDnnKeurpxQPEK7i6SGIq31eMKrUfbKU8x4Mk
XqlzjnlSe184XgNGDXSnCCObZZT/fmJop/STTDm+XDx6bAvBdS2Q35pQt67lek9y
J+IM6vTZ98YZ/wZP5cd5aP/PPjVrU0Tqj+x8sNRv2qvBKOfiQHkhuZzsGajga9mm
SU75Xomkq4YfG2OIdSjL5dKQ0yVuG62O/iTfKXNT4K4Ug16v+eVJ4C28Llqz3q3E
HI1CiScgMGUAWmVa1g6oK/jXEzd2hVCoAm/vjU46GB6P6lEwqJwQDwkPS2nKhTLg
ppXM2gTsZvfyU7O61LP6opuxfeSonaktznFPkNcHOy1gE7yfFXBywzEkfUgdc+WU
bhN7hYJpk/R8OzO2e/AyFbXL2XupLcQ0lxxIxfQ7TyzjvYBwcG9+gyPaZc7yhEMK
CbRBg5uM1FFT4z5S9EzqBWFzDZWpX4bx2XZL0qoq7mNGJH/T2NkvFLfGfR9Ky4Ot
amcjl0cSBEZR2cNxcUqkTIRQmJKcyiG/XvgJmYWAkQT3MHsjqAdhTw601PDLa18t
i7ssX92DpSebHYeHkiJTQXjgrxUgLJVAsDmRB9tHqlRuJn/FFpBOiKYmk8qaOktC
AUDsWck9fa8Ajtwjl2pYyj/twt1R1g4Fi3jTCbEcyuVKuKLLtYHMg+vRdcIvkQTD
8cQjlGh/bAIV++i01oOhL1FK4DaoHj2mva0Wyic3AVRBJwUcsSrxUVPUmMbh6sQf
rExwywvySrO9MzbsKB3Ifs60K6UeRG78RYv4d2DyuUK+816fDYwKzD8DQgV9dySu
E/uQa/zHko6LX2bXdo7PqRemeTXiYQSFr79so3KNAC0MEZ0d1CEWRP+Cb6bRGYDi
bS7bx7UsiiZUmYj7H2EoKt1nNpG1rHFJrwLE61ZLw1oNajOT1AwUJH3nYgo+LAhq
wact9SxacPlkzH6VRZbhgdmQtcWz3mNUuY1ijFoI1llMCtztxdN6vtg4DgaPfW08
ox0So5GEzbQL/WSuF4jkf6pK+pnxDG4c9YALmP58AWT6+CnWJ0Zq+pfzhqq6cpka
w2OAoLpP/GYfJgAiJvY6QP2lKZzabSuZqdXbGimWGLO9Nye3429sEj8c4b4PbIw6
ccUrH1HZLsJlbzSolLfIyRQRAAETyT6oqz2ih80hC/K9Pa4M0S5mEwkg4HneXkc/
NfZJgw9CaOClZEBnc9D2PNiEn5wohu6eTxrV5glnvB73DsA17ybniJPzi8ivXUn7
VbDWvaWEOaODI0jKTIjG+9+KziXBHilqSjMscbXdBk1qez9eNGJRnoUvXsk7qMtc
0Kkt+mPZ3bua+MyZcU+LKttDEWlyJbSglh9B5l9xHCWU4VWIV0rDAff4P65EGfHQ
CCPyCyMQ3CQWFZdh85t2T58tenIe80N5kjlfbehZYAQGeHEq55LOWAg2T5knBg1K
7SOOdq5V15k+tnrqvxZ0cmulLEb/3CNmpL4fiIeEofd+J/H1m7aI23BdTy7MtNC8
LiUW7RxLBF8pRs90ZgClRqARPYCCbt3YiDOeEw52n9BpxkNMQGex1TH1nwCyoOh6
R3wbg9kWnmn5Kkj82dznRsZaHcZukG6XOca01b+8JmM5PO5FKYZBcI1Ng4WEiz4D
AJSpmi4Y/c/Iic2BTBFpF9NqozIiPAWR61I5EVqobDA=
`protect END_PROTECTED
