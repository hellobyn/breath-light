`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHBgmP4PA4j8IwxvMq3vUJgUHEHozz2JgS1K4O2KHmx35rMYkPSipv+/u1DjoHY8
KuRAKkO0R0++KKWk2+hH07fJjF1u90x8rSs5sTiwxdwoqF6g3hKyT1JAybd7octu
cy6FBX5LoRf6V8gfmOT3RRnhDy2zGgKaVDu2HF/d/Og9ozAVEOSdbdfBV1apaQCt
brdBGkjxsWn1Vs7sOyy/EGYNNxA+r+uuNlntpmdCEj297qnyPsFW/EA3/zHfbC5o
g2QOyo1srlSn0aLbQKFYuZrXyOcMujc803oI31O20Fw+rgR1p6IRDXzPnKTZmW/9
U8iTsBB/aq4mwiBIgp3nE+bcigvHngZyQpL8BU0nHXAAEiZ4jqGhEf1HS3T1ZRQR
YRUWGVz1q0k/eShqjgKadaZ5xJ/XAT1bP0t1uunVJggEkPLEojcMd0a3t2lJtPy2
MYlPtuWozJfFBjfdxvDrBTDDwzSuJVd0DGL21zCsQROqMu+PejUBvmhxAZ1sPLxY
hSukp94gkVIHtJ6UvAlnSkIETHYz8qfCXPD1NYnnvqEbPVQahyZBAutObyQdMB0V
ob1WWR/77X8O6D1RLulJABgbuT8np8oQW0fE2Dl6KwWxaYZV5RpCHxaz9HbY0AfM
oHJcd0dUVaFVLu98CofDTemppriu8kittdGREId4nSXVs+DBRf+X95bT8xINg7hj
rEhXjTh7x0LBQCRHrt6qa+BaUL1x6MFi/Bgriz16ksPPdbBtXvzjf9i7Nf6RloYS
SiwRmE1npzCAW3k9P2+vPuAXoZPceIgd4sWGBLW3/ASrcprmlee1Jl/+TdzidgEg
ImDlGSoB3e8t34RxeEYS8xtZg0Azq9rl3Bbr2GtObLaDFNxx2azshTsOaXg0HxBa
I56q+T9yayWgVqhg/Fgdd3ViqufusgWaSkLAX5VORcH/Jbg7lEJ3E0WtdOe2AtBx
eoD5CCI4C/fbszF00BdAUa0qQUP3WmS2YjN5BMURVAosvJtE4e0T9N2KvJNdDJkf
WyQWeblGLor5urxD33fF76KwjCJFqvK5Y5sxeQLYo1FbQpGun7MMz/OwTLc8q86k
`protect END_PROTECTED
