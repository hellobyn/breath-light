`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7AyoM/YbM66N5JUifjxsGEqfCFLaq2HDqVy09GEDcUWJvIIrnPy6NKOXmw+lQT+7
kGRveYsf7Nyo1PyiDei8/B8cL8KBjsAxGUlzkrxix6tS2nVwlpcSdAMsDWoQCvwR
3Bf9C7oFgKhdS6TUTzYBbRgvSl+uh1+r9AqF1nzYgnYRQqEtsF9MThqF8ce1yU+i
yBAYv4WRGxmz2U8z8c4o5ckM4S+lZRpLDgYKwGavf5+AEEh+Ch8oX3AEIi45DZrF
6LBtXlyl/kjHJCgvOrjt8a6qAN31IDd45sEg7cm97iMDioWh5JsIGC3VG/kLAlk6
L5ptbi9jjxDuW4vEhgV3S5FIH9lKnl444sO5AayMSVd+bD6f+QZ0Iy6RN4uf2Hs/
ecRlpdySPW7ajQ48C3eE9ehkXX8pCi+PlIwfSV0uwceT4L8VLLPLvQw0ei1Z5ANp
DSqvZMULwZMB++wAUe56IdxpgHHOGF6HKLCtRnKCBpLvGzCj8J3MRMWTFf8onQAD
mUdmE/er6U2/HgQlYwtNDoFvUPBFXYGpa/J3XGaMfX1Qt+sZqGVQD4nr4QZ3HTk4
JetmRlZZ09wGVTLm0aUnf5gOdmXZI86QeCcGt0hKcikTS80oyPDDGVt0jZQoyp2e
KS4rYsvDw2N5rODYKz0SPOMovz+nzZaWlIEtn822DvEmjc+Pn11T3lATTmdMYktd
0bODXDXm3pOnWyoF/cc5015BTWP4MqtVlWiJoLRJ8ieXIVY0zdmEGtDHJzrdIc4p
yeFk8RNuA24ClD2KIhnjgheWjaVJY+TjRspT0RSVUsitTFkml7GWU/cVcuxBP+vR
9lpNoXhr3CPDm29pwu31dUTpRQa8sH+yWvqIHsMOMkPr48zCvrfotsL0p6H29c3O
1kjWs7hUcM93g0BKNm/81bieSOeBPwCL4jWfWUkZ1iHcbq9fOpTm+Q/Ne3aee/26
hCeAb/fFGMQBSRUOGz7Pt5Iasc2ljLb5zbexrdDmflYUoG0Zij1xN9bUWupUgpVv
pQwjmLCCSr2OuU+yKw4bWaibRJc0xI22dv3ckMB03IgI85yDfQRlGVNf5VMvC+Cw
YY8dzR8feaeW/jCouD2mHWw9AEulMWY1OfFeBBcybNimgRDyW+8cMJ3rWn0Ha9Gw
RR+xqCLR7Tnpy0XOL9C+NV3FqaqWr5XQp05tfqSt89wiLt3pRe3aFnRQ0i1gZlov
h8tPN7MuX4O8mnac/QmX9FQ3uT9ibakMcDH1kAvUNhS5x1P2Ae+XWuWe4OVxP37S
HdST6A66rFwOooWj4Te1bkMV6JhRku+QvBOzxq06GWaMOpP879pwqeOAqDSkrARE
r0qYNqzV9M6ymA+OPx02xBjrLBUmX9SWYazcw2mnHWC1pNuw8vtU7DTzajjYmnxR
JNIzZ1sHtpvmrtIR48Az2NTa8ZRy3sMcOQaNo1RaLJY1SdjUlSZuCOIJJmTwODBG
Cm7cEwqC71mT/uIgcFIC2J3GLxNcDydLIdOvR8gFPi+ZKhZZ/khkxU+DX+SeRtPk
Ikc/ZNcw7ArWGEt9LBHN9cIqMePwOmWNUjpvgM+CaEPRI4bsE5ssRytjodmR52O2
3mCTD8ywHFKQGMZYKBpht3YPRSG+B9xan1jLyyv7sRa5ZCjz4/ZlNZHVnWnBYKoC
OsKjx/30cdSdSsPa2dt738PflkLL7DZCNPkyngcJKYScgBH46IZe8BY5ktRzGcKz
aZO64iZ8ED/UFjsR41jDhVeBijTtFiI1tkJvSSx54l3I0pSssZS+X6NSPjQ1F5Mp
yocLpyWcHfOzOdoerJsoAEBdTCWxZUwKr2KEDPRwF6DPM8rolF/90lWYx5LD3Ovn
DMU5YMrVyN6zQs2A80vufZ7UGs6Xe67h3h2YskVVxj1msQZlDwhyGRT/qn86+8Oe
P9OQzbNnDsXzBv/misUveKlbn8nIgNTeqH9sXWJSzGVqb8uvGPzldCFNcVGwPrLv
/Qa1H0dXw6dXqc/G8J4OlDf9AVD+9ZJaomjwDyo+HslsrP1n1SOFTmqgiUsLps1C
KUsQ3OF0DlsCgnKz8GD7bqLLc71o5/sDk64dimp3Uf/HRodZO+oUrId5jSuSFTnx
M2fYlcXuyu2ofPuu+rzUI6sCZ7Dvm2xvhydW0uwQAtpJb2gQrvsit+lkF6Jk4pkN
c4VdUaYzdbhkS0sSyCqGkidv0IuR3HzE4iAHJUKt7YMP/92T069vh/YMJ3Oi+8qq
vMxqXrScKVD+Q0pWYco9lXgWt4rBnM2kvhApH8QvtOzvK464oQqZlAOZAfMHiKNt
RWRp//+1eCtMS+8+QlaQFbNc1LltEy/nWt3P14RVr71mVPR3HRBeAOCGx8S666ru
Sdn0Hllq4nfi7Xc2dqubUFv70W6E9sR/vZxJVqgk11Xti7kMzbOtAhkOV75JD/g0
nIRq4/XlKwFhCIDaA2fDPDkxT3vMmZSybZSvEnElHnD9yAcL1St96i8YeuS1m+OR
UCQunN8TfjGvZ5CqOm+uGU/TduZjzvC4YcrChT+nOnfXVJPaxigVQtl1y+YiLTBA
PSLxS1/rP9v4gMa9na9OVMQGiXj1PqRksqwxJoK85y/+QTywlH1Oa3Eq9DiqFaoN
q2sJcg8KkWxGXsJ7aTcLnX9MEdS6s54QaLA2cNtEANiL/80q1/c/QJL+4iqfnTvn
vO0xUyuFBV+cqgEhA5BRhU7GLJSw5EMTnfRDzaHg8e6geto1NcDgKBXgRGjNgvoL
OlWRvdYmptiU7RPNjJouIT136WPtVUIFShRK5+COdUp8R4JtnDmggUJGfLDKq8rV
k8OwNSrprtsnSiN/rsrH4fM4vvjJFT9CLDGgAuBBpkKYIW/X7eEdNoE3tzyi+2Cl
oy5aBCKJ3TPZ+Ncj+vFnWqKdo2lsTMDc9Ggjw8FgK+VXAXa2ih5vePfp+4dTZUE/
Zduv9tPWLbdJkU5yjfx4BsG7EDzcWuREPV8obXI8CNPipadJc6RjaKhIyN11FI0j
lDb/VAVXwtzY9We0eiWC2OIKHlEVB6+Hm5CqgnrrgjF4W2UNk2KLBIXTLudglgUx
4IdHALPWUBzigKJt0FK2Mo7vbdSZGZWtbgPGohnkANMmZ7mWByUd/sQSNoSWHt5V
L7RCz3bkfaebTdqkKeAEk2lF4ed/nM6snFLW3ms2iTan0b5BW+h643ePOoYQU20r
Xy0Pq+dbkB4z338Yhb+hsCS1WO0PzELIrJ1W/Wm4qgERM20eTeuYC0E7QhxYTZc0
UbrMbn+WGa5rREevEn2hx52nl7Kl0GoO7k9TvQ/MXLz6rqMexOo04IEuE/g9+xLK
JJiV+DHZIeJTtzXXcD7/m+lXm/MfNGgcAqA/ZoyA6hLubKXEVW5UDlG/4NHWKEdF
HjGXFMTZRMBQZTObDGPEmFKXSq3I980EjZiCxhwHmw51MVw3fq4ykqGsoLNdpkmo
KEMU27XSwkObm0QkJaqWO5rBsMsmXHj2lhHGro8IhjAXnrH5E8nKwk2iBw1Xlig3
W4958pzf2rSTLetAxIkj8HpG0PdddkQWes4KiSVd6PK1emrzOILfCkGKlwOZK5l6
eCeiLZzTCzdX1AE3ooKwWzCOvhsgFvyRb8d0UTMTVGzjBIw42YFeOcR8PQOSZOsF
UFyjf/Tz1gBqS8SkhnnPzyM3kL/pbdoOtVPvfXK3wxAtvNgjUJ63BRlSB8iq8P28
37UXENxbZ/xwR4bd/77c1+XhxMdFmSQ8x771hnEybJFxUeR/rxGdZZfRassb89dy
7unrtlqTuTmtJjdyPF628hYHc297V9J4VYFTQYvqpfI7pgCFTadH6k0TyA2nL+Hh
i53XMTQbYWRNhLGI0pNcufzuSZf2GtGYEfNb8/ByNPZzUl1pTAkQ2zsCiP0yyAoP
zdf1SWgGyTIoF3V9/5ghXDJ1ibjtoM4C7NmTqB/tGBMI6abmJsGs36HxwSU0Swyo
58ThTmAU56Q3slLF0zFXHerRdgA6DSqLG0hl2yOMeyYlMUyKz3H/h2erLb5uw6DN
kU9z0pmC9uxdeS5YNlGwdSbG1AulHhpocpo0SK3KYzXKWQNNdyZ95o6H/+gH+C2t
hnyLl26Mz+QINiGD74tnLjqzmIhG6xaKCFl/7YfFyErZyhPHGsbxUyVQ9oLZU8pg
c0e+SZ2cq6XnQq7C5ZlqcrNVWWDr7dHj2g3xCvFNCXa2RQiBFzpU5JRf1GkFUpHs
fs+Z6QDweIpy4ykZh62WMKVHwsdvo1fqj177uOAQN4gqPwkmKw+qQ8axmk5j78oi
55jF3AWgCcE4XBnapds67luCGq0IGbk8hTMnwMApKFfYynIDDtBZrcncfXVWXwsn
7UiTB3/i6D/Dkffjjy8xSdA8a4+av3vQTk4VhVelIvv37WAo0Cj1gqmDqDPFPv2s
9u3Lst6zTUqS6a8rpF98to+0Upk1q7I+FsU3ZY2+3UjpDRURB0c5SbSETCG7eXOI
g2g9OfiPiS8sdKVOrHcsY4NmIlW4CGoCpEc2EgoYuH5+PfXrlWAW27fR1XNNV8Tj
Wdns0uDUpEXpqsX8akZVcsvjJs36KiWbcuzj9BvBj4qnridHTeHHsWg6dX8tdcFn
LEMxxWJ9KPmuQO5enoqTSIz/vqNuLkd6oj+oRUm+4zjCO8LIonK7mTJKZD1Dhump
RrFTRUjNF+wq55TEcH1d5nMBHwmzgZNKLb4hK7IuMPUIC8aVZMl058CBaPci59qX
drSn4HGXTo4ThRRyj1d/nx+rnsx9Hhpk9M0n3wRM/iXL/3b1671AyjvPqLXBz75v
MO/Lswb5SjoVAB3v0QW2ihQPlk5/7r10bYSnXzKHblqzacJnsKqD/9tcpKZf/XFP
6FV6damWqq+CZewWAFrOB8mp2K+4jsYv2gvzstVxuR4bgqJkKtVg5fRhyvi9o9Hm
xeSL7KTOpOI5F7Wg+fF/2VSM7Vf8EcdE9m5wa6utRygnw1X7+bNCCPbKqWEV/ydV
1ZWHciazzqaTikE3SkadKSma1utUxZbjC8U3wr64FnhwiuxvVH36+5MZk7PjB6k6
AqiCo2YAfCK6MeEbFS1G59glbVA55nys8AezplqS74lQFNJF0tRYrmOsK7pFgrTb
q4fryfngqzHmAESweWNtvm/MINNySdOXlXqU0eP5QyeY+yEaGnajtniBKan3AQx8
NUxFC5TrrcB/xKC4FptvvZHyU8McDkkzqRdnrCoEe88PPKelrDPZA+QI74iLp5Zh
sNd7+fPyoebliAsIdKN3o+K7Oqa/rscb6md1XdQoh9TWR/Me+/A82yXogzeMlqm4
rCNEjjhaFUXcILdejZn0tnVxdDGKYhxVpk/wyTEArGjaWKEmWyqBNA1/dGwZWfMq
48wkEqZh5DaqmeCD3c6qHDnHGZxWIP1PPQe2ZIcIJ3KJoVmHPGDlcl+JycFbl56W
Lo/3/lqal0eZjjC5leOEzErdj4G3z2Rp5nSvYg/hhcr2a3Nj7uQRhNh87AoF9xWn
//24MPxL+c4Uwd6UVPB/HQLEu5FS3s59dTnv+FTNdDZXadJbDqidHUzg1dPJ0ldc
6CA5ruMapEwyOImfbhf8OuTpcqlKPnBY8zJjP/pHLAcQcvCbCSSIMt+hOfMfdwSd
PV70CNzwEOhjuWdWn0CZ5EcmHSkoM9KxSKMgBMcsQSNqKqdtgaW0GejtrkCjmO9N
zZ7mv6DZh9TGqIgqvuCwJBlhNoY0rFgMfIyHZasq8BmFrvQ/we5A0H3rRnRLUy4E
Y5/SLSZNzyIMQgvzb4lt+pvtv1h151qydnVxjlxkqlKHO2WiwYpVw2OA2bHfl8Ac
4cvZSuztQ19Zhn8S9Px+a+dbnF9zFLhgmgeAywotwWn/BWcp0M8vCUu0ep74u1hf
VRJ+eCn/IJ6KK0FzfvLJ359LctFJ+SdrO/iG4CFoCLigbcI4Woi7/OKUUjE80Bwn
8elxcn5ObFtaza63OfdZ3dV3yjTNof7pNluS5aNaLhq7tZsdrn3XWrsLvrSD9rXN
alCxa/EcHSDoPbWWbKzaqXL7i6yLfvWGSh4oXzkJnTuud6+Uk7ytm8muvuVnl9e9
gGbyXS00hIJhOrnYLNfse6Xk1dciuXDQyeNruvKau7ofnyyNt3VRWljbR53Ptjf7
p9BGOm1n50Ai34v63wreVUXg5mc7dpgXWsDVYOJoCzMcSLCagJHcYL5FBRLvhlaR
MK7za9yW5MaSrnGCc2M6lvRwmGxurwjACOygGV41U7vpM321K8hq9FD58o8mHiMw
KNNZp3jM6VPyiscs/qvgvV6kh6M6JNH7vbH6fZkreSpnfrxBtvueEDb6CCGs+tCm
jPr9FeIThWgUoPrTc4YQykpmOF9zoPNABgn8b4j7odEuqbWEMnPqBAj1fs6d4AfM
HqqxffmA2RhTQrydFEkVwkVzZdo0lhY1r1YgndO3mj0rJeLUwzNKVM/PiuG8dmBG
g3viN14SY7ej6QROnWbPkhM4bzp2rfQUhFkNsVnzJKgDYK27YOJh68p7CWirgWcK
ibfCuVMEEeFeaRGli/242LsJoVMpTco/s9LVM82c50Vr8wO5UpllG8ShbyY1hi3F
peUwH50jDc/uBX4ene8rwZdBXBxfGChNd3kw/fIe5VC2rj5R9RRnkk7BzKyWyVr8
YXkzYNt8VVHcblij/wNzKiCIGOl5tiLhIJ8KuaAD76g7gqoNtB5OpA+3iLJZ1P0l
UGiFLL+F0DLkLHLfL96vDgMQXI5zdEa0GAYNG54iUzfTG6KPHPu3z9QyWZi0fAb+
jayPCLJ432YBIeScMzeQ5rGv1L37OIFq6+sHzpeExB2DuznKnlJ2nKRqZtA6IZAB
Px3wwD4XDbF5dyMvZ/OX7K502rgHBOtjrSpSCxR5o31n9y5ly6q5GZhM1GY55rQw
jnanfbwvQN3wBYMHJnoygdBhOnfi7CPdSBOG+vMOc3IVsUl6jEt/UxUHqaZOmlaP
u6JAasdkje9EoNKmJxSxjMGH4dZkEZztz7QIuywpQsvnst8TujGCz/S/F666/LQF
ngtO+fqnkNng+DkzuhnZfXXPYnzgbeQKPdUc/dkrv3NRsy5kEg4WLxExd2t0oWix
b/hcfg+BQryJ5j+hkaDoLOrFTFkDJ+AyzPtxU4uURe77Pch91YPGCuCnIGS9tCH1
UdRayUU8dWp01uLbO4w8P5JvHf7RY9hKzy35BqIVmtrhj1egQTvv9A7zV/bdTiTI
u1EwS/SNQ8IOtg7NelvLz+ZvC+pYHp2AfJpQ9zE7jXfOPbx0S7TT7k4zILOe0IkL
Q8GhG/BsAmuLO1x8c6IUK82X77FsDbvb/PSgW/wKpbXrJInQ66CbXjQ0/i2Oiw+v
k56tgwMd+1FJskkhGrATInvi99qO7vggGvcQNRZ8kvNq8Fyr5jHI+lEiRA+DvFli
ZSt69qEQZOD3QEmrwhp5u59mOb7eub+6raY99beEdBbm0K4VoN7BrSO921VOUiIr
X7USplMk0ojJsQVEkqZums94Vhsx6BDVBMSZd0IF6aY0KzWX0rQ3RZwJhFuGZIfG
CvFdRQrwyYV+Nc/KpGA0Ex80ZTr7cfUGrLTqiDlA8gXOQCQBavo8vaWC0jPMMQ9+
7GYKi/biFW46N7cGquOHqpMl/s8+MWN/PQwR0fQofbfBnkAQuHesA4twMj1w7KHI
dtyel45HqglghjIhtVDD2b8T6ZMNkr/3INoitRKcuoAcDmBnY1dKx0Erd2mucBKW
xv2A60K5tN4JnanYoZK3M4DVPfFKl9wIuzIWGcGuTlgt+JSafiWAPv3+FQ3TDRpy
x8AmcFEYgJdDvaKED+4p2wuUx7J2PyBOEVbNIkP94vNXdNQBDnXat2A/rni9cuvc
M+9TkPFIqn12dh6kjfYuXKLJb+gH9MeBRlDIV/3MWblN9/zCz42ZYNqHDqsyQmk7
ymO0LpBIGR/E3CEUePPriXRwso7PE1b1vlWIa+oPT/6jvxMdhFvsTAQvD44r02U9
pgGds5ATgRNqUNrCqVXIJdI9DgFNyNTchcYAUBUSDn9M4enAnTzap9+QtIVeTszK
IWjgxtyiXfgiZPzQee4GuTVH4zu0+oL5SwcKO25e4xw8zoyLe2l1CpKxtZO0i0pJ
9mcKK3KC3EXRLldBzoriwrErM5+NzadfjwvBsMuv3IC9+tNoH/NktGUgb58SyuuP
fHUywjwLUKtmJDD4cJUAfbCQPZua4IatG/QJKgxgCP7WbTBoqguKVFgvvq/qltbM
yDC+oYuAf3CTcHvn9OhDot9Nw73NCKkPOvFNMedoUONj9V2xkpy+SWiLHfioClcY
JVHSW4aHJfvQDIuSS3qPnGoWIJoioOyByr+L5q2b2sFHe3cxXw0qPGQazd7e3kEg
cNX/LTBHf972ClM4cLDO5XowD4eq6tkMFBiB+AUpLObBVxEAQn28q1abErAHOe5G
BwwkgKCbtNd3QyEatPOiug6LAgl+6kYsnmyxoIh1YkxZGKDZX5jbT8T1WGQUj7AR
uvme6xq4JVd3EABPqoCAwiTH53Fk4Mgln1b3UB2K+lX8Qwxv0bWfF/0K6d2rmxuQ
XBtZ2NGbRofxXvSNjFQ1Ssc+B1Ws2txu2ZtFqfsYx94Yq4uaRJ42KTFhhD07kVr9
9Wq0UrLprHHdsGA0VTLpyqeqSxoSnzG+f/isc08GP2WnyKBGFi2SakxUreg9/y2/
0GKipJVisejU1EucJfig3yN9G7YT0mUHrCrZN5RmiSX8XG83wtDhHL2T4iYUbLx5
hp8D0Yg9ycU4DuzeCC6d+YarpPMGJiQBt4aTlGSCxkYRdKpM6byyctkrcIge/e+Z
MzXFw8yJKsUZxoQVsO2JL8M1YS3PK0/IL/bIjwG7a1D9IaHC9oRTnivTU269CRtC
BpLzcTQcYXTMIf9glmddpKMRvUpCSLJ2qmtRU+xKMp5BabPJWs7BP7fr7UhAeP6Y
+VO/m5OKlbyFDoZOerBwFgJGzNB5vUECGjA7lYoGfAHLewIPbKYL2wAPGnvN7Nhw
i3fuVDepdo17BUU8skhRuJ9GrrX+MKwR2wNokXdiHE2x4bP23r4ACD/q+QXi2kvW
PD2KL4jsoT92H14xzQXPGVbom93Z6j2iJNQXEhQVGaV5ZoAKyWMr2KO+N4rgxngN
93xEnyTABcabq+udcFho1ctaD+svOrV0RNTSyN3TdmQsBjUI0xz3L+bfcl7hvgGS
/z2lzWgKCkQWVSY56uI1xZeqQLfeK+71anC0NTKQJvcJwJtHen7cGphSAlKmkUXz
fk5G5AQCy8B9eyD8iAHAdmEg8685x2vkAXx7NrxQb+XxnrkkNM/Rddm6AYdorefl
t643mgdlNFmiwPGG13u63Pavw9OCudJrukXly635vy1+LUfDmjfSuE09MwNB2Ntq
ebkS1C5jvqhoAkoPOJO6zM73CAiLsNUlR9Pewcjbbstit9SqsrsUyBFUXucy+TO0
8u8Da45j/fBMoYwFmENtek0nzn4T2gdlGcTbHIyioJu5Wi+ZfBy96DQMuQ3dNAhi
EAormo3FSkpxxEcldGZ5uNQ7C+J0LlwLrluvAuiKMnFCZo/RrGpoeWKiebu7eQix
y2gjQ0eqve3LrKEuzEhtxJ8S8g7I/o82M1hol0ivjBEQq/1VnvOZVzeGOVL9o8I9
haJvNaxJo3u3t9EZiKum/iayxc31RDu3SptFqFd0FDfKTTwd4lOWJXMTqp93+SGi
k3lvoipU4ijYGwNxRrvWDF5FSz/HS7zY8k/PkIEVKFMU99X2NeVpcqxfr2rTq2dC
zYFd1IfgaVgNhtcZ2qjAv4YWlPXeopiRbH5kDRBds7OsKnhRLfD18lxxBIbSNvlU
JNVeabu8hjK6LRuYQCK5SNE+GVpkmGBwpekJ+qY4v9NUuN6zjFZDfCv5cOidnHAS
P+Yfcn7HJLh5RVQT+Z992dN6XDngVJZN53dZCKKUotSeQjOgIozWahqKU6v/lVJ0
oLZZIMDlJnXT2NSlo7Tf/vMS/qWTIGEpFAJA7Cc/4IBM/3UkCAtIJSKWmkjOgWyJ
c8c/CS8C/5CqrUcy1umoeY1rDJuAMAmxAA3s6b6OkfLbm6Bp5vkb2jt4PZPW7zVl
9VpacONKCEwgRI28d1Cvdr7Q9sw2YdCMacX1TRKZE5hYSsTgvclOZ1/YBTEDqmAw
JC4uUZ7jfmYUvlCibUdojTABi/s5++lWvh5ArGnGtEbo8kWio3ZIdtFd2tq81dTb
GhzGY20AryPBIKLHYrLvplZffzOukgWWQIpEYfC/GVn+1aHzNqN+6YODPSx6whJn
lBuOl74JEI98sFszwOnmL3q/BzpykE6uaEitKDOyfKEnXuNzwbcccNPpa2cOZ45l
6ZK4iD/lW3nNZVhcPecUoffP9XbPSShj3Cugp5QVw4E1mGuHm+REZCsWCtQm3Gmh
Fk9nwtBjDQwB3Onim0c0LNfDSkrinPp623ArOtTJfTptMitNET5gRex2EDAt1ARr
GjYRjS28Q/gwYdoLJPlxpcG0LC7ai4dDyRniT2iheCKy+2EhzwRDF7q3rciUc1rE
AkxWyDsjjsCqNeCSM/GbOCEC/fVlhDYX7jX06GIzSmIuzyD6MKwtSKuFdcbhqoHb
0AfRMP5p6GCxnpm626UUMm+0qltA6V4/N/IuRlkGrUcd5lkGt9S+M4EWTsvDBHHB
yU9qttzMbgPnQFKLUbaVvY8eIBhc5eyKxLQG/7f37sintms2dFWED71xWqEZCFVB
qwUPMToKdLkYmG3JvoQjwyvkqTYvK5yXZkHiZeEV52g/wa3zwaUISmnzm8Vj3air
wZtNMOsaK/sIa0Xcbyz2JfKQAoH1n5H/5zBGJO/B8c947DZE1GNKRksGE6sb1Xq9
PT/EZZazL0l6c8rn2o5u43/UH3EGJIEbxMgEwbXZll4/rzKI7XJsBBPdvtN9Yi6S
LeUdAw8eEdXRjHSScWEpNgyRNQObtLCvnkT0xSBEtbQ/Y+6rfIrRjmx05a2KDobJ
AxvoSfmoFL5DRwr1c9p8hORX0FWi0UNo8LP5QbGWW+ya+4pBiL2oInb9+1Q8opRd
vnwOVVlmnh8Cq7Jx8gK5Bhbp+NgU2YXCT8fqEKSVVt5uFNLGWsoH8FycX0xVWPHu
6tpfNJfejFHkht1s4N0nGH0pEhbCD+2UWg3S/b/LVfP9axBSN5AsLPYJQUi0jAZq
8eXBrKzlQjLXbHiUTIP229tN7+SK2RFPfPHe4peMSL7D/fvRJBjaD+uocycpYYSp
ZSuW3DCFmdtablqX6K9RjuZeupLkXjWGHAa5pekcL7Xn3sEqLRMt6Pwi6eCGBfVj
63LFnZym5+IudnXYzqIVMCeHRMyRpfUYWJDiT6epPtuL9Q2ya0ZxZn/1CbajnsWR
KBaxgePdp60Vp/K6AKA4UAXhvzHEWpiZsyvQ/qZPRJq9bXmaQaWxYqSnhjXTSiD1
G36wSvjwh7whdvcqz8L+KkZ4JuAuwQew8V8oFbOfBb01Dy7rXsn1KzwpkljS9JjL
7h9zhYc5yjXqWgtVHpWpEr3xK88WqFisGbh4ryfVf44v7GNXdY0D876eKNnfQXVY
M2fYtnCgEf6mD0mRfIqv0Qbu3+zs3X+6mGzbNdKXwNmIFV3onheA8SPW5tNrIP/G
YjAM63uoUsnRhYcW62wWiQI02+FQjfUl8U1joKgHOd+mWzn+NXFsc3+uRgXzOJhB
KO9fLR8KZtjws+N2J9N8VOTjtXraJEn5y1eHoEcxQhmKbYw1tZlLTJ8G3NqA7qnc
N5sUc/bu1jIjVGDbiojbRUE7agg5cnkPLxV4Qw052/NciGs70i4h9irjolU0ulAA
f/bpmFtlXyRu8211dSLBFcatKDoEc3eL2QplGix4f1Wlim4cXTjI9501QC43PTpu
8we/nSvzOXCscocVO03jOwdeYbV+Wog2DdumhyZnNoK4anCBQTVqYoM7FTXQriUr
Y5RzoCSkrZhRHYl8niHBSWeN8gPqDafk4Luh7y2Q+7mlfGG1UnWouIw8r5V/fPit
ogP63oQRPe0WqOkuBGMcktYPsN/FV/PbQKCxeYZuN64IPVEcva6uLzADeUCYnR7i
so9qXKICfPYPsJrtzPTn/YPsRWgaWX5claFnLINWluxKzLlxukq/rMhS61RUqZzD
MndJ7tXAwWF2bce7ol4gu036D97FHH7Y18eA1xaEcreBvurzhrsamLMmvTHRZBwJ
JjkY3hYkmdzcfVZvrcDX9fH7t58bEtXd9R5vhWuqLxEYlfLWpBzBlmQ5KGzYOvR2
c53FEz+U56u42f8B+LMd9WsgG3yUcllo1k6AkrWw0CqjUPeOu4lOBPsCRNsjacfR
8/mKE9JKh3402iht6EA1zXa3QbnqofZ4HVkIp56ce9OjCUO+XekEOS8vqh5kBk46
bZZX9D9nRXKkTp3He51mh0Yd3FCfG0YPgPogKfXWPgF15PgaPYUKujlYXEBOQ8ch
RsiVxaDTKGVb15HOyFvwTt3ceWhoCqLkHR1u8JcdcVqh2VKlo0NeTn6oCN2o0Ee6
AsF2MWjlic63/kJibFCmFcklTbX/exo+LHkQdE1KqC92yQ9GwUZd1S3aiQyRbITJ
qHq6vanQAcyVmc+41mekPltEhyAgPm9pUxsAbRn5kVnXWR89ltb2cvU8WEeEDwtY
DETqXMFbdoHGSOx7NUg32BlWvThiDYa0YuJiPXofHKmZ4tMBPp6PkJMRpeOaWqJu
2dcBUjzv2OUjLf5f2uLhO/LOSxrS2Hx4to+VKFpNC7BacKS19LeyCpP8dPXcG0BI
WWIUTmr+ijxvVt/9JuvZmTpt8ooKrrKY5bI/TUVF3AcVMa+Xy8E4c8/jZuwVbJFE
Wtm7moRi0fPbgCUIii2rNPeA0oxEZQijyH1hz9o471RT4R+wF1+4lYpqNyLG5PmS
6rZ6G5WpxlF0h9sAhO5q69dGkixXKbcBj6ynOuhtZIOvnivqX3GoalB18X+uzsts
6YEoOZuQ/JZDL+QcxBVIa5nubBOgcy0QC97ZSSU1SIOELVgxwU2ZwpbhJxPj4jmK
cf1+Glt0ovLU9LeGMZauVHRNP/HfGQzwrOJsNJUZQdM1v9/VZ5TDJzImLXm6ltrd
4oH34TpWD2fWXa/HEywdQ/siNOOSUJMMAKnWHjgN5cLdmn7EKsPtpq19sRRPEpu8
TZAzNXiHY/sdlY8jvkhzOp/RlqEsl7H5g74kCRf269wG19kLRFoJ6ZnRY1nIBH/x
6iCKStpl1hFZsA/jw1qxPXXsapjvAP+PReHIcdDKn392g0CYC9AhdrQOO0wtQPeG
3SfgenwfBSLKoXfs+eKUXuTCU72moXTSLO3zrAHsNtFvbXnbN/hzV6uTs9nnkabn
ebQL5wxPCM9fW/MF/NyeeP8jnXvlUou6fBq9H/rd5k8BRem1eNLs1yMQEwsswE0q
HnwPr1+rHoWNJt+cYIkdNqRMqc90Rhy/xWNZotTc3VhkNDsROM60EIU8MIYQHF/9
jpdmU/Yi4E6CbmyanRtgo+DLVekwQ5cHwnGhC7oBIoJ/klAQaw7YcBXUfYsF6V7p
Nw3MHKC0NKoTy2g933NOuRG0ED6romKz6T9Ggs1/QNvhQboBlSmY7/wQb0K14hiy
N6Oicas895XhVQ6VwOgS9+k0h2MT41cYXG7FCsaHGFpOBN6Xj8U4DTZYYt+Pio3p
raUNmkfGacG6DWlWRM3Sy63PYfINA5P2aeNPgsTyC7LYXLfHcOX0xgPDFDM5S8s3
UnTr7LBtkzw3wTjuFUfrhby80i0ro+miST18i6wlERXCn0OpbUmaSBa3/W+k2zbk
mgDYJpIEUZrsp0gnSg6lXwgojWvZz8kwlQXVeOodqx0LyTmLA/2VMGNNTFKfPTdB
iFuFA2PwU1W1N06bSL/R1CbWkjwGdgWedHR16YwdcMFJCJshTtvyoOiKy/yZvXFp
tIrjm3GdxCTeUzXJmT1FydWUyUP30IJ9D85oyGOldt8VvKdlx28kPJaVcLvMD14L
XWWy+jxy1IcxYjXQCKTGQY/Ko75YBYosasK3fDPAM42s9gyuOXuxgCUw0vsoDLVz
7BQli5ltkhJcwJsaNjJJtTmlb4Jh8Sy8d1YCJOm9MpRP49y6wRFClxQYgtdf0SD+
C/CYF6Uuf+nN4jJyOH4KhubOLjPKJoiLOx6EMwIKBo9Gk0nwEOqgIg7QMiIJfkv8
fwMl0lR2NByyJ8+OLM/hn2JIICVdOgkqWp4C+bz7GbhR/t3wwdeRkZnVZA0GjsLj
5gjxSvryd5uxVuZcMcqKNu3XdYkxXHgBKXqJvYn9NeiLb6BrOZkqYmqairoPlL/H
ldIgTvb8iQljrQy+GkrMbj/FBraU4oskCmnHDR3LETj6/bGwUN4f8op4pQ1oXf1w
k7kQchM9JZd4Pwt4XlRZKrhyuSpYJg0SRwCSe33D4nX52pI8ome6WAHZLZ7pO/Hl
oZoDGqpMBZ7IyADN5tifGlXu+mVzGPb/tNz81P2SaeDYxWB82c3JItcdTcG9fsZi
//4RIhbpiIplWMAwUV88iuezfUH2oKJUVBpvHWestS1IQPo+yRkQ4Nsg7Reu/zR8
Qf7lsc+m3LF1n1xDmPk6vSa8qkukTWoAN772+qeEbYsC312r70LpvMRKUrh9suzu
y/r7dzk+3M/uvsTOkGatcAGncWLSEhkRtBUFl32AeVOk2ZGfojbsBqHy2r4xIarZ
94S0EgsHJQ18AIHlsNFmjVZQTunpgC4Dw+01rSo6AkjRkBjZxjsZH2D/vKxaLdCe
e1Ege6i4mLnIc5BahvUfR4tXMdOmE6ssuDyUU0RRy2KmECOsjBxaYlYDqxN+AtNn
9zTMWzKRmkpF1z0FTC+6bHqUvnF2k4lk6iBfUmMjoyMZy8brQxOXgXofrIZJQqp3
RCSCBRQ35BlyaV+hM3ZFX3fJajj0ATUm1ftN+pskqjxmkk1qz7Pg7Fi6g8Dbpm8/
KM1QAoFynwGw7YU2QJgFA5hJZzm6n0CFNQdWI1bc6/xruF9KOLT9orfTlTCzU6fa
zK66GQ32s7n6daBogU2Pdx8t0LhlkgO3Swip4b7czV2dE/bx33SnlPvqHn1ro9VS
7cd+as7YUtyTreoms6uWz84d1ZlEYjG4ntK0NhvsXa2kA/Sdg5OVmvGYr+AEa6HN
+fknTOGsoy2prmYX9i62KDQqMZ+tnoGtADYDbShsExKP+IF6vJDgzz0LkVe54n2G
zpMQ4wEZxbSTz2dJFAaBqGm4OdaTmc4s1Q8HhXvcIVNqAQTuw+1rf8P1FQXbXmYJ
gWgKEGmosMBwmcIv7i8pr0G4GiEV1wZ/uBlIaP3xOOFMQMsSBnivQPigkj2wlWsw
SRfzVvfz/GxRbsfyWCtzQhHPaWGNdP5hNPAXaPrMg58H3nfb94nMtxuuJ5l/qWiT
EcVCl0GYafF0wx/oli4k3r+RFMqKVcUhLWi6ujo7sbCzHxcoxLRe8cKjXx1epTwJ
36eJ/VEPfec+kllcrZTihbnwOkRSzgf8tFDvdvgRtPkpl0PEUCMjsC2uuHtnjKpK
CSTPMK8D54atMABg4QSkpDjpEj3gT18KbMgNFppPL8xsSW5V/qyGEUGIXCKTrdd6
ot8aXfA9pbIuc8iFRvjOs8wVLRZVihcBLodev/1QjAn9urtGPOVivN3VgjjpLmVd
I8xlevbR88JawEw9PTMkwwrR84C+RIc4tHy8HAnxE6uuI5jAHWpUtZ5jPSJSb0o3
72vrSnKxbxkg5bgb/d1RtuQwmJFqtAyvh4heRHtMjwRqwY4OPw6tTZnH2V7RCVXO
Et4MwrcPzxKXXJAjVRrmxInoxXKlxqkyE6JUhU9+NCo8RHYsNWRA9F+VxmqlwLdA
YIc1UuMSVZ/RT9mmVrl1tWi4HtG/jwNb5EwMafYUSEu4wtExIKsqu0qldDOp2NUP
9VIieU3/+3jL6LEa5veahB+mMCVCLW9XZ09wwbzfIoJw5q2gCQyTbwMisxpRQaT5
QMQavWhSCey2hm4SUpPO0xpb9zCA8bNkWSNt+bdP2DhE1aZZjObpVcDiT9XIFsNK
y/yElDzA7GA/t7t1tBO7PN3YwDwsPeWLiDpYdNSmsG5z9HhugmBcds4qudEhPW0A
tYwUov8SSFxM+mqtSnkcOGaXUl9iWxxQquSolbqZXcexjuM5cSYxwkpxHH95ZN+X
hLOFZFQ651OQm3WVEwhfsFPbKu3M4/EjO5qK7c2rr2hzgiweqUXbYhZFSsrPb/BW
gUDeJV3c0wYHF/SpRruV1KQTd+YOb0BbFIu26EZTy4qkESYuJYDbVrWC6IRnxt08
Er4sfQL2Cse2PGun3Mmn3a6BHqF6TOxYoP0z6F712OQIXl8CO5itpN3yT4K14Q0m
LPABFZwSGYgC7cscZFQ25CzHhcnqSVB6K6t1675mpoKYdXz8j//lb98mh1TsuMur
pHd9LrIti90tzdo2EhE8QwRokCkkp9jmaQj8CddFLvWLHds9bLU8NRgxtA63VIaO
Q5cnpUkxtEJgRQhPqJS/fxArAS2r0lpbqm7gp2dK4cUQZ+03RWvTFWZSyWjj4+Q0
0RjcikEktKMCnadT69zt7OpYyR8N5wr0Qixr4ZRyqWzjjnOiZ7C5kqD8ljRDSfKV
9xq5t0ehejjK5XHpVPP6zY5bDSZXGulGnLakrvwQftLh53HcVKXaWxskKWtlPtAT
AtJ7HVwTb530TcemiQCupZTZ8nuDb6eBEnpEnOkAMTteoUEitIRMf9kPh2wY9Qs5
1WJGucKztB7LZ40rYHn4qYnDypvWaHEPkMMS7HIIp0/3LyKH6CVypssE/aFBSJX8
yOzTAjQQ14x9V/3a14AwS4K0iTu0nMU8ZUBagPUusJrTl9UuX6dTe3eKQAsYdtop
GPnIbW08MuIlAr+bua3Y1U8LBIzqyghrtXPauxjrBOv/mX9y4rZHVRFK13JFSV8e
oEdIbw248HbVB9UHLFtstxgTPLf7ZI2SEVuIs1D2A8t+jEonjID84v4cVSQsSrUY
bE6MiYCoQhxuMRGCRgBH/WoST8HmatAW76g5FDChZ6DCmRLQdwH/Gj1Sl5yia/2n
66QBjfqZOmRfi5I6gUq0s+T02fPLpOyAANxY9mO+rEVDCcY0ELCgGEc3xw4rUTSX
nUUxtpXphsIGnrirtb75IfJ2t5R8sTITC0R9+tfjYPbQmnhjp19MhmuSM/P56Ytt
i6szxsptAxEIUewj9hiK/1z57+RDlABFiuJR4aMvM2tZMolaDur4PouefloyabRA
+eJ8+7sJwXInrHHHUd0HEBiMHCdyYXL7En0ll//cgjKmm/AoPYUaGrsw5VzvQZ/P
x8rCLWYqyHW4nqyXB6YWboOe3J1Ws7r9FzXLUvlFPCMVYJR4YjYlHifEcroujnsf
Tuoz2yi7mtOpdUI5f1GvAFYW3sPePfIEx3VzEul5Fgkw83EUgPJEmE3yvOiqZV+w
wYuh3CZX+3PuE+aMVG16nsyuCup2clipnfk2UEwC7QQlE4X2SurVzqEGRhD14Hr8
/quPokgVk5CEDGGkhHRPKqmQHb6VTnL7r7cpXVZy2sO2qyNWtBmlsAN0gJky8E9w
qAR8IN1sGfRxWvUmfUQ4jCmtqLJ4sNewzUptbPb6OUjtjSZP3ZYB0X8nuutqIt9b
YJ1KXjdi8KUSeQnlRpVaebcfaHU8ckP8dQMkSL9NC0TxGEgulbgjp95TmIl6cNAR
XMoPYdRS5iMNstAM8VVjZh/kSW4s1PbQIx3AuXsLOCQLSDog0pQdZDrlVH10K621
4MzDtyQqLzIF2tCiGoMAVZ4pITxc4bF5GzXH5GfKaH7wUz92M/Z6u2U1gcS6seJl
GEn55ybD9BqaZvnrirHBmRHsv4Kh/t5hGdBCCQIVG9s82uZwLzrSQp5roWpgGWUD
FK/BHy8U89TPs5Wh8sEmeJwcE+eKyEaPNiTySXduX/ZcyH98jxQ074UrhSnRM0rH
NaGezucBvnNIrJOMuiM4imuJtPSwChJJqSf+Mp/xvrTytAVL+NHwhMHOAyyK5hLv
BpYz4tvqX+haWLUngFDsQDApYw7xorB1RTBSozjDtxoF6XTkJiReDidKDMX0Hokw
5VrQ0knpjp7Y5y/3mMcnv0N8UJ6zNcQRBwF/y1Gxwrd80lMn2gCMpSe0/8WalQIO
eHpRtxjXy5RVtx/3RMBu6iHT+UviFp1nIImM+FxwAquJzLPRn0LkZuxcZf18bLnd
lFF5bt8N/QsxXXR8E6n3uZ55/gSYQ5+IsZL9e3nAHPTDJpOB5Y4g5n7WMSMsIsve
6fd/QrvJw1tKlCT4dUKBRIwhwps/vByiqkFUv8cKXNdOijkKCYpyM+TlqNYub+Rv
RfOsY+B+xGkLMpIvseDf39Uu2cY/AKuRe5juJAWLNEQTV0prJOhrUX+P1cNGhBzR
WuYsNiImZqncRN93YpPWSj3SCWAKtxGIgvYBDy3DkxxTStDJX9pFgahXoBYbXLL3
ZLLDBvnpiHDa/b6VH7e1bkRXmc7rsNdqURwFljjqpuu23nIcTy0LhPn381nHwB/R
wYPesIrpoCarSlnDI/K5dbwu3UKrxZZGxlBad3bsrucGxceWTts3iBbArPCSOdyU
pP9+AvMWoUx9WjwdxFDOKgENKoFA/dh9XX5Nn6mgDCyJWqtZrgvNIK8MBbQ5SOt+
nKBPqVNf7CxPup/PjJpTumyM2qT8zvbqG+kgO4kA70gMZI5NuGDzpZvmJpQ7/chV
v9QuWVSeXbkkFmXIvA1p9mA8Gx/pcQVAXLdT6TYpttjrybdxyErIrQnRk2gVaixt
zcvKZaOcH0Y1UUPUq7YhyZdrj2zEuGWF9lDenYPf/eNu9bmS0R5eHk16GPk4y9Eh
kpwh/9HUHZwlhAAvyIIBr/RHgZ9GugIoPNvaDbTmTuTUGZKvlVnp7OlHW0039tJi
pCq305i/Ailu7e5EjYAxhRwDZIHVbzgXbOz3Bbez/E8Pxe9M3ZSkqsGjFyh3r/x1
XV4CMl4AWQII6DDmkqysQj2zml0JDBMzoqZe7I6qrKUSSdyyO78NyNESLwRuo7uA
VnAmoOXTdESfYG/llyA+fAFhqzfgOphIOivNexWwZzA7Sq+i0sRKA2zlsPJTTvYX
Z8mcU103Alkz5JYzHCoCZRpPwvVCqmd0cTO8OvrRfLY5rykbNMEkCzE187wW+S72
48MnYpCXknsBazr4vDyWtdIke/tXEVO0n1kpx9rA6Z4bmIOApE9WbdSTOCvnfBAO
1ks/7a9RFlG6zXE5ragIM3kGJB6zUmcIUsQmR3FcoGVqxXeTKb+Wrui+x6P+3F3S
8JJXnvNZ8unoHPqX1la/G5qd48SxPAPOsL6h3nBcnOXh0wMJoo94rxD5SyWmKSH9
Ud3/idQEfDjkwIN4zX7S17JB2AJFhqw1eNtzpdpyx1FIISFrQ9paXkJgdl0lJ5oE
qqO+08rA3X9VfNILg6TMM5p8Zf+CngaDnUV36L3rO2ElkAMkmImWDJm7JA6HNK9m
hctZnYVuG/fBiqMMg5K8PbxMfjkobQaf2dnRhlkfMmT9bR/6ebox987JLNIdkQjd
eq/50NViVMTmFm6okr8FEcbmFxw3rhkx8gk7ti+7ffSoVoiy+/eUx1nPm8orX8re
0gXYLFDuojRmmM1baDliHRLn2AAMUglTTkpA6gg+Tx5SLZjVUb3cFcL8UCX262FB
FHdxG9M2VESf+15eZO4iuPLmNtKIUGsdVsec/Dbd5Fxtr9qJkmK1jEO0yt7iSi14
l1Gr4fmPfICVjfiWlM3uWnS8fn3BfbU56a6svX+wr4CCKKIUDSXah+u79QydXUdZ
cUZo+YCPEkEfONKgpmD6p/EiskEqTrnFrIjyKJjAksS8AO/TCVkMlZQhpvLpULZc
vXGclW8Q75rw8Bfk46kwBQWKhDk0Bvl5E22BCV50Gmwc9GahOjDOJAHG9An7cB0O
JJurQlleMgaN+NzinlbYMQBvPSuihrcBnMbyhBuhUserpD2FKFZL9OF7gBqGVn2T
HqH63qTikqpBB5sSyNcl35s9E3sJdTQ8lporrSMRH2HbTQsCXOO5A7wzDW/Epe/g
qcnXZzpBfuAGk+L63sFHOzfcQJDW2jZMZpBaBO89/H5KrFysf27714HwQ03ISrAn
7dl2ukG8jJt8XSU57wtpADh8BxzkjGvW+45rVBVIVZSFYdg5q93w7cY2kKXOkITz
pluYP26bGhkmLgYdCwml/ssojIkYr1Ma8qF24hQhf9D3W9K0dBWcqLbwtLko/TXv
rb0yOWqih/bkmiZ44SZmnbH/AP3H9uJg2HZ1h9e1MJ/S0zGE6YBKAwMi1GDbrrZt
JeK22ioJmpIOhlfQDmUhzciKBJexyrd3A1D07FFIZ6QrVg2QtTLMqlof4/ypO8m1
wq98Y1OPfvSM6kUlnBk1TWWlcKg1dEMnSPrE54R39RL2agUk2qD+f8EEtFTxdqAv
pg/RXHgoQAxjKHVcn40rVxbfCFnTXv4AGWuW9VyWWzHeLVGnh5YnmeNEZYJxujLS
CufH6f86+isAAWoFayhEovajGpVPbY7h60RKvHSje6tP7dudrfjBBdO+1KPHiKA6
k8Ap0oUDxKN4Cf4q/dI2dn7n74Vb384FBgxaxvaJan6gS1gg4ONc42ap68wANfN+
svlu3ffb+hGf4cdfIj7Hr+X1AZnoI7uuQWfdzoAMK8yd5jLkwVWwaHAtw5Fub/wd
zihP23S4BmyZ320hpC/mgBPuaTvQ5O6a6bk8xe7sekilFifir6nuiTxFrzMiMZPZ
2S4Bg7iIRIMDvPiNta2U2dH9WMXL38dP59P8Qwltm3omftU0nh5MjxQgUoA1WIfW
OimjtdFfFWxAAoW2sgCye414w5I1ZUX1GDVFKVvDBHD3lVz45a+Oce6HXs1un+xY
BiGNfExSxoAD1rmayz8TuWOEr2iCjEtqjObEsVdtD7cCA5qWtVsB+hwcwiXcqw/n
dNSIOF9Ln8V8lvZim2kLvgewvxEp9F1Ps7SRRmMPCk/rbph5zCfiu5zaaofa+npE
iSTmsWaEzhOEC+6q8IDKa1blWf/ZtyEoKznusnvQ6N8lErSOIKRFu3iGQSylpsm8
Ku1yNplsstQOb57wyfuaO2gQDLPFPqlh8cklGqFSczesx8HPy4/UGvpaNHGNEJSX
nYsASQRn3Kq89CvUiry9ZY86ykvAwsa8whdVldLuC9NBInKYL5lcYM4n/d9okpzQ
uBbrXld8Ez6p7kj9KoGloNMhimWbRnEBRJHDtbfg5ZNMqBKO61856gPqm5i7k0oV
FVD9j9j3JitjvYYKh86vwCGT99euh9XxGwbK4+xeu6vsnkMgaig5KtV7Sx+tRaHg
yET9NodE83eG48by7OwzLNbZLi5S36CvE8sRRWwZHfcaNINcoIeY9hGtvbVPXtp7
HK7iFWWlkZ183O1KLsBeZRdZpdscupwBQIuAEitfxf0qjAOGfr+oOLEp1j9o+9sG
NLnOsUiA7bnUOlej2g28AsazdfC58HaH331Wd3tnZrbrkDOhr6SWL7UvCOTgxGI4
`protect END_PROTECTED
