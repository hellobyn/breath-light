`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1ZwX+fRArMFqSZM4O3gmtmlwDaaos0dssrhkdcqI0iSjDmVLAIWtzkTyDdeXNSY
60X7XUJqzjYn7bYFCYEtNavuacrZkOxt5Q3yCCPMQJTCfPx/BN9pW/cRtIRreWta
ox1pQNfFZJI90yMW2nAEglw8KceprBdgvR5GHDsKOV9ApIJxwyCDWhc6w47j3k9R
lCFwcoQLAkEehc67TloOauHsGzwLtNMAB6TUwWDGnZpo3w5lUm3XF4jIZhpz5rWQ
LTANipw1Fz+BPJj0EFn3YxgN0wvPdPr/5cvHYMYNK5imTWX8lD8UrBTtLxprNUGA
SGtiU7IUmJaZsJ6T0EK4cGLDgHwi30UWBWbx7rNP9O0wHwyBxiPerHiMtvDVyM8b
AFZz9XPaROgyzNeS0iuhVisfdtqXiM3xK21g6r+3NLtAWHVmiIlwfB8Zt8v+OJ2/
kjkumshYgj6bW3mS+5PXyj85brWyl8RVaNBMTFI4qoclEeEDnqIqsqrotOx549XT
NCryz0K51oMHloJ/mTSrA5dD6bTAMPHHdQ2oySB7YKa4FpxS5IaOVxVzuCTn60wE
4E5/QIqdyIJl1PmIJ12KXcNi++KvJtuNHgrRZf4pXVwui/FanccKpD1u2Yb7SMyB
47EyGmnE6uc5uMdznVztmctNQ/djHWi3+TLrdcfla9STgamR5cTMFh8OWbotba//
Yha6sXMyB34z9wTEPcvaXlkvCZFCz0pikRBonNC2prwYvD3fk406lbX2mS9CXNik
10OCbOZjWU5QVQzrmSjZstdHLkJfTK7xWn77TXsqWl6AbFhh5UGqtKO9HhkS16ur
2Qn6JxnLRWAnTTtuZGS5iWZtIF9lCRH1RZtAMSIWsXlGLsKCtLl4leyxGXmDOlgB
i2rh03mghsciAnTMAfew1pYbN+fG6J9RBb56WFerAFD1DYcDDeDJ8FVZsVOEi/j6
WdEvKf7+5dehMDh301m2PED6LOon9OPLC/I55pVBLge2et2z+bLqr65YGEmUj5C4
SiK9/CkDDlYUr6FKJjqE7b5FFbxrIXEv2suOMS9ZmqInaTmERRcIQSiEoR/GuH14
aN3k7R24ANXjmymmtzzHdaY7Q4T29L0PGkG5cX6I1f+ZeGOPW35zqXV7LC1Ehqdw
RLT2prumfAleCUsvnF54Vo9WU73PWvjdUvODhw+T12hpB1E9dY+Kc/Q9+jviwr/e
QsMRyIIk36FHA187ikEoEge8zB3ClOndHqRIUzUlZl7Jkn7OJjsCZU3Btm/J0wE6
+VNKKYN9gi/KBf8sSuiBhiliyfdWvYrJYL/83ISuhMNvboKm6yd6A+aAG3ucxveC
gvMF7J1LHhKorEfDecxhjoEZkNhvcqFnQpQDY4FRnBsx4wta2Hj/JyX39MJqjusv
bklYYiyqCzo5cvqVTFitCwwmAb+R1zk6aPq9hqZSyrCeD5whP4PqL6M12rJL4yve
+oi/PhLSctInWsPCKxLaU/KclFbNhqDMQhlMZTuGhhgj/6LlgzKIlCZgpbc0iSmg
kt0Lpi8idApURqAZSN5Rx6dMgkTKvTWlRsDis94+Rsczbow8eOHulyiOnSw5Aa9M
WJllACxYeVxtrrXAEQgKrsX1JAdhrNGqdOfenqrs8Bu+NF3iJ/FAyF6GfuFt5dHL
VSK7AakOs/OqTzQMULxnw/Smpy3pfZXqPOwG7uEc9oIf4NvgObWP0k9m/66uQZFy
J5NJU4lO0R5a29g7fBHyJFUJNOnN6Jl+SaMegroXYqaTHH97zr9N6FbiG8+G23Be
6APcLA2OFwN5I/QslqekwEIauSXwAEjp0GunI8SpkBgXANN6xUSBTvcmPOF6xEnB
7vM4Ge/i7lww7/ZWoM73XDpCwLOc2W5xkgu/eLgYEOYXd+qcrdiQeKR8FCpnJj4P
xk/M57qQ4b95evaRWkT6bzgyAsdGg6FvJsFZMUNCE3FVMOFxGRI3ccuZbDLuuebR
Xi8MaMnXitaIj9GQ4D37T22ZLHEIkefnlG5rNYlCDhJJPiSRj+9FBJNqR1ZfVFrA
FzAjbK9C8Z3ADy8+ixYMvZjyhSkMaRGbflZRBATDLE4Ld/22Shv084CXSU+H/kur
Dz3Ufduois2/120HvA0MZpaalPj1tsSLBg34TQ+BoIkJfwbqjQFYVpvi89Sx9/wc
l83kAVb9sVPnaGPNMt5Tjc9fPtnKUXtvYpf/dUlTIDvucPSYA55ANWUx7J8BB2LX
QyyYXqznvyQ/zkTth4ZYzqrKZw+3f9tTjRAOU3yQuGh1Ud7c68U0Rsvx1rUKo76q
fwIeQSRWJZdI7UgE0Y1r147q1ikHw3MzVPPsQ9ijPU1pIeBJMTOUsOLc8gzRLFve
GCM+vc88UFjuYUb0EkH6he+UA6mCMsKAJUnp23XUuhge+c9ozXgit3z++FM4UEiC
VQ/9S2Esw/PdHaUQkVVS7YCZpDAA9sDH7XaPF3rN2XIKsUUPLKkSWt4nlhKlcRdi
hwPgf09JQ/XBNSXNm5xpc6MTMwSdgZUUb37r+zcQwbBhIppGhdtAbeD1mzjpWcRV
UEPW4i+7dX7rx4+X0lPlayOUEoWkxaK9srYagil3Zi2N8GCU3LJ9BPFJWt58ibgB
D/u01xKTc6WZ6iCn2HPQF9nx2b6pMK7kt8xbkg6kGYU+ZM70nKVBCDUxLiNHIwli
eJJCJrlmlMrtcsk1VsJfThGOuMHvwxbr65rNIwIEBzS5AWIW2orFGGkWmDTMcCw/
`protect END_PROTECTED
