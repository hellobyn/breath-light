`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVC/RiKtQLspW03LKgcKGjFYI6c0t0/xwy87355/QKkygKPuoKEuIV0QhhVfzAnW
aUetRArP6MjQfBvgLutSF7epKRlEmoQkilDWXV7A+eGeFtUKj3cMNTp5F8igfCOA
NF3wnfqW5Ap2Fzfyti/DCvVkWRPwDhn53rFjcSkHI70s7m6XfI64nYhP61A3MOVY
EGl4iOzynGk/26iRpnepVTK6Tdu7us75u3m0a7Rng9rcSfA/1+febPLeoWm80CIC
uRstdIIzdNZptRViELoXFniHgwE52XzjqWcmwhRGVG1wF6FTDam+exdCTEYO/REj
NXGh/8PVN3jiMDymYnIULOid2M/ldabqW75jBjKFP25mpo10JXdEQ2MOBg+97K+J
6ysOGSWVZAVYyLOE30o5zy4sGfV6QNArmhBy4r1i2M9d8fivIFCLwDiZ6qT+S1LU
t3RjbJQ4GPQyIl12kKL7AbwhhKjHscpUpKhMV3S2urqooPypButLt4xwtzuRNqQB
tI/iS6CPil60MRoXJFn8dGifui6xZ8ene4CHZI3Emva7dnFFpBTxq0Q4hpjGrvKZ
lP9jydgLtavyvK+hAAnkyzyxA2fug1dCNG2WUEfzldfASBKuupJdcYjzv++x4MVo
toHWnjGLP4/Zze7eGxhVmLcva+qT1L5PITprOXfJ+WCRkBiymbhcsFpMMrLtAGBk
Du37cH6YayhCFMcbCMJ9usGAnAax3sCtsSf8mzwuWzd9y3oAQDwL6UExIYHhrIbY
nYwivSAis9DtqnUy/s/b6hLN3K6ELeQUPzQ0soOi02qRPvBi4TgyyuAO3bEys1f7
Z8C2Kfw7ZCQdWKcS3m9OkPLyQ77HFMYWCB6kbeSWxnY/K80/nerVnOz2o7GRfFSj
CkObqsFwfcGedv68S4A4fJBVQwbj7LyAcwRsn3gr2zDV/N3RvweOcvqygxLxLDjY
mMV1IyDMkbk4E+0AIzr++cPvVTruHeVgjyM5qyZFPt8HGh8jmpME8bcCs6JDo4OS
KjwMjcmt3uudX/cjD9Ghrb0l0oHHpckVvQXGaytseCyrGBVZdSXpmvN8V1m2FQ6C
iuBP7PWKtBBtChB41HFcBoi2i64ATSNNZHCI2xcHemoRX9raKN6KYtvfn/SIlcOt
yKayBxDG0RqGNZQsmjOkZ8dfQmQiHx45v9gi80yKUets3iu6cQdVFRZRf9D6vqyb
Zvl03957pFYoYFmtkliwKwKCLdSScW/Pmfxe0FD+HKOBf/F/6KY8I4TG2j+7RZPa
nccwR+LlPobAr1Wl+6Bug2t7ZuZT2r9CYBGCu92+wtvDCBSzCzBZWnJcPUfubvky
FugGfqVMXRz9Cb2Tk82AL7LjvF3JPST4hFQrlOdatFnCyeGHQ/IS0ZUeREkC+nXC
RBRF9V51YnMYVGBZiYmheAuoP6xBVAuLsh7cZYd/8ydIgri0nCKr1Oc3lOWKPBbS
G14j82OVWUlq1c1d60ncUK6Nf1I4ujWLhCcqONYnc+h0WFg2fXJR4l27g5VnF4dQ
Zo/Tmhh2hVgAILGuU5KMjBJ9rNNYZTbMsbuPld4zVsfkTOignoaP5f0ypWiO74uJ
9huBvKJgkKDZeHnoQE3o/plBU7cpvl+n9CV8KB0IcBq+rP1J/fD1gdjonNED89qZ
+BjLIW0AB4TDEUb27RyMAElihldFMFO+qd7r2M3y/FqynEsIkxP3L5KuzToMtibA
94KMInbop7p9z0euM7jWpfdGpbVqKGmY1IjuBjfBbQGn3drg6o5hLP6GVo/6TO+1
abcZRzrnsqKOp7kQjkbNIoGJIJ5uyyQqJOOwXOv6cPAv0L81SmpM31KIId7ioa9B
efIOiRpyyNP6+3fp/BnkDM5Yb4ar+HLXnHJUbF0e+eg7pylhwtLXPDuFJ7xlXy0t
yZdE2VRBC6Pmu58EF+vh3owOOI4jcawMoZbbpL0UbMjy+iJ3Su6Yyi/7letFRFqC
TfbQBLr0MTLRMKYUExxGk95CHAQiBLG0LRgNrNfK2PT/FQhuDDC0OesMhvV1R7/1
S95eDZy7OcbvD0v+gdOjdp8PLh625k1vW99T2CPftbm4VsVeIK6+dFUrFIFWqtaL
W3Uyf1l9qs5sEhcAhoZxvWC80pl+qbCKXlnZsP/koOx+H1YDTcp3jpfLEg1hz182
A5zxLvDtCf5nzNVlin6v2SDqfoSkPZZUQAFZKlgOZgKp9m33gAOlXl9ukIbi/fK/
KuUJIoo7N5UspMF/XKoiapyV1U6oVt/4huCx2XzVx59mIZxzoKmu/OkeqcefNdOp
TgNkAdc53/SaY+naVktPmwvxdEn+PJmNT+UxLfXEUumRZC8yCDuqA1ZPf6ILhbij
tNpymN9ED9FJTOsvx6LJ5Alk5vHDdtrbMXEBL+UOKE11/oa7zcK2hRhu2imAH9YV
Jb/aRwcoP3DnwglKSdLWE+3ewoSjFwEkTstvnwEADx3OKjqk8d4adwTwpOsoa/Uu
VuPN/E4OPg95MzrofRr+rw==
`protect END_PROTECTED
