`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCa/fAIQDbPd2lCApAkrBWgLxGWDRxlv46xuWwNugQfPpmb8WiungzFhC2CCaIFn
Ri7uaSoCta0gCLthxrjxcUYZlKt1PCXOkH1FQIGmplzv9jFWSKmo/BHNOwyPfoM1
VYWi4ODEXRVeX/u5CxB6Q+VHNIjIjKZNdLuN40Xfe5Glhy6xwqmbATBbv9FH9Wt5
/h4EeoeekNmEI+RTwn+3V9oU4p9MZZ6Iy49eYgxh1hcSuvLX5zt8NPnVd7OeQUIf
O9m073K01YuC86iQiNeHxdOLw6bpLHNceDiLST22pu7YbKWoVnyFpTzrPot3SjKt
VRIIT5LwUKa+6z+QY6yOQwXbPrUMIcBPU/SPJqdj1iQ3qZHq1XXZVYxu4wWu62Ri
4nE+E8o6Gi5s5IZVpH8UyFEuzjG69kBFfpZt4WU8TfdTXac+fPcySFT7QDWniAUT
afyyhfggJSILzzAl2Yor496sKoreU2KYoD/SMsICmvEap26Wo9/w10JYi56J9vqk
DyFu63m8g08Zu1Bh58zEf4jXtqXiQuNZEfQA5WtYUS+5RtHNQSYYSi54/ZwRMyfc
7uulLWY+xex14wvrRe3scM73VYXA/yEgyf7xdWjUbncREZCTjNWUVURagSJyQR5A
YthY9eBwg9KAgiMGhPliA65Ny/Rch3MVBqFU4/5FHjoHytt9EnPZJdO672HbIZRP
PMV/Th+1kZsjKiUy2JUlAbF76D0XaD8TDFDd9nP1ch4yyIw4Lx1gh5aPm3vAFcxs
iNQpWvQxQ5PdpCEMsMSHuhrA+E6uZVJY0iIkcF4ScLWfXZgvHgV9ZmD0BVjDnU3I
xW6maGcrtGr+Cz4VB3ZSU9y0r1OJMrY4Ql+0CIMl/2s1+m6bly+krzi6jqvV6S+n
xotMVvoz7kWWIQdrERQQqLi1ESWoJ7NfMOBXPx9JPhbZZAf1Fhk+lhDRAa46Sb+6
YSt5pvFGLjGEzNsjm62g+gcPeI3XQSgIwTJ/SUISYUqKYdYvMCYzq3n8MXNTBkYf
62yBWwaWzdNLtbdD1l+VWpdfAEhx/4vvP+NKHDSKFcIAXmoqzRCSdoHcfnRA9CDe
QZ09sXPcJecjAJFuuSrMHP2ZmGE5xUWa/L8wDPX8UbALHS0vLOWOiC7vy2wj5yww
iYy+29LC1/y5rZ9YMOmG3+HxiYSCdIrePfz/Vd5XsKYDuqLeI+aCR25oiixlLmmx
RsE/VsjCWcwF6QlXkg6CIUG9zvejnQ4rZewUuaEm9DGrZr7RkK2UysjWtjYZY0BQ
CeWlOpN942axo16O/LnREOw9hb/XSCEXB6Tihqj13i0=
`protect END_PROTECTED
