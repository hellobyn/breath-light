`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQPg+Hs/2aXweyAslO6RppKz3nWbl8i8BerE6rqD7WV9J0Slmk1v9wRIxBN1c1Ls
06pvfaM/sJ1GpqE3MX3iVMGGfb9gd15hsuXa19Ej6QXl9bbVIh8YrfWN5qLhYEQ5
LeVkMA4CSAW/aFAiKOS6iGu1e18SaCHvTFlR8tMe2OxwEGREmuelxneMEPGjIaDo
gF9st+mPuK976LqcHbK1pbo03DItcMUuacym7WQvbkPO7tQBpo71fCEiLauT+bU2
XuFSiEXVBXltcUazFfPUXDuFRO1ZKHjbuUxOYmEab0MKiNXZt7P5649MEzvuGVdR
IfJQV2qwea9P1xeYElgLa+Fs9E2udTXDaE/QAHoCEH1JQrVhU00IekpzFg3baxWH
UL6mZQiCmwYYucjjqG2Hgyk2VQf1HgkUQAU0+WRvPZTVKWeluwvsZB6xcdYyBsX8
MKMfvd5TSelrQkfgCH059huqB9ANHM261nVICuUEkpkfbBfVUq11Kto1HyHYMRvF
bkWqMDxn3Rg7gpSPXAXuXDR5adXfjWhKtc1UAo7I3FUHtjb8oF9yaJx2E4NV5KBw
GKxL/UotYNqvAiv59VuWgDg62RaceDUbcnI1mNppGtYBTNa4qjPDedszT+KNwUrb
oEkTx5G0RfBNkAfSxQUfVGiyO7dK2CgrucenVV6jc81jHvnVYMUzwhMUi7Fezfnm
tbArlSKMc7mWm6slG9UYiGkPJZi6w7RkNQhp7VbkLAoFxRU/bBadU6ZyJjDm8brr
ciFgjiIXsS8OqkAMI6GpC8ofaFKDPhQGupzY3VGFQIRVmyET4urIT4QCdwTeIflA
HrJZOiFJANxQfQgkzqd8Zgur6lKHqGzPz66PnBcFt/rF4o9VUaJEh9rzyFY4z6bQ
JRersms6b+MVX4fCEotu2TLK3/VniQE9wzi3/npAKa5M8iiL9mqKmSfH1R8ew/dz
I4E5r93pgYMVHSl/Qq1jZRsQkgpPHrnvXoR2je5fYJmEEFVDRyrJpxnsMClCp+9l
yxlJuebYk+wwGOKWl2m9ryIHRvkwOrLUN4MXHKR865nvateHj6JjErgVh/xWzbcJ
dYf8tloY537rpYQCPkGN36A9Xo+9a/2YHWX409BD2eSefG9LkPB3VxM6ai8Gy16n
hTY7Sxvec/qvCbhs5YXyawSnTG6R8zPGIROjyDf82+4wVh/5HFiHeQFQRVc0Vuub
L0dYUNBv4LAP8EBZ4zEfwRJDvVcKY8wD1MiIHWttX1iXJRb8Qqjbvzf5s+BStbgp
R4j8shqZydzQoxmhg1dT8ttVLkApxZErEy3ZgALG97ceOg20RqHT+KvVT8ZqcXeZ
6V9JdR/dCQ0LFD7NehK0pIoR3YmZNxcsgSdj1CIsWDH7SAtiq+HoaAajeHhRpkeR
TmUOCL4q8/VUEJKpmvQjbySFQJlS7VtnKcApsXkpIp4g4m5WTB1mYvsklRICUWPZ
xYN61LTiUfPY73X3JPz8MqKBWVPdwpVoGj2YpYjxlhMDif62fbbYQClFF5lLfQAf
fjeyCnfyDLz4f1Rmhpmhqpj1TNXiZCIH0vNPQDgwahSDcWdYtBBSHCMnhCpsDC3t
6rxS/XQDp80naeW/RSUWmqWWKoq0qdxXo2RTp5s/TuFDu/pw1T5U1ODVGcmTsLLI
CqFvAmqWmrZ2+M/450IWA9wCHUhj/iNuvXSI8MRUZe+sq/c3O640YGW7U7tpMVbU
sApXuR0164ETFF5IZ/kakfF0oInszeuT3/JmM6KCqOaVcrqt31rJLQwEFIFyAiJ6
1idKG9v4l7rDbUI3OE4EcEqGQ60Zao1wdbZRvbmAJ5q1kqbfz7kbVDWE2+yCLuW2
xbP4XZdCrGBZ6v1yO0kS8jL1TTHg1MgnF71vzGA9iLlyRCMnvZkp+M3SJkN30EKg
FldRjxDmka79PXUo8+taLUVxVeud+r7AwdjBOxEHaaetqlj5HmAW9nmlHnyneTmX
klsnOf70CWTo0TiuecdHkKfwKghWTFxSeu+fDPLgXNh/3J2hdLaZKdM/Eqw0ikb7
NPGlolavgewMf9yLorH6EGFqh4Jvkl+NrMmw3sxVAogfmrCLoTo87QS34aPoT+Q+
dH6jSSHS+avmnsy499sqKeE++IDrHYB+62IsJYE37PrZTwPIpYaw9U35fGlEbDPw
5HkSL3WMVtL+9iKCw25TVDGYRhizjhr/k3nI5pqCK3ATbunzptuJAeFhmiCNDdhJ
p5Z7fSU1vaG9HTsJv3z6lQIDWZ76UeTTBadjmqW4zHIw86+nvmHrE4Smu3rnIV5H
pPDHCAB8ioIkNk5RZmJTFocvPZSUSe48jCQzDAz5nOJ5nY31XMQIafDXgrLUdCnt
fSug58zB0LpQr3oBpiFhqnyDUdymaAq7/f+xkjnU7R8eeR76KX71FFh273j/IxPi
zPfAYP+NYPYadWJWMWVODRN4Lf5xOPCDpaOWgaXNlY+zAl4mQaS4brA03w6XiVo8
EJkgqn9avfVkhj71GehGrh7SvWI9ZP5wmueILVmVH9NvCBK9FdeISCS94/6FHIAr
qr7paclkrVzckwaT6Gg3HY8L9ALjEG3HqDI0MwNjmc1SVWZCQsHz5CJRuMhlQyv1
1BOBrpHZHPKQ7cRoUNkCmVKChWQAJHKhs0CxI5+ARMYqoAHFZq74VO6D1I/yljqs
42fl2Y258fBDH35KhDQILkVpW//SrbTgp/4cuQBKoQ2Bm/Rzdda6G7FY2o2QJNe0
lLRUkl8qQMe0BVdFBCUQRduwFR3kd4FNdZxy3TsBh6IgmXFt1hPev8Z85lFXpyAD
G6C10Qwk38ohsg52D+LRynVL5hKcQsnT2/x12cDjKv0=
`protect END_PROTECTED
