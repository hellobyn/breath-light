`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhGITLMZww3isaiSSgC5sQJfjkAUPTbG/17dGbM7seCSAzL+oM7ailkxAROOWbr3
KBt/Tm3+3JyFIMkNNYDB/DJB0FgoU7z8JzbSU0ucqH39uMdARGksHWf7a+orU9lu
lbBDoUwKxe6ljI8MnJaAjh1lezE/kO4qhnZtr+VOMSLoIVF2k2oP8XBcR1Ftsjei
SOk3c3QBlEjqDxZUUtmKzw==
`protect END_PROTECTED
