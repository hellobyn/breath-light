`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3CX0FwzJBvd/JhUXd6WuOpk1tVzC6MEULQiT6lxDp9sXgOM7py7pzWLJTBnH8Ym
Re/CvlD8q9yo4w6fsj7+Wh8XqO4GdP4ZzslDj+bKtUWW5eK/oktsBOyJxyjwbGls
rlQ5NMUJnahaiaj28LK53//COSccbmxsBg9ul7+SueYpUjlwyQn4qXEazk1ywX0F
y3l/k2P+N3U0/M/M9StbD46qvGgWq9bihjEK7I5K2/rThXE6P/wMHSfVqF429J3Y
3AbSpKAVjFADgj0g9MlILHGw6oGX6yWcAHF2WahNWmz8vJt8QzyHtcZYUXst/FnQ
HenWwfTCLC/wtIx0dpkeNvP63ExYFK2+nLsh+pHNkSHQTUOc4znVa/opUSRnBboH
dCYT4M9hdEFUxNJkSnMvUC0Z5jPLIRUScwd3pC7k8oD7DeQFxwlFaNHCvPhsJNuI
vJ3LmAiiHovJOPMz/5eRvpdbY5ibWiWB2NcgCuWEKj17gugfKoHTfMuRPO3leai0
Thm4m1InkvzEeaIBDYJbq/Cxktp25Gcyg/gl+4kEaftWeOU81wG3PMiMWMolY8vF
fsck6iRE1M3kGAFysTpNxUi0jx2zIYvSAFr5PNeGGmXFp0T8fqK28hBmQhj53Bn5
xLqimEbE+HzfN/afdzg402rxgGIM3Nu9ywM5at1wcDHBtuCJjWwMKqAQi+pxv+ph
Hr9/XPVnNYeENdVzW/iDB4dRQsFaRrrTIURav76veKcauHxOSvRCmCiJ83bKKU8I
hEGry2D5x8BMxLetEQeK+AfudhFzmQDTd08wZe3sAGE0JtVZ00gTakHTVbTk1AgV
CMNwWvBJzhO8Sh50qbw9VF9ihauTNM7q7V/cEKfruzFo6D1KXKE1XqFaPVBHD5pa
9srjWTOrdFYN2JVOd9wI/LEXOcEF9ZtEoWV/XQB9UClzhV+NamDAcBOIfco9z3k7
f2hEB7F5UwvhlGLVV3aGjqtKJiZES3+g+T/yuDhzzVje7GrwR80i76RemGVC4H3/
TQkw5/Ls5WTuESaMGYlRk+fJhR2JQMeyh3lnsa0kaUGgUUNGv3JpcNaq3He2l4hu
WxpJW9xEt8zDPDVLQHGp11q8S4mMogKNAMvkLjeRlzfO/zEn8Z3p9Ef1ATtKsoQB
llIup2DOQIya+/wj3Np3b8fIWaUn+uMC1Q+4UjQEL9hXd27axG1VCaS6i0Od4eIC
sP427hvoYsVIX6g+gsgKdl8l0UcrWOZjiDViq0sLvMim25oQiWw1IwA8bBbru97U
Bo++v9ZDMqhJmAQeTJ3vQx/g12s1Knh9rBLBOGpMQf5t89t+6AxYesA/aZfgrv57
Dgsi++R3vQ/7q7ezAzMxNZ7YrOJqAZ2Q3lsAPLdKJDeoInkSpGTFv4zz9lgcVHaY
g9GQdIGfuZGqO5fPPCCfolWIy/TQCaOjQhSS95yyaGF1AcpnK6zPIbaifZd67tYY
L9Qx/nJkb4LgtvO6GdvAXdv4l3GA7u2cLxwmNpt0PYI9mI5VIg5o231yy9Y4qtkg
54RR75fRJQumgRNTRcR5x2q0Ai7olw/qrihMfr/XXGeWlD9iYcGQ5PRCvSqWuNHQ
FL8PzVOEBppVoKDt49ZjBOvbBn5VFHRuz19vI4pBmWxxNLk8RPGCOe/CgiVPecOI
gbvimriP40n9VkoRlHLEs5YLNsWai3op1kJUOlTMo19J6qaU7STafhd5ILxZnFA1
UJa+Xlafnw3lJK5EUM7aR9H60qxTVK96zQxnpslbPR77PBDGPmGD4hq/1ox86dHV
YhWAOajrCfQvLRQl8lNfZBGSzcfc1YW+fuJ3bn6xAMiIK2yU2ti1HiXOOEt4VIEO
wGkANShY8CW3uc+etzxfJx3h0SqoLVnsT3+e/lwIOV8IterC+KKfj+fp+777o4YN
v6+N7YEjIbvm5GW2FgDRWL6BeLNOmmDIATDyNkdIS+Hcs8jfAMrXaYF3azs6Yzxe
MohKcdA7REnbLgQdA45ByqdtVUvYEUc4Ggu+2jmhtj5rJlNI5lmm//okRv4BHlMd
VqaxFNtkFYnD9gWqKZFdeatpoCaZ+jEGUC972pUhuJgl0BACxmltn4EhtMLtT0zI
h1BqMvy74O0f6HwWU8z/rE0olrbiyh76dJXutBhm9ceQGtxcNqf7cVwdyQWkTZcl
oRn10Xlj8sSDhB/xrJXiYLshGAkDAe21dIm16K6xfoWy8ATL4F+o4QMFj8Gh74cz
nDDSfDNB48VhqyuYaPDMyQaLD0ZDLy7ULJNV8ls6USjZO7Vdm8AF/61cBkleCzF0
cBvbqld7Zu3Hi6037f8KgRh1e0IX8XQtaFJojfX/wFrxdQKZ6hPbUJoKjyZc1TE/
dU8Sem9jZTvmB7uoDEeYr4bKK40dsTrJik/hQZrJOBa7BN/Nt+icXBy8jycCkSUH
o6AoQsg/9JCWHHhpbNxsBoB+qzQa+/FMWmx5pblqoPxxXrKLf5WHFNWF5pnUdYg7
vstqD/lZ1klWygrFxAIIev4xdw+JOTP8R7U02ipGxX9V6fw3fjXzaGnABR+KHtXY
mAUiL1kP6VdS01ZR1CvhbgA3joYeHLKyuHNwG1HIj9OzuX/hZrV+N1Vq8enxLVKu
ER4R7MZgK+aGKf5PTRDw6GH82MDlojwGsXGloXrjypykX5Pe2lUBWXsFoPK0sfQe
RwLli8hktR4L3FwBoCehhomFiq1Iq9WlqncmxkqrfwnTI4UjUQ3k1uMb6b1CDt6b
oZez1R9mm16SUELcKGkudl8Evln5aGZB1q5rUz/6ghaMDBjgAtXVczX9FA2cJFvG
l+msCrYFCNC4RnpzuvjV1ldBihgiGGryC+OYSTIkO/ZZvGAO6RZLXH+8oOKMtRGW
tad6hX6QfuECQzQS+tK2l0jH6DOfnAHO+e5l79kjYMnt2oC8Ir6lQiX+PcHXtZ9v
CIRY7JjFJSAtzad9kZ4Ns1s+dlC43sLc8tCYGqvEOlEX2gT3L/M2Nsrxs5oGTZNE
`protect END_PROTECTED
