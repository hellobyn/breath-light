`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8GBUdPXqjNNXHqkZIqEXpB9COOoGe3YRqelaL/GT9UnGuPEpkypn7tlGvVgOwI2
0bm6HX4HNWqQoXlOa++Ag5PT1FrCk+4bgAIKDQXfWV5COYgmVi649eJ+UnxC3hFn
GZqYfCeh/MJOBSjuSk7Uo4wy9uIqP1V4BGq4Z3f1/g1ih6/Ruex8TaOxmaHI6Ke0
hgflKGbPhoii9DGMtYkxVcbfN1Z/QU8OuIbzI9fzq2A83y7bAtrP37DoDkXFPfBj
AgnADR7Z6vzu3NSLq4qaOV9eTTcbetum/hBzo3RxxPOFeaYDITUWy/99ua3hMV5d
c6drBQqfBEVjpX/NjxPm9n+uxmieGsyUz0USPG9hO5s6ajKQdsQioeaQYaHGxfEB
ZSiTUS4lMB2mssM8NDBZd93xVy18zlLewp/vlSi8BDju5mIxaid/7FTRGb2HJOaH
A+VaWOX/zQHmBtzzMZ+NNyLkUHA8TNG8irwRwiWcz6walD/vRnh2UuMO68r3jsK1
YblC0PjkCwcy6DjpnYZTXqP6e5xH8ls4sA9xqzl1oNB7Iy64dOmlcjyuNOCNu2lE
JMAcZ49rmcak+/9ffGwvgl5gKStd3fwEdJonvbe7DPKp+S+uxWAyBvOMJFmhS7Ji
Iws6LQ7prJLU89Ue7TTrFlB4gFhLx52rdzI6K+wxcbnwVFxnIydXy2Ixr2D9X6ux
mwQDIWd/uA2sByP+LpJPoNWNcWw92NRdhVEJA3fVPMQLQIGqzpq1ASyAmnTKriDA
nBmfrX/vdklRr24XUcje96qcKcX+tb9//Ta1+YUmc1usn8ZPiMM7PzNA73dSpXuL
Ov3KC7Sa026fNZu+cNczSVL5mf5WpsnkB0lVGPFVx7y5CdZOYtBzwC+JwmH+IWtc
wVu/XAsvh/ZvG62UmIjrLzpaKkHI7ItmF+9dA3KMQd6hBBdi2OZECwr8OAhDhLOl
wVd/5hEP/He67MEwTxeBsnndKj+QuDQO78GH4JV+619AllxxoDiAR2ZhR1WbJceA
Fmx+adAZ3ZOrSQsN3n+Ha38jCHlUURze8BQ0a7gMs/MOwzOxTnKQL51WfVwJ+pyY
zZE8o2KAI+DfWQ81+8PW5/Q1EJStoJlNO2Ltn5UC5PrQmykicsnIep6dQL2NiBEN
FIjHLYcR3RlJYDd8+iL+FOBdj1JvCdroa8x+mFOPbZBx1a1MF52M2dbs8ibe3swx
eRWUYdufDCt7gCR1fQkxpQ==
`protect END_PROTECTED
