`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDfuY+iplgOWFt6vFj5NOH0ccmAPU/Hd3A9Vbx6zJ6wdvJDqjMYw8VW4M3LBg2/L
4f7E37I5QjbfD4Eq20uqVrqptmbGzmowZ11RNUFqA6qzdpJeFGmF3ZpOYXYR8T/K
OUmIX7IaI+KzzX0nqO0EnBOZzBrgkN48lBYUGkgXAxBldW1PnIMhk1Mn5iy4X68c
xehSZ6e8UvzNTeZ22CXce2oZvttq5/UbdDr9NV4x1sraoOeE0Xu5Qy64F85g1pSb
E7ogOs7TWorzCuenqQQwjATtB+UsvkuvVErYQpbn1Jmoaft+3nU/wNTsbDqI1lWF
5KC1j8Vb1JCxw2usmlYusUA2HGWSlQr4QGL3Li6hkReVSCCPi++qlAAO8JCudRJ7
BszMykDiUMPaHz92F8vndcxFFMaj675qay5ENR186eOJDmq4BcrgFLeQi4VXVkfg
zlpapuAuuR3it4ZP75IvDfbnkF9tG8sNEy3QFfSygjosdzchQOqBNgIAl/y8i+Lv
rD1N0CnaIuAEaEL7X28N5pxyKs19NFMcwcn/1VYgdevwQg9ZHqOAB68J+m9SbLlP
eTNNP5Z0zetHRJc+1GcKy2+CbW8IuYaqKIe6MB45epiA7o4iG2bi8a56jlxQwuQm
iJH+qjCBAQ2Xt9CpnVD8t+BNwYk/t09KlACEzKIp2EMAamDenjwxkjThg1sZtOi0
J5oHp6hbZ2x0g5pgi9oeyiDLfeh2pXThdY/JoAEetscqjaW+E/3N1Eg9KCVBWYZ/
pLUMEPS3ZjjTETbwCCAx8HXdmpVrqEnNyK7NxiBjXeAco9Sp96Kxv90GNhfvqJcU
Gu9i/BIG9JgLE8D0LxXvLaDCRhKRTrGqKeU5w0lTA0MQNDNkhBLkuFaS0YObWxcT
fKubcT/zA7Oocw44jZ6JBiAUpPzFgBT77uZeTurTx19k78SSKlkratADm6qhZ84A
qbvWbg1tjSsYEbgt/HJNBgazXprq7IgKGchImniTPBgTYb8uGkny3R4nYjD+FFtk
odMpQu67b4q/oTHeRZdDhKfGrr8yTlMfukwaare35yYd8bzEWxqp+NcKoEInRCXW
8lBYoR3LN5RS1nL2IZKL+g7Ta2LJ/sHMrODRNoW3S9QnBBCafeN6L07bVl+1cD7U
ybbs4XthWn57ucXK477TaqymAgxngEDLM1p/YnjZlJZg01vEB1IbExYBzOuh1rEs
IQ9slRhGvYlDQeQmetZLEr5WevOZ3vahggyRAePGK88MBqQv6Ib/R+hhO+x3A2rg
YcUO+obqNDYX1Ipegdtp8oojobPPG++pJPhgipg1eBGb44SBewEh2XsIlm83lz/O
s5s4ANzyntuyxbP0RL2hI52G1FQaiKDf2JqCnd+yL05NiRlC0kq8zcxbkPsL5ZDw
50+scEyb+0ye0MBSW9KVwWTMcx/kDh9K6hUB7aYdtY82kzV8UGP3TF0LEjc3QJsZ
`protect END_PROTECTED
