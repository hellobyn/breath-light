`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtW0GD4UovXFGB2ecAoEBjc1mG+3ljr+FHSFDDRClpkURfuHJ70v75IPCZekTPCF
imAwyZj7vL+uJjsI3BtmslR87J1e7dp6ta7c0XXosSRAUG2bagbrsSgu1y6u7xkr
jm2lPygoAsVIj4jp9mJC8kGyGx6BZ9R6G3e7sxhJYYBcP+C2zh+PicChlCxX7w+6
w2SPhFdgitEeXrJ+v9cCyEEjUJDfM/o62gendUdl6auu5MY9T8Xgl7JsRxxTO5Qd
ObB1d446gRlyO8cFQ4gVHdEbyC+FCdATc0EycD2u2fed5rLwqe0/qWy499K/ERQL
Qd461ACXzKwk8b+nqr9yA01abKbDDuVpN4Rc0JpNJEsmYI5MC6B4DyucvpkpWDYt
ZCOs5DnkTZvgN7EJI38Kh2jJB99fP7Il6oxiH93OdfY6Z0gLgFPBQmqf7sW997jp
OVZV9C7DB0FT802981a4/v/YLtV2I4NT5kyCDUS83sLFYT6r8nDvwQrCmZSyDCkX
uYk7EtfByH/DpFXMTTOGAqkY132jQ3p+Ab54F9MufVD/79TEYz7c0IT1zEaYNc86
xz+zYK84CevDJip0MbTuf5AQrPWzbbewkd0qd8JVuRHWevgS1y53izv6/5kndaGX
2Zz6R5XpPtxHTOZZpcMTP3Nue2P78ECVH4tq39pPFl1aIvTeYiAj3qxm+zWmn6E7
lpSPghofMLvbg1GFU7ORsxht/XxvuxaskwlWIKVYcWegqFUp49L7KR7ltmNF1NuN
OJeXBA8pVHP492+oIi+nwzfNDbsjyrA2L995tmsLRZbEE9/FZ4sjUNc5CkY4FEMZ
dkx5u+JQwulUYSJQkEx7s5ZZFej+ov0WVyFBdKlpzVDUXcBNnaxOiSvHgI20u117
cYhYxTYSmhVaDJano98mEBFIIEcmOjIdwvJjRip/Qy8=
`protect END_PROTECTED
