`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hjpT5ny+uTXsYompuIoTYfrMYVJ16+51DVbF06VPtg4N65GA4wyg7pwWH6HOA22
gNGse33XQh8aLgdMZ+VR4vHUo95jK5CFQJvmI+vnMqjDoLqcVJrT7vujplzYNC0L
GTq+rFnduy8nxBbDKVGV/onUdXmN4ryu0rEEYwGqGNNTqXQrfrS9TTfC6r9F7KC7
Hui/yEczvHXC2hr/8kt+4hL3IzaVF0cGKpFOsvx40fIrzKyGPk8peCWRDvggfOpm
z/mtO1lvAHH/lI94LbA/6yOeKP/gacyQFYofUPLgLUNmZFrc1e5EaX3V6JIWjWND
tB9otlPa+TOOp0IUEXsX7+onq1OYZ3/I4q43/2M53CvWMfJTYG94ZZTz/sTiSccq
ugH300XmRJT4Mnq+iPffx/XpuUfENPdOoCY4qoBA0roo+dDHjCm6eMF0Q2Tf6h8i
Uznh7aHsC1sEGmpsALZLJ/ZjQ7esQrCYFr3qj5ynUuwnlA9cOyu06uHEECfDVfe4
fQe6Uptj7HgnK7YNUsguDPTVQclBrQ20shT57rMH/9oZHgdQOtdI6HnRg0cVEP4f
WjIr3xYr/Z3DdLTqCE38C02VQBd4c0JfzLP7jcYbhfeE1grKY+XTl26CvEOFyEZY
V0pk2Iia4uBTULPMIcZ0CiooE23P7SbSSIoqIRTt9e3IMDq2SraxFETABHjPyJV7
c8YKkdLoPETQci/VIvLl0eDnotjsazUKlz/Li+SDByDB2+8PCrchkxwY9b9VA4+b
7ZvxbcrApNmF3GlM/UQid+VOuP44IVsnzQZg12UAzPrSP0Zmmf2dfd2x7dwLKZd1
FW7TIJjv4SXj+4XN3XJ7tyQDNNiqoEpGIHzqnVG2sUCHoW6F7aqH/LhjzOPmk28l
X1C51FYkpySdQjWxgUEPPWd3ICl2cAMoNGgBiLC0W5kGqb9f18iemLwESoL+jAdK
O1xVki4HaWqpjcfK9nTnu7SAtk+i+Q1bZ73ZjJfySCsTJTUBirZzVGuHGrCkLXHS
FTmNbVJO/tH0ZGhLlDyw0h2LQqTjB7POfHR7lAOvEkMd51s8nafZG4IV/tz1JTSo
2HD3LC2X4zNbuxpec4eAbOnMtpyFKvNpEQxY+fbceGqPAvi+Wz48ITZyxuu3E3s9
qf2BxkArVctpCCjZdAGtzwpmSBvPY7H5juDp2rk4sUAHH60bZKo40SeTBtM9m7v2
7AMempHB2BRxwIkqVUkbw4y1Gz0GPwyHngq/GHur4631UnOwbU/Nyz53pBgwTDze
TU17jBrYcRzGz62S70j9laMQ6xFYSD+R5n0IuoXqtpjePXcELRWBbaJ7jDxX/l9b
MjSTFzlexVz12kbB/hdCF/bUZtii7i6qxwuc+MN7LoRu+RuGPPig0o7jX6g2oZsW
nzv9Ui3FYmHpuHI9HEToTJypw9P8ye2dDDbUIqx43hnBrnjrh5/WLyeJBxxlEd0n
S+nMslV9AcFvyNQfRk0lw8LT0ygBB0CvcTjtnYIl6MBhxS8eCvGXKwQZeVfuZzRb
r9GFsB2CgPSq7kaTK2p5y2Wo3cBpQpsNRoN4FPWVnxMQZ9A19N4zAIBGXxvnrrtL
49z1/UuY0AYxK3Cxn5GxFPjuvGOzv33Nrvl8ihIKGzpdjDW1sF6lJJc5kSzEPDhZ
KpqeaW3RekR50NI1DNultkLRV+0u+iYw5CufcCJKJPh3cNAgrDJbPZd6najhO9+k
nTZ/RSQyZ3XcRejM53PKC8GkuFpyy4e5RDADrI7Paco2Wu8d71YUbEQ4E9an9ECZ
sDsLKUe6q7W5/xn7Qz9JQh8HnV5ZiUZD7qspajuTD7322F62j42bU4x9yTEE02HO
k8Qk/8AODk7bH/D+pVDuO/r6Ndwbw+1aKZg4kI7tjUAVZbIN1jgOXb5NophTNAo8
nSac71ho9qCKfZm4dvMIbV1pO48YdtON4tNQ6bqpbgDdK9nZMqLJ+Jcn0oVcw0ZR
pi54DJnI02GKFSrIYUu0A92xBusffeFAkfDt0OKg5k1P6FcQNr88LQdBP0S8T4Uo
ld90xsQ2T4WYr/zL/K1D51Bvj68WNfroC2IZj2pBDr98bfz74lCvbVARK85hJLmt
InLNWVfyIQwzEXYG8wUOAlt1meaHqG//MYg+Wn8MvpHY2xPcEB4xqoFdKltRvfEE
8cewjFc08brGEjcZZnMQjF3ZMYhGHi3b+2u3UtS+q0wzW8wgC4Lq/s7mpqvqNWFY
E4pRb+MV51E24uoJLfpcmrH3fU9RTIu6++svcSDL3PURBt0g8UJnO9s98Gtsc+VX
eGx3Snzy7syh7w9ursImFUgFJwVrH6B6w0MtbAU8LaghXBns6kqNPC7pr7LS4dkz
Hyhc64lzeG3rLVOE/o9LiX8hls/QquyL0AwP0GYrXAPSAp/BStqPjAgTvqrnxHem
sVNVGsh3pyPF84ztHVxTK1o7O+Zlj5CLEAZcOruB3rJzR26kAPE2YmeCX8i7g3jZ
NpWCWKP7nRO185347Hf5az1ZCvrZ9F4okF1f/XrrIXeiaVGrW8aTYdfe1Pj80ziK
kphBfcaTS/94ejhlAs08RtDaMypbzZbYihD/MuFb4CajrTJeUJnZG8bCMkKOD7s6
yCoGmH/gLOo5Xh1dy6VKtqWlJWpzr7uwfnzxyS4cFNQfSRypXZw6TRgnjSzV4b38
hdxWhTO9UUScrazd5IOwL6uaJqbWApSorO980vOPxmrFEPlV831KRqof5RTi0WM8
xeEuNVnLngaVzFIuNCxVmB7UEqD0X+WhYc6a4xoxE0snCQteZTrr6oZ1X2Qj8jLp
kA5QjDhlzgC0lq7t+qrhEbwrEz8y6BZ2+HEJCmsHvh0Qtd35OzXgCwz01k4M+Z+M
9k+bw6w78On0cppyQznvevkXFpDXzZyzRJ9YtUSodnoJNl9EsW+gTGBYCQ/tZj7e
YOuqiZzkF78RKcKEzJIatdO+xKhS5kYxA7Ke/gqvyuvjfX6fcH0exf12QmmpQ06b
PSndJlsAg7QQIMJ8q83g3XJoes2bM1m4bQOXpf4ObrXVou9Zg/4BfhTfB50IQBc4
TJpu8av/eb3AgMufomr0DzW/IMC3x+9RaT17xN3lbm/t5hcAd6phVBit2fTbmw94
dq+kdc27CNFgGlXAfYav1F6uCTXgLjkBgmdFBz/UiqJpCZi5EazrqJt1y09QYydm
YRqUJYVMmNpRcrVVwy6nFLApPFcfhJDycpjbT4Dh4/nSaAqJyzgr6Lc2LZJ0fgM7
rGxRQnHEek6o/cPYQG4JM+sscqPEF5e8QsDZN7B/gj5Sf9vddA0o+WlllgxBulJG
MsU7MmiA7whdkvwmZbj92drO7qTqgVbhbof4U41d4u2ybq3JTvkAuFBsjcCCl99e
/rJr/6TSRAnvPL1CaBqbfJy1f/4t8Uo+bDeDWNkojFLvOOhibgz7bQqOoM33h28h
vY6MVj9VWbK27j16lGA0mYjfXHoRiAYtyQ12iA2VOSJAbGgxOPVgEJHjbsnbzYHk
cV8TVCQ2SapO1q2jOsKDWabzDGCUHmDR/Azc1uyJ5GjpPuQyXHsXr7MayGnAcdsS
P6QNRywdiLnIiq4lSFf5Wmtl3YlGnT7hbr28rRCFL7xlzx1PWpt2hPz0Oif1/9V1
skk3uLjOJRUYnMha/VmTvjaqi+b1MOAwpmYGOlPwygxslmmIa25/CLhsw2t34h2H
/am55jIKQ9GU7Z5MQnzt6k6k2OgkZ8qlU+8l00xHefK7GcIzmDXDspeDCWE14eyv
Thf+Zn0RXsvEyJOr4mIRJwVG7PUwM5gCI23gBWFXHrOeSxupLsH0mTNauyM9wQWb
/vP6C0+CZkD8pcAumTQYlCra0uxID3jXHu6wxfAd7TQN9w0fKosgOUUUTuYNoRiI
HaeGvKo8vfkCxzC0LHd/OiUvFbMPmHBVozcrW+I8IIYLkRS8gt9inga5G56pR/cS
iLAmuHX4DzwwGt0KRVR+Or1KcmbVLDJZl0kj/W5uIMyKfRqW8coIve7Sg+/Bz9wM
UitTpj5GyX3ZsASMMfJmsAIVTcfiYNmdfdgDobEIjrrnLwn/iHIiPsLTNxlxbBYU
jgoB4M4zb00Y2QlpmB3vp4xY1toM200nG0jv1+bn+4gXYQwCpot56LTdsqk7udCb
eQWqL9ETZmMCj/TXtmhes9Y1ur6qlyFOnfwQ8P7kOsVm6MDBxnLNefGwVjAvfViF
Qotv5KTStbsQEmqh8kfNy2V/Hid5bkxCa7jk8Iaralt3CQAn/fOfMtwfECCpDLzd
b0kpyGtZvYBSdyyrPpB1bC5XwlI71uf3HLJBnpTcsnu/F0tJootvdJLSy6UCnq6U
fwbLT4nZhsFVd/+Spye+zeq8GO3+OC1iGl6N/MPJoCcm+9j7TGod/kXHF/ssfgYa
847K0VrWOMIEdnTrjzofnYnr2l6af6b7oNYzCIvmGYfGtL5hxOHUP+u2VcjJS8SV
hEFNRH8D58YCBW6C3Tksr36IKpax8LlIvWMquR73N8UXJseTSfyDo9jzAspRQzSq
erXaAPtPsZCwLkvd41QZR8fKZ7x410i995J6YHqpG+zFNLxd4UjPG+Q/SsUe+Abp
nP3bNbYB5ZvgneBhC09COryt+efaJnxdyZq0QOfMPbR+EiGxu0ZOaUS0qjz5I0xG
mdH0Pr1n0HNA3ZHWO1i0UpzZoH6xIt41fs1C2DguafMVUoRfjbYJR0xkBh9r58iv
tU6dUKybDZaEUQzRvD8RhPsCw8f1tm0K21ttVBzmKmGaNzr/ZR3LcZZAmZdJ4yN9
C/DDE0+1dpN14dGcuIuxEfXDvzgNximK/aFA375bg9E0JvoSRsNRhG7NREzJk0+/
cB7NBvQos253JztxiCsbZRR69IiwwF1Dyq2r755D4R79vOwMbpCh+m3SSV/+x1pm
HXEBVSKDecHS97sAMnUFveUXgBZ4Jz9WkDpmRMgzrRRHpP1427XwiHQqdc+tjLOq
Uf4lID/mcAQiFLJul2BQyu56NJQSth4gSD2O65XCHH3PmHhdrgxy3yf1WAoM5IRg
TTX9yvbu+7AI4jy+5yp+vJikYF6Ncz94w7oeI+KV6vtE90Arl414QnDZajRhTYHL
wD6GSe+wjFv1XjBTVWkrk5eKkXowA17ZLYBhYGQ3vN8mMudI2GEMWvEcSufDfeld
wO+yapmQFrljHMCoR/v7sjI453BhUMP4AWIwnJQgNuhsJtUMAiGFacC3KSdJntcu
zCEhVgTYtl4VKJU19OIhINw8w7MuGU1D15ZdwdBdbewqRt70MCKDN3yH/TgvWTcE
8jbwWVCBhcSN+brDti6SNo4rBSt5x4wliyyx9lIMtOvF1y8IoX6imUNloA8H7bJ8
KeF/YJyMg53jLXLqJC/10zRqZQKtosdL8JnsY4Hx8EU1kduTOWxJiA95D0/7S2yF
AjLEPfY99r13ksCHwseSbv+xyss+wsNhYTvEVkxp8mNUjIr/wXIQApx48fO0Kqlg
vYvfS27B5YrSwNdHqIBhXLPAeaebbgu+hS9K3bmzkHvz9vpjwG5twqSG7Ih9GtHe
9b2MpwCDksF12ryobyywWZXdnQAvAAjeYnL1yxyAxxcuHgrFGcKdZERHePe3s92J
TYmFos5pgWF8TTyxS0LnJe4kA2PQBxtnvK00hfTs49L3a/qOwzOr3muV4hOApQR9
W/Om9dA5aAfwvX0sVJkA+877kiU4+OigiuyQKb/s077czAILjsGMKVY5o/MA9aUQ
oIEfN5Vur5j79aXh3MTVs+n7a+HtOWIctd9O/XeqET5WMwioZ7xrKIiBLWkiN5vv
c5m3xHNjY1rBGBF7KkuIgg4R/pI0YXi1ozLvbypN1/uCprnmwffPSUWWtxkVRJvA
E1zXwlN9BHABpjuDX7uAcNfjDsnc020RLFpcEp+g191Nrjc2M38pHU1wenLuqypC
jn5dpJChYa1b6uU+W7jqMGDiZyYJBb+yLauzWgWwTqzErbdg3Y8liPCZKMoW57Vo
htP0g+TSS9kWGbXKJv+4z7PkOcgxl11d1w+XbXLoa899lvW2aOHWnVi4ReMgIM8o
UitXtsXfkOE4BkZfbWoGGROILZyzuY/G93KFTSt6N0gMu9L1g0EWFouiqd4XyqoU
3e07VBUwdEYofGFpnh4EqvPn8Mr7ZGXQzRf7wqCV99tzlj3t/WHlufs4cJSAE6iI
3w1hGcG21hYoOBNr3kz062CJGF9ngu9EHVT0741a6+DXaMQrF6fgpF5kCNnCo9cJ
vJdp4rOr70iMnzASSlKCNO1XMcx5XK6iQ7/3ovYyNlhqUPTjLf28q/XzXA2jd/21
Ja6PRewoYwdUGD9F/9E+GHYbpxHlcTtlTnqalnisNPgCwoz0MKiplpTiZOBXXH+G
pG20txEjH86pd7LaoJYZ15PH5nERNf4LpqWVGqq0wHdcNSRXs9B24MWLpQFPjIup
kVgQD41qLak3AZtZjTlUN59s5oJGnfYBdQ+YsPl2xPln8DzO3gYAXrVhuG8HN2YH
69CpqS2E6+rGZbYSi5vMUw6CWl8LAqb/20YOCFOXd+PV/YntyJ0k0pNHmXHhVFwl
XYZsPLqzhxLyrZMRCs6EDulAiBcMeUevW+ppNNtWpW69VEVjRga/VUsh1BIgLlgN
ZGLyWGOr1++1nYH7/kq5q+xYqe6SNWgzFFAhCpm/IMWC6ZebidZd0A8hlgZRILqY
aUyPqt7H/ixaiRectJi8pckTSAEREE5qza+EfiOzQ/xZDntIBna2OH8xHCDngM5T
Ev8BuaDC+z7pNtzqnnEnVeAMxHIv29hhZRD0nZK3F8QapXfP2WhqzmVM4cVkOz2x
dXz7MrLErSJniJ93Q2fGT7Of3C0IYTGPLcZD0fqLHlNWTEzaUmLVE8/KPPGIZdoF
JullXx9YIllMU9ic0xFCMVoCqLMYoRT7cU6NQMWFX2UWXJYTp+CQtapFeov93CdM
FOyfFyLMDceL1k3FlyvLLbcFn8ikuNeGjc6EdXC6EvPu4aOrbW1wCUho2Laq+x33
O9GnWuOr690Qvi7I6HeaGHoT0z3cI9YEdPmH5jbDYsmggdQI8PhkzNS1koJlZVyI
7If7uiiS76sLo47YG4qE75Ei0ZWsPehi3m1H0cBOpJz9Yl4GwjO00LQxG/YZlxy7
bQbykZzD0ia8K705wCOKeJMM+ZYeQiNeyGZN/PnnxWzWIjC34ZYwizJIA4vQ+K7q
MrwJhZTldfbAFlaPyFZx3jMjST+yIzLf7Z1z/gjC0HS4TaxeGupcEyEY8rxZaHEq
3/Ixvr/iAdDlZU+CjHAkwVSmJvCHQyJ8ZCFGx+nxjX0AS9lhKzLN9rRXKDpx4rD8
iS/3464FHTaLnjZ4Rq0+lxyis4zJ5neqtzdo1tzl2RHC/cN6c5lqb5PSWL2FxYr0
vypoNMrctv+8Jm1ECeupAYnN5bcJpOCWMSc8SsbsHvp6OAKli7kuDQ1SpfUS03UV
/T5EZnWThWXif5QRzcYAUwZ6UYe0xpOOcQ0xmahjdpRJZqt5+wFqoyozWiz+DuR3
iysxRRumgz4Q/a+7qyWcLuG4oHmwgBzgRuWG3356zkbMIftu9/wVax3+PpiJ19IE
J36thLBJsih5JXR6zu/4PcgqUl4LCgkLZDMkhmFWk4QuSNTCeWM4ifpYqoFl+o5d
2aSUjs0tLWs6hAtg5knOtCn2ZgVTBP2XMs7tiHutIQApT1nP6l4nnSybihakGM5G
jK9uj+o46rBpkV1Y3NgXH9/MrQQQ3rsNFBrt8DGa5RTb7fcCYOjKGhKywbBAoiMa
nXdMXrnTsTFXgxpVlKGoSM6ugY7WOeGjcIPgcvk137sD70WRcMTmTK1lH9dHrvRg
I0NUEnK0elraw5iYZDQe6vp+wuOlgJGCTw73LUVhckFkTeKkb6LW02t3/soMCOSl
jaEOV0I21/sjla4ZZjxTnRYFBmADBKMUcvkPoeqM51ToLQ8DRO1G3Uts1pWA2l3l
5SJi33UIBZsPztewlGbC+NaF1iLAys4j3g4cDy5Djh9UHZvQ/fCZktZK2Z2E8bP6
jdCBarB45D7lv0THHZ/Sb+sG5EtYae22jldlNbKt8/IOv67ix/QtpiFnAOJ4PrvU
wR3zhszfNJ/3w7oVuHowcctdmA9vxZvjzEOuYQDozepVu3Dt+Z//fLMZ9CjUaMER
toFS6GRpaMJLaLYhI21RfXy7nbu+Qh4ECplpWmvtQKS7nKVq785MH8Kjj7hHq/dI
LPHqxjd+UtUjf9S1C1IMOPIJGjcLvyZoffYStLNG61y5DfS+8VPz6uM4jiabGjOT
Aq0hkLJNq9CPAAhZvfn13wIX4/FmAKMw/m1jkxmsisF3x4bafX4nliw2eIyXShdY
VwRp5JxGE2lP4QZhyacIZGXZrSTTQ9Je9IFh5dKMsJfJ60wyviHBJ3AkUAGc4bJN
SdYEidLe/2ZU2r0FdNLSpgKaFMtWIUmhyIT7dZvdb4qqP2OqakeEKbz9m7XgsYuB
x+2iy/jfI/ALm1HNxKhZoP8C0zaaZZvN4FifUzAlzDfTRtweqAxicUSlcDK+Q/6U
xIBYcrmMZTZH9oDrGqXkpucUmkqBhjaOMFAH8oJ1ZSSMowPXpfzShFsfwSh7IwI/
2InqbRAfbZFdD4xGIA5FsyAQ8goVPcbI/aEdvvTlKep6hR2jYhQrNlbcDGLWC92G
U4rRr6vshNIUkQaLPit86USfUK0tn0OOKsimY/L4AcYGFk7t+RfaF2WxHkJk90Ps
UlZ5uif2N1F2wAv38YrXKInseyfR+33OYH7ksAWo/j2uzXyPaEfSZpL4XvQyRVaS
zcAEN7Kp1+F8yjzeggTTuQsKG5NKgz0XSxSvI+xmnyjsz3IGIvxz7eHVDly7aZjL
HFy5XUTWblRVVZceeRnHHVKjAi63VRtFxSMjfnY1AiHYb3/v3R2A6qQ0RDeAGG6x
qHbi4XJDj8iniTsVPBmVzVDV0mEEvHPm2+1rQpY9tnpMp7yln1kyaRYAYm7yeuUF
VzJcTU8xEaK8rTeflp9clXTgt4k1X0kfy2MtXVkPSIiXWDkj8qbAURHqghAbNzGq
cEphZTRSIQbvh7Upoid2vnFofPhykH/WJekQM0pnfSdPBhXIlbIhAfX/FQ0FIpab
r+rbdPtU+nDVz2ZBgKjJxPNjaVu/UOcjRYt2r0k4fu/nMQLkyP+ePNZHooSvGpYh
Trb/v3MQsl5pjNKSkYJTMU0KKVlJiUcB++U7fncUPpt06N4qzziUHY4NP4Ffo2N/
8dZ2f6FNhRgVbMkydNh1oa79rJ4rKQkm89SR77R9yJIn3decMCuCj8LJCXehgeQd
++2H6wOca8voyScpZ0eRXBs96jIlUu8/M/6lRfTIgOBa/qH2W0/9Wfym+K7ORRUo
fBh5IZ9x+mpzxPhi1CyIBNiI16VmaggDGBgRRQjAqKVsAd3dsbAuQznL5BzzIbV6
QRGsAynp5mJONz1DOGp2hm5TFiSVHGEZ6oyjUrTvdTIYkdSgduITS6J1AkOhru9H
DpLsu6KnAeeIsLGF4/IpWrFseEBJOXY1T6xwT1vx7vzuVRwEpeCFgW3Afqz6TMX3
FgaIfxOzDGyFJ52OYtE7ik6D99sSyiF+RXLNV//956whsSKxXPFnA4jOOh6gIdfy
gR+KWMb1oRVtLdl7zpsOcqXSYjp+amijcDVskphg+AOvZeirckcZo+U/iKfToT+8
sHlbAMGBnzvHWTOQ5g0EVt1PuGfYxXby/yYqQK4fCiX5SD4K4Zfwi2wsQpQs7P2N
gK3sP4OFUNp47boTNP9vC0UlkEaKNaGo5vZm8/bxGlCcuzX+svxTDAKyWoyxFgqs
Tsig9/Muj3YfEym5ou4mn2xKZ4J3Wvq3tErO5ZpWBK11E1NRH+67FTSgwOOs4Ghu
LHQ/K33Wny1O+zrGub18Wy6swBaRIsOSFwKqszFrr0nkouZddsRZl1tKlXTKbtks
BrS09BJqSbMJnisVCrtIT59MY5UFdnFTwkTBGu2NtY51e1skNc/V/fh++Q4A7YYR
0WJrpGO6ej0gdJVnBB2HDRYjVgX+4itmYEMn5HXtCxZ4U4znEtdc0/9HkyM6+AGz
Cdc8b4MC4RBinWPcWgVcOF39z3EXHDiJ9iZgXwVqJGFauylMCFY0miMYuFePahSa
UzNTanQ4TqLnvdgZJY5rPIokow5fqAB2eXlHS56pL6sh7VZmzgWZcceDypNHAoYb
6hDe0FGbvG2+OHs9BDuN0VPMT9CvuhdqRACB2XHYUpuV9WC/mlfJVODGSmL3oYti
/6E9xazx7xa/GL3pSipa7KR8KQhjrBob0/fylkkvzvuUhkbFEdOgF0rftmNxcIdD
0QJlug5PzN6+uWUdGdE/OSCItmajXZhMOP4wrAlRUqPPSfwWpNRNrULu6hcAKYb3
ELad102P1t0YPQc//qWCWq1bCjfxPdnIXvEzjk11+DQSDCjkzueL9yrbIUFvM3Kn
BWff9AeSOn4XOIXJpEG6tl7FWBxmnCMFIp+qngv0mkUqbID/fMk6GPEN35N2z8cP
lXoyqmthNiZPJgvBHlY+Gld0+sJLmcN6ww9WiLzE98TndTX9qy4GzF75V0DnnaD3
yi966BkY3XxdmIAVaRAdOAR3fFNzSS3/M5IRBKfpkTasp23CgQYGo0corL8ozZdw
Jy/JakYVKFTaOst3evNhy8c9QJk2scHCo/+sX4TXuGRJaBeBTiRoFKvEKtF7ANoL
L93nIp/3G7XPK58rvoul32sIrAWwDjiqEOp17qzyFuS4MMuY9+nQOJyLBn9Ghk8S
XBZVpmQFHaCmw98lMavVlQULkfupb3mwuNVhaJes7SGLb1ZV3BBI+Yt+RK6KVO5Y
lnU7c1D4PoU8eBaKJCs2jA40DgiCigNZxctHxPGPuXi286iohskjUqIU+GwtwQX5
CR7ztPgPDl5jVRsZSdz9f+bBWmGDF2IUvIXvRAr8kP3qVN40ox524hlSUPzIFem0
dXiXjvIJFOEh00Ycg1jyqeQbTnPSHwetx+t9urKwpr/pRsjPBfJ5Y4WsPr8p7KQp
Sjju65Kmrrq6+626EaaMQQUo84fWSa4TfvhIbexSs3b9COrio/K8Zf0mG2I/1AVi
N2SIpsBwPG1teejFhyBiC/GzBMqwqkbv8QR9RLt9ctzRGnb+v5cDcG8WfQCyjoM+
/4NRb7gOz0g698x8Qv5NwvHLLSLU0sJLVsvRCjBpw5vvSgJE4LFuqvM7qWZXf09q
RqInHdr3EaLp/yLmgV1BGAiuFkELZbSu8j3ZbMhTSoptegaIU4jRxi6FS09oX4uf
fxNLNDyEfn6qjOAq5B4OWNVMInNsusXxdJ8KJz9XUCjGXF2H6SUdB9mPeePeDVl4
TKlwWHmYNvIp4W4T/nXIpULnl/idwJ+nl6kyZndp6xvJGkqLTJ+4uT3CIdSbkhJf
zsxrpZYTXB8FxaPL2n9dXBlu+rSF3ydCOSlCuZdhsIHB16vbDcnTEMTrcPQUws+A
OqqCRC+73DcreJzjo1E0H7QgbF/WNdEBTV8TTSv0V2pNiuBYmKSzGIvYJvg4CcGR
FVa35ynbkY89GpZz5wXxTNUW0PzAPgM/BYqMefRPseYaGkQnS0Jg9Xo/xbKy1fXT
fqUdk5VI7A2zv3AQYNQrDb0L1ETfeejwguRYWlGnuHoBg35hGdKGeFyAoBIau/tw
1JSM9dfMpXVA+Nzr8T1GCpr3LVsDjS+wwjeE3FhT4k4WoQIG6FcS8LlfGkWhCuRc
K2jzxwsvrYJX7vVmlr9sZSgRGKxLSUZjzcWfGVhFChWtMt5xboqlTkp86HZdLxNh
pHU4v/TGEB2hL2Tye/79cYPO9y0EOr8Zs6YZ+lKtzbyCjhRGysfTI1PPzph8q/7f
NceDWvOqT/jNZ+xctjJDgKjdYuwsPH67tVuYj6xtAE0Yie/Jaz7of9Mt1qS02SwT
IF5yWnZzYBoCeBQzB2/Ua7FDupY9pIGcp9cD+0W+8wMK/l6yZHrCnVzHECvoXUoU
9uJ5sRmleFutD2bRx2gBP50s370JUhjh0oicvMvVp++4CpENF2Kl0n80nGKNfydX
mezCagW74aw0CinldSqLNpUeuP9l2oKb8fok81XmCI0NIXPskFDSQkQleT4RlRmX
WXZPB/DVT0ecZPr+1EQaYZRq+UHUZSGIC4vDJryAuj5Ikrjs5xJbrhRXty/CsGHU
owUzac52/ASlWjhZDtmWOBsNkc2I9MmzsBXDvveRNI5IVRWUbB7GZ6aFdmPT5rXn
fOu/XBDds0YMwAoUU9GaabBQJJWP9ejAznHD6fOeFrZx3QFZtftKkSJtxmSFhOU7
Kb+slLJNc/s6ba+sSo62NkL0jWc4sCBJNch85bGx70nIhszu40tfG+1ROSsJ2fmf
1QwcUVZIFkD32G4fT7oc1Dko/F57uBKJRaM0uZMaP8fptiHaKJSEBzBqC6xXTjEy
pVtBJ0rDrNby+XUBWyZyhmkSPukMLrVcCOiEeFpqK39lpgPftkCeD6NOhnQPYv2o
hx+GRWLLm3+x5MZgX30JuaXyEazHMqxLdLT6QeslV9AMKvQmEl0xERNcSaO8kJqf
6iy5w/KI7srsv4pLy1pIQ8Nufnjh9YAeDYgKXd+apuBFLOkPQaZy99FUtSLgWzXj
bqi6B3MdSSTw7xKh9llG4+JmAtm2+x3AqognWNMpzOKvBeV2KsvENr71F1ZckfKj
nvWuLLQRdVSXKPD0RBxXNtSX21hHw7n41L9Zvw86PGuP55o6lfjMnL5eeMQIiXFj
ZXz8Roa4J3OTGp8FxA1PtlK5jA8CxitdPbgaW9eHBRVkUjQXiYQMvXZOmaq3E2Pj
mJSKhRAccuvhl2K5pBdPY5Afg4hH0is6GMtJV4twrRdJjOTnQu5t0TPNltSPQMoI
S8kLNsDTsrZEgEKwlGX+qK1Mj2hv5/1/oG45bjZPeTkLnZ01U4Ji8BjlO4DgvQsp
FZJ78kcKYg6Mj80hUVgTdZbezHhZr61Cb8dz92zbTSHeG4BNPI4O07AZryrP3KrM
907DWJsp5CbhByGIpZjpNVpGKD+IJn9XpjOzINl3r9Tm8TmHmv1F2BCLV4u+trev
LGaGu1Zk6JR4qQwMl83adpgW9bU8JxdEDaiuGB09SSDMIXLOEDbjWvQWYOmW5etF
vg4vpAojlb5PtM5bY1dJljW22ZEjYuZKKkvFD2OgoJAUiT1F3jSpeTjowxgKmzpz
IKTw0TG2OfiuqR2pQz4m96QFK8xc/pL0BBq51ECuGcX2HYemoSCNYZ+9/LGZPmL0
8LZ1YRxQggx9UVfeXdErHF0zXrRKmme9U7646TV6OjRlNUBC/5sbCFOnDeSSIGIm
i26oGN5RKRCs3VBM+MsAIxKlvJwK/twC8SE7TbpdTJdPTD2YKYrclBjF5n8z2pN+
TsaMjw2ppUu3/wQMxiNqfXbDUh9psNhBAEERgE+le60EjyCxn0aUS+S9xGIyVMW9
U48c1LtoOHoAEIJzZObrC7JUxDlm6gWeCM+xQEPwzibzKsWMxg/YIVePHQeOSOwZ
SQGvio7PHEOBZpL8ScSlO9Gek59pEVkWZDO8XsbFXdboc9GJFl3mZZ/uhk79b1gA
Z3jhp+JdvaQRCGG8SDW23wOQJW/wgtUMV5gEbUWLcqJv5mBf82dYnSkKxg5eRKCm
vY8GGddwRNrFDRXNJBNwC/+PaJeJAjO1/cDmoNVS/4AEEhTDY/vtTB2Kf+qDEIBr
LBxKl2FyoGDN5Wgp4H96Oatfw53J2nHlQJdCLIZRwukX8epUt/oVHEkhyYJncLIl
cvWExFl4NI+oAUMpPXi2PI943SEXPnCQcoIx7cPKQbO5E9XBjchIcHNoM0HvvDMC
Zvun2cOLQqhaenrubWV0YP3bGmT3DPhS8gtEnmPZEWgUwLRcRNYtheNTG2QyL6Nj
kJIapz0M0+CmiEtSlHa1K1lLL0LXY9uZ1QYQiel7Nyh+NPPyakgYAVlE5J0fFqPt
uM1gB91DsCoXNiCxs1FrgobRCMG189GxMR/J4cOk6u/ZwXKXYs7qqU1xBaIHXe9n
OlYYmd9Awj04VB9wY3qgOBQ2/YgIt2MNkNphnIr93jz2Xs6o/swBgJ+eQYe3pRj3
XR4b7iA/T7D0yOzu3I1gfpsqYexjlaAL7XO61j9rycMVCTI7WowNL1/GzE68eN9+
48pHwInRMVAvm2kspAoWLX4E4QONIFq5nGvjMFloQ1DHQuVnXqK+rSPQKIZ4JRps
NUdJJld02pYyxmLQCGxjinbgkRF3Voo8aIsDyRSFQH5eO0FWRg5VFE5eR1arLCvK
/dHMylrVHFB+Cpbc0g//wNo5dlY/cabHhSMFx51xdLrDte12/SsYlU/KkQbCg1qR
0RJxOolLp+VhCAmh4adiJfTwWwLhNYFcMdWKwMrZWJJ+kLze9C0HzbhfacaZt4ny
EfpBsThJawGrLDBL7TAOBDt0iGlo8IR8tLSR0zVEtPUss1Bzlayl8btsUM7F6H+N
0BOu6gQexBbXZpVMHenkMmiXrnhqWfXQG2G4znEjC/Tek72puhDGSG3855PUiyfo
Y8guUyqaFe0qkU8Bk+aSnoV7ey/bzXq9QriR6hTXxEnG8sGXqQdEMYKSoeS6JNbY
DY5y8AR6tQpex1+xkVk6iJ5W0p6vI7CSOR+fO9jnLyr+bu8uMp460yY1PQ+Gf7/D
oo33LswSH0G1d5GYIKrOHSLE/QxRCnWwmHk4ekVowvQMUFpo0hE9jpOpXQP6ucse
5lHSczHd7Dd6ch2m7o6q7NgZHWvExBSx1SEkeqVtvGnAUcRVIkNft5jRm1GOJ9zY
gNB59mRNtkRJ3R51cWPfaQrp9hxNicHsoRTqLDyXpzhkAot5UZ2iW6Z3U+/oYTLv
9Wu17qNPqPf5d8an3o+6BFspo/wR8RhHDuO1Zh5UjG7ronlx2vLQgwG4jb8Dgfuh
A3slUrhqkWfHDLeQN+LEy9bqcn774wTTxiXC+vPke0FwkUGsdWA/iozMMoxK5mJX
RF+qeIO2ZLgfA217JxtakjW0H3SGgV2KjdRvm5Q6q8U5Z5voy6OHAQeA77dicTTv
0yjiMx4ZHCCs8KMK6GgrQinMLrNdlmDhSJl137TOs8WBye8r/x87vd3XmJZ6onQ8
H5AwR9+3X63Y+8s9qR6vVTUU7aq0C7z9sBuGFx+UubZOoPfRg4D+iYMi2qw7HF5T
In3ZlRZ9OxjT43wVfXqcQcMlJpqO68qIYY0iVYK+q+f+y8EbQL5mMfna05ICm/rg
acwCrTg45mXFzxLm9IzxEfcNGyaAF0GcfDzd4UaFLSL9Wh4rr0oS//YbbHKg4Heq
J3jm6ensCrO51Deiu/E6TEF+Bw1kuekPpLtPViEBejXqG8vLiPP5iz3KM+mkUYFp
orEuzxWALWm/JjXZkKJppAhovS8FuSnIsuzJiNhxkVWp/vwGn6Obm0awp4eqSyHm
AP8qjOCKNLdmJ+N2lMqrFKTUobq235xwys++vS9Ks/qnAY8ssBQJUIS+xVcaZ+lr
To2e8GpaHwViO7jRxIbDLpeemX/6zVKYk5hThPE106BQq1UvQtMflqUAgcMCklZK
Ddb2f//k0apAnh2zUf4kE/UeetIMcClVva2+dQwynA5yMlYuRfLdkFFk9tqt2xBO
de/2RO2PZfoQ9nQvBWI7lRVhGXohFmL3BsOiyeGyiHWztmyNmSLxjw1PkphGWoKR
gqqDj6zdzsMYqB1xiWNOPNANn6fD5qhSMya+X9T4DXzS3aGF+T+TmsXKNpTwKQmJ
S/omkiulAGDZSUmWxFXIzfaQp4xM9LjzT3xXxM7+odYExFr9K0UilahMe26ATiOV
MCrJR30bf2sXy4mPT0ifnLOaNXFoXakpAnXJaNWRLqa5m7EM7TwYzsP+xwigGAkh
O5i7f0MNf+PZhwDeXh/QepNyVn82O4M9XSAtOATiDoUOL429uVot/9qbptDy1KlA
YDRi421Va7i8rlUC/IbmK/dZh+n4VaJAxJ+WS+67mN6I8ocml4wUthB5rETeA3eH
V0foJ5XL7RTe4fqX2HzVC0rZ9OnpMD+ACmIlYz7i+xgAgA03+llY2dEwg9ubqYl+
0Ahlmy5BA57nyKiWOLChI2OAQnHhLl1O8pXUohyUYn5cvUak7t8tmjVthYH7NwbF
gourcFY1+OLpwgAUB7jLh72fuRfBPERuhjo7gyVzzbp3vecv778O5e3K/iiy9tU2
5mv3fOfn3RA1jT64zPmiYOKhr8wUjPZ1gR3suf2q9mAkujLQdsa0UBqA5j2palw5
r6A3f2IwliDYslUhKWFES2r5Qhqr1c4SWEYF/O6upYvRwgq2rW27Sd4xfblPVIBv
WhukrCIsLsm1vwJR2npugyIsUozatksQlJgTRaFqq1AbW4ksbkTISU1C8/07C6ie
Rds5Sq9WR8FsdrJg6EVDkgs4SD6lBMkEtrkwMHlAHCxCx24nYK6XFstMTpkULgAG
d9NPZt4E6KI/QUjO7Eo8Hg==
`protect END_PROTECTED
