`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IzwLQVeMV0uM9rHVK/FjOO80PN0fjwBPjUhq/+WXnqTOkU3SlLdrAmg0VykUGlK
As1I74Ebpf5nJkjneNDSow7udItwG+urmEYPLLERve756+5eVMRklfuSQvRvzdeM
J2Ci1/Q+tgiyvlfLkicAt3EiFX/d3Rsm+xwcSGWaMtNT4iXdbXMzMztvfK4p6lpL
XFTGJZkY1md7Nc2gQXwARHOe1FQd1ybfqwQVqNRyrDerxtrGbZl6BB0QgICqjnuX
5PgHlF+VA/jHIWgFLxkIcIKhY4+dv/8qPBgWd9OkYoDI76ugs6m8kWWzTxrN8fOM
8+WqSRSDm0S+FgHm7US8lWeCe4Ia4eJ0zUmDj9S21xUwQJbx3okzAQ0vhv6dftmp
iaw82niVTp0aiM8dylSwi+WuSE8hLYwibfWWbyLA7q0vhxvGXx9UDBoSQLEP+dS0
G+yYsD9LueGFEWq/f+77cMcX7TeemNmWDplXCVffTVgrP7qCYowzfAUPxznWxwRy
kzp7qMfa3AXllO08/Gr2eeTMaZZQTaI9L8WJ9iXIUABTwggj2caFLQGMnt1hR+V0
Ht3nevKx/blwc4aIgORKpSMdbWKsggvqRRFsNl21Bfo8Z9zfbemi0APDBSR9K8oh
TXQTrS2shfKvBZR798T2OSG0Q8V/j+9Lnz/XGbwcvZff+FbIy0vONPaD0DgEtscs
JKGCnw/igT0mdbYcPVDdPH0Owqu/lfc8tG8fijJ0B269+dJUWDB25ABfiZ5QIia5
6U+vyKK0H95EVWR2LkHXpyrM0sbVeK2DNJAhrMrF0LG6CathdzzYe08NYaIPzG57
WP/MpWLp/502shloHP0sVEpjSy0Qzot9WA9auL/AuJULr2RLfQgLsKodlMjZ3pj/
oxHYOQ0GbcAKAWEVogE9slzsM6ltDpYgqVTs/h/rfjC9Z7U/16dcUgYXSObrV8/+
GLq5Y3tSFfItwUbfHgVDyhU0ti61QdD44ueMYciNUTHl0pO5nPLiZ9Regf7xvrQk
xM5K5lHoHA0kwX0tYlK+sxrO5tlCa7S5JKFqT2VrjFZ79p0W09hd2enh9p59QDuk
1LSz1EHcHBe1J/fMmAuhlHH8UoD56EUHJ17DrtECN7ucOYccUgaJ59/hOsfGfLLm
lfil5FYUriFVySCiqtbDljgbQd7m81/zAxNObpmYffOlRUGZwcCpKsrOjt4iwLqm
Ny7EEZ31gbcm//VVCkfy3lRRcYDIOkc0yd5Y/Vaix1zNoP5nk3XZklUUpsdmnlNq
pK7R3gGJ61rOyE8+96oxufbE99RrHk5gozdvNzed0NDbyCjc05SNTTFQHNT8VeUg
Lc/5hnL3Hw+QrSghCff3KbnSjHZS7Taltk8/eJEtY84kkBshZDZjmKUbDel3q5Ra
niO9cQv88nKo4JakomWxTbt5+MMJfo1p3cDvesFg+ajbizPlTsc9rZIY+KNKjdoE
n/fWZ+3/iVrl2qVIc8BzBTp5p+bsLNL/1Q4xrMaKhYeVDqSvvYBnB7sUxr0rhtuk
1hjSAucL3yacY03sc1hcOi7UWJZGeyzRL3RvmhRymyAEklyEOgbLof6d+rbpYrI0
xmrZLTB1uv+KYTspuX/BY1RYFRAAjXB6Ah8ESQ1vxGDMPFiHlAozyY22gKNkt1d4
PAXSvnpsVyM6hlEhkXvdz+iF21YglCPg7KdHXqi04xlVGBphxqyAqactEKveM7CN
xweD21RgV2BE/DC2w/OoB+3gt6mDrIS12115hMcmnN/1GB+Ci5VbLG4QXCLa77Ji
+Bef9V7UdT7TJ5uFbpnXYnqG3/ZDWFMdwsSSybnYF/qKOwRFSgXzrIPWr9Di4pOb
Dx+3YCbHrnYZJenkI+IvH83tcPFlrZ0MXuM3Yan1RmAw0gcdK1MEbNOqi07zcEmI
MZQfmeBqFZoCTUPBubQEWCTiz5qU4OStTWKTsxjn9pHSLLiXmYfrcHD/bAQcN0Dx
9OIEtCMZKCS9g+TRvtdsM8TBi1lt7vTOAnWvgbVwe3UQt5ER8COUcTjMmtWtgfPB
vR9t/sh6Pw3Opy+QJGBHSuzfcOtmxU+DybJraWbR88ldTQEqaKykLLgbTv4Czlc/
ET1WmHi9qrn5ifUePSSoEitoZhoyKrpqugs0HjCKAkYhspL1D5XwuF9kn9Q4+88Q
nGKWlZ4MUT4OQQHgx6S5PEetrPduMQb4duQH//a40GKJMDvyKdS+WPK9dZk6Jh2J
rC9Xg1esDbl9okmtZHtdBGqphyVr1+mqcau+/auWp3JqQigMAbbp2Zebk52acXJy
9fgK/xLUWDfyU3Tj2+WOn0wX2fUAM2sfMNcuydERIguVXhn6Uimb8rR5lxaOe+jN
nQYvVgy4LyRa7F9iZBidBz1ZML6ql8TljnClTYrskhSoQrndx8nA+GlbROtr6xRt
/BEl9PLWZFsFfm2/O06XngdmJ0+mTdry51yikCr3Pi0GaKj5Ziq/IFS3ce0w+wdO
iEzurBIsL5jfvf5Q0NVN6NvD7gm4ZYqIeH4ULiVEB0Y=
`protect END_PROTECTED
