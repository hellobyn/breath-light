`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwp3HChzJG23VRneOCLz2kBg+a0DPNbE9LyJRfJO3qiN2qiWPzmiA3B4YWUqp96Z
Mep1SD2Bg0GJEav2vq7pd8LtCULNS3vJCRvI9zoU9OO6TjqY1AgZN/vb5aHJhFf1
uWimsKiqp7xRSAS6SlErS/9nuGO3ei8B5hX37KRere7ZenL8m68w0GPrCyJm1Gl8
dmLnuRxODAeJBepfubJL3mvj1WKEDnNMtJS3kTwL/h7SyckpViWLaiKeZNEQrNoI
gLlWuLK6QUrTWaovMd3yzJHtT7h/PMvXK/pttmE0bULJAoHmXETsd9ukiORcvIUe
bIxUFdwNnANQFruyLe9sjRWxo9R2NB7ajI0y1r7KKTaZ7rFSJP5dYtGDNk5lhXe/
RCY05eRlMW+HIiCVbZjmDVGRAekqyYmifVVjjVBv0V+wMWBjlVfNmT4BzDF63D2M
kU7f6fB8etRGY50c0JNmibmqxWXcU/1h0JbFbW/A2fdf6V9PZhwM8FYKNxOjckJm
eWXtoRWFOHAKCg8h0pL9fti3N1jnVfRZazXV6bopktNt000sbJG9bHz2IXAaqdm+
F0rSjQ6V2rxFSNsee6fahs93kMzOQVDL42SkNob/2TqsvbyKDDb1InyUXpkae8RG
AqGpn6XbZMkV49B93CD3/4yhcG0QATKq2Aubzitg+ZIxuJKvrUQ+vuL7TB/vIQSB
kHtjDzSTdkeqI5vf0zsvultqDRTBc+yKwcvDZUqIkvOSPG56FEErAWmjh3w0C0Jt
3b1zhYOdApyGRPAEfk8+xTPUXAnP118GNpwQ9A08ItOHIWERvlwOzKQafyFvLI9z
8GK/gkBx3NihfYWgR+tgQtkUzKqVE+IpWcunKAjA/9cDz7ovTb6iYWmoIGIFHsTl
7bGk6Ma/4PsBFO1ACeupr9DPD70/zfaGMYKfJvieQwFs3JURJnltBw2BCNpllUdN
MPi+wrDxHvQn+KukIj6fhnQtvBRHcvobqggMMEGdMAW2KghKKkWH6aS04ptKs7Sy
KJ8RYr0mdplUR/0nN5js0rbPz6f3tJEKokrg6ZGQP+zP5yeoNb9iaLCz93I5S+ca
vQ6JR2qy8mLQD0YdBWfu2hO2O/7f03vBTfF57lXAy/tXYeyevo6ZZ1K0GWCEffqa
/7FUbQ0T6wf6Tyu54KqyVA074wdgL9HS05cCPSgr9LKRYPxSiaKV5RrLEr1tO5Ez
gVpB+qJJ/ET2+ttQyUeNE9eLAzw8KbHE1JkeBu9an0s6EoiQvAXzLZhp/T75M0HE
2CuQUoGdRP+Wdc2skDVNo+W7R6+AlczwnlHfEMi6M2w1FCpUucd0cuUukdc8qB9w
r5YrXkATBUH3edL+Oi5OnzdUfH4a2mEHBxTHPkya71eeUD+e1VW5mkosdrEOCJbB
UMQguZig+9H37XV6DMjChw==
`protect END_PROTECTED
