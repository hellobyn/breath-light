`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XoHMq4XoZqgr+Cxqmnpxr1hqbZ/xkCRtRO4Nk80eYRwi1mnYOZ+wCc37bwV34XK
PiPRTqujijz7P/AsAvqwKOwhY9FD9WxFnFnNmgyvc+06t/nXtWMQZzgrgGiPEgpI
kMJYg2AeDpcDt0o7LL8HiUT86nfO3fC22nbC0fM6r7PRTrrrsRYXIgaupUxNCnxk
0rSRxNTFNvwvxr1P0wGPDgq12hH0uZW7QPoKc9UALGh2zOj46dJuzj534TxvQpfo
OoHelY3jU9zRHRffhQuErIGOpusF/mpONO+BMGVdjoFJ7nISiul4+fKeDZn+Azi+
Vr6Y4ha14sS3ikhb90HIsZ3m0Y1YY8ph9ydv9Cv+VAaS6VqyH/58188XbyaOHhaW
qjfC46cvamKAykJMSPDG3cCRZG1DjhaQG/Xy1Tq9GnqALpc/zb7fWRcENSNCv1pv
6wCQJzqZXhsnxpBXrAo2idxVL9Rhf4Ro7nsffp1HNJB3OReHJa5RWnRPVH1nOIaT
0ZXfgvZ1WfGlCqVOdN/b/gqFFyw1gTnO9CjcOMLjFnL9FD0tuu4zn1kJfr1llrfC
V0a1sxm7IjUEGm/VyYd4pAEM3SccQHqL1HEgeUmH2/lm+9yzx203xrNIA5F3cOKt
J86fpBkEZMVf/NC0nqcQQBbB818zrEZe8SNJqzLkRAOVaK4Hb4pdyKSG5nvxusPE
12lco/wh51hDTHwusenVNo6NcgZ22So6L58A8yVq8kP355Y+thZU68QPwyUceWsg
FUlR6K/XfRHqs9vPdTRXuG6bMFqe1Jsry+Ha+AIV/Fh6Bivvr91X3PXU356gwPRk
r6vN0dYvaUcsUE2qBtL0jgbrLMORQwdNyy3wBhN2B2dFdIjACpl9HJUluN8Z+Ra+
Ps+o2SYdYo0/tnTINvtYUov7G+d32Dwi6OCk88qZYdMfxYxsGQ1wz38YMDBHkLmj
x/2dnhSuQHlUfokrZJ1TLGdP8QFsV7hapnWLGJm0O1opAP7cZCRhGpTQGNFscYRa
Giv4CfHTtQgrhLQwErlikpJkw9LSRP+e1jDaDHqfZkhJ0wpJDPoNK7wmNEVft5/+
IO2T7JBxetEeHHRT2eJD3H0WmwuUdRZQ1rW/owIhYbZrtseu6sEqRrYJeVL4Inup
pErnZ6titfXQO/ewkxjHICnSMPioJ2obNuo9t8rb5msq2DTPXciz9cO45C/tm/lr
abg8qPSsPd/nZG30UBmGFSX4nrJsUshjSfXNBTia8EGjUm0/TKDUs9C89MkbqBO7
YvGFgxJOy0qLsdAdMpjWiiAIN0unAj+I4cY+wdJ4fvXrMBbYDqqnmyuGU4q2HksK
MXLthcaWaSKGPlrp8gPI+HnmIbpgN6I5poFrxopaVgoX2WZbUK85c4Bk4YT9rANz
fS2DQ/4UJ6Blfv6Qd2+MxAqTWRFq3YMG4AvG35s7qPwDCigb50pjBiIAVPYZ5JfB
`protect END_PROTECTED
