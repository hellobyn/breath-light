`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rujFgnYxNuS0eutosArIoiMlK85bUZzZVxafPgZ+87Oqp/1NEkaBcA7R8P/dth0/
hfvcPw9kD0dNfR9anQFWv7nR4zH3CDAxtBuzU6LEHNy2x2DAl7evAIXFZticmERH
ZJLbakUfh7EmgYxD9Lb6dVpBYhGH2KZRQ4+pdodKEPZZPxMWYaJj/hAb9xb/N9Eh
wOAhsTOmrn7w8wqpYwlxkeB7DstwkX8njhcll4wB64FVP7B4Z3hJ0P/GnqlhvJbP
CCudu8LpwW9W58+evHaPZa52ry/YGod5AW6wCM5blViKk8OPQotMUf7kHgnFAyWI
6GDuUAWve5irRWaGxAvsBpbGCSAWI25hIamtwqO6fpi+Rzo/vqMTH8umbzht4TrL
FkGvo2kZW/Ble40LE2ab92/myFnYLnF00INXEHoRufK3UxMfuC06clfbd1hVXxMx
Vwj1t8/K+hRfC/1No8bRURbC95U1QGtg2/13rnmxDSDpq5VB354+OSHvqwca9kvp
yKSgUIxkva+VoSOReV50J/JD7QiTv9FRqljbLjxt5DHiVPMUF2s1aeVf6p/I+ccw
Qd3pYq1V+DbZoHfdJQSjgGqgFgdcNNYszN71n8KLHAmeLfocxz8WjI5phoOScv3h
2ufMkwpoOthY7Hf/XX9XXthYjw8kKx/aqtPGxJepFTxpxxh03CCZAMLHqpGQ38hM
D4vHe7r6amw3LjRAyq0BXBjxJbAY5cVQhQIgx0c+n4Y=
`protect END_PROTECTED
