`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
giQsw0GKThKEZorf3g89Tgl7Soh6ZKMRY/Aj9muod8/aBAX0HDhrjkKRWnNAf6Vb
jo/UPrsJXNkvot6GZ+7onpYnmaSbgf81ClIgZC/H9t3W0SMeSx/2dajXDQbh3onZ
F/8iXxpZbc6Rp25QTNNRNDXdyr1Vh7CrIaKFj8IaI8DQDIn9k4jpXIYAlptBJg1V
eEowdnSeGsvoj+FqJKqlVa2UZWpr1bYWt8zqbuBylw4dC52iFhKh8+Po1GG5iWP4
VsBgVVtPm6xGic8sChIyucPYBSP/b6ahCS5UXy2JaBiY2Epzj9Xdl+EmkazRDuyn
fYEup1hOXktHTlSQA7t65OjsWsMx+oomEgNrfVY/eN6Eel1SRJgqY+JLXF59e/gz
hZ5xEAdoRXZQAMc7VhtKo5tISNFle5F4u/cd0ewj0tv/OKxGXECiQ7DhfaA+ZRjI
Z01RicNxtvRYI/zz5WfW2jK1hSjHwebRMAk7QbPZxVWnrEZjC/hnacvH+JVg+9+n
`protect END_PROTECTED
