`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRdYlDRPT7fNHpewt02hOWZyHCm9odbLthHZLsgyJyJTwpUSfaFDuH7N3QnGWveW
pGBHpAbdHBxv7zQFquJiEiOPd0eDjHyKcjz/x9ZKaIsQ1lBbIq5e9In4YrEHS/56
Ypq6zq1wPL8TcaECAf4+J48gm5YWz5XxS7n9cMhoEkCucNUV+KaF5jwn2YCqlVk0
yXazkTj4dOI/ULxDFYjlOQ+TGdQtd/M0ToyZGNHhCOZgNGJOR1jWvcWffc2lYe4G
DqquZuKcq6bUkosOkNSmlw9OrrG8qYuNRETk45wtIJIOyk6AVNm++AwckMVITzhE
Tg6zvL8UIsgMruHSOcaGFlHbLIHt78MIbfdbaBTfehadrjGR6l2gWJ3JxMl7aCjs
3Xdm6MRJ1royIMirp2bCZU9S/+EiqbZ3DiGYkEeL17jg5RnO8kXFtYYhlPJ/V8vf
n3YpBLJbmawxGiD6jFRkKjB5J+vvnfYAuRyLg1rgF+Ys8Fyr2BlZ3mkQI0Y1TXUI
cxpxXJoPxR55LiWQHXI7MQ20blgp0NCpOZ0THNV6So5jqlzH5VryPGbW6Ay3bg4z
JPUt7S/mZK67L2RK2EjfvyTWgsAQ+Zu6cqi29J3cfpYrql+DFePR0B+A8U0K6fgn
RWWuezH/SoWG5AoneqaVBmRPH9c57FAJ0u8zU9xi6WdgovTK2St2zd5GkqykNCPe
ZS2FoqdeoGzH07lP1ExgIIj5c3da5+8D83JPYcPIf52aYWGWXCOJ5MDgY5nxAWlR
aKQVEEGN8SPn3fjlTezU6TM8cBHjJxRqyQ6lSXHBplr1PDgo/26X1eA+IUVTp+3p
ga6/ccpOspnOdH17ATFxQd+nkW/R/ccOw5Kqa7zPbtQTyTbZl2s0GpAy1gNFv0vR
kKabdWCPgtgXE56ppti8XtqZPgGDuAPc0m5eQP263vWRMNmfagq3G2Op13NZfCxJ
rQsVYh4SKtHNxo5W3Pwpr+Ys3LZskGFkN3mCQIptojz5ZX1oj2Z4NTgE/S4IQ13c
LNJVf2YxBukOjz6FXmRf4CxrYZYbxWfxWxgAorVcqdngpmV6T0ZUg+GIxmSLRd9G
NxUYG0jcINDJPWwd+SLY1TGYvHgQWYZy9hvv6NC8WTreEpXPJouiPc2bfgOkFLgu
TtzUakYalXO2JIggSpVuAGO4feLK2vc85e98ECZGTvrdemfaLWSUbqhSKurrZcRq
oyttH7ZPWiXMNHprIII+EASKhym3BSsTokFOcYvrd6LRjtSGDiXbz3ZjCPaHtssU
2b8YBLzg7VHOQh9/HGXVzyv/fijYhJfSp8m2iONQwdwdguBolTN+RqRSHbX2n3o9
CT0Oxr5xShJw4J0MNEwHxsg28ssc4FiiasJu8qJdnVCvlr4wdi1z/khcbKUERb4H
qdR/pH4oUIwSRPCcTEKhE+UQ3wivDcVx9uyAaFXmia7uTQFn5k+xUdG5NRRo9+03
YOcKe/pi69RX5RbfH07rLSHorHa2AEVwO6IEeCu/T6RScfbmsm9zx3ETKHDI1OZx
m6b2ZrhVq5lpRfeKp2lu00bTcDclbsAsBmNR+w8c9YrOZz61dpLmTcOo1M7Fad9N
nOouQTdUSKnrmjdHQ6VUDL0qVgmN0gG7CiUkdrmHdlTZVdbvhaQLb3bvHB0pHRhu
Yca/C2TXjiymd6h8TMYX17VVphSdTje98bm2Q/V+PD8yCQ7OFPcPJ895YmuytcYR
+EQC195qReiDMlBxlxEsHk0N4TMqeEVVmZp6DgIIOT4i0hZxefH4NhYP0UaPv//m
aMtWLjZjzpoWuAwB0lw3qoI24T1p9lE3a/Ky2BuwOmUzBs8Bi2YS6C7wr8aVkSgR
5frgfz3Hunuh1bxuNuigZyNGRnCqwshFedg0yT9jBNWVofShrQ8IMR0AFCQQA12s
5TrTFJpZ/OLQVVKi2HApXfGuo75eNwQmoqPqz8Jeq8eqzDviO8SZUwm+chfcozrs
NMAfSTurD/Mn25OXNuQmc01uREFa+kq1Z2uM8oen+3fuKGxTizk3hD1+iq6xK8OQ
kJ+ifP1xKaNdsgPRAWkQ5Q/OD4VLRxpBICzO5v6lI/dN81fYkH0vGQZwpXLJRYKq
oTxKU2BnLNCIDYrM3oltRIZpWQWqW6lB0ApsyxX+NYj6VmOrqP/KykuWnsMNlLXS
HkaWgdVVi70/KOTXy49cfsz0agZi6gdI3L4sBv0z/M7LA0SjnZWxLM6mcBrcoZJU
bx++qdy71+nUOKxImqbggtLkCuwU17R4EsTCuXw3+7pac+UVkAXXjUCpt8bUsAUq
zAONoO7q87jvoQ0YVvPvdO+lUXz5uUwxmUIDb8oQVPsP2wN0epkhEno6pBudbHO1
ZgXEwdW+MCmqEPC/b/ItvD22CX8m7/ZNAFqBVCC/jrGNF9rQ2lSi942mgJQTDJc9
V4M+v/OP12r/jxtUP/z0+51Qu8rZeXSyW5gizhdRZBBxeXbJnUmyaiwP3+amzi+W
C0ssdIGN3E2s1H401jD9mHKpR26D2Q/ADqdjH/yH1Co04Kf8/v3hqnAex156+eUW
Ak3oIzrp0BOMIVXC74o6DHv6eISh5zVLbec647skO5z0F991wliN/fRjkNxVAMp3
jG0o6uZmCbL8SuKNvQiWOiLuNdb8h7rw3LHo0ATqT1I2rPAgvdxMlEkjDgSJukPs
MdzZETdb+75cAJUfPUaI+yvub3Rmd+RTeIt+fuywY85rnDzfvhDKyjBU+9M4547M
pVSRsGLVYzVrvtWen5INljZxnRUCTGEP/Fj6xrkdKdeA5JUgDgxzyy09kQQCqEmj
LaZa9BQP+ja0suD0ZwT3sdlnB9foXak7hfNW20LmM6TcZ4HLbpVZ4Y/Zxr9yVF7h
2+qX0tFfw4Iy1cua+hBXUZVUgXJSBaC4gxX/wO7f2grTGpZLoXEcoFfohDYdBgz4
AxIHmZJrmij5NtLhSvLAMLJSjY1M0C9ZmqpQbLHI/GBesWrStgWMQ73/H4wk7pXi
mWbNM2Vy5VMeC3Pds1EgKdC/zyVrrCNQNvWgRSR/Tmqp2nJWqowqHd9mK19DfVAa
fjzV7F0ELYugmdAdANvN6CheRbgr9a1muSs5XjmD0FKR3vRP30PgKpIpR3mihgjd
BzXibmgz+FuvCB9GPpf54rsBOBV0fz/7pGmoShpwlK923LHsrMEcnP7htiBY92py
PJkenpgrLUxkMq0sgUnj5XUEKvepGcFwVKDxCWdhqtpIUWdRtV6QwC6JE6MYLR4E
mlOBJrLSS1NGOJ9sd9ECrWrQXe+6PosqpA/U7A6nOZtKP3B4eiM5O1WWwZnV7J5M
qX/+CkJgwGQ+pVVoDZUr96klW49/9uC9QWcS35+NU3pZyBn8MgcM2RV4NBJvElOV
9q6zz9bTJ4v3duvmFVxTfd2uh6rkCNKWVR7HUcZ1ijrgKhaigdYZ6yAm/MB3uksP
0ewg9m7nlSrRKLZSG1rlifoNEH4yhGNDqQmHIsv3yo3wBC0RvzXiQ4kFrk39LnAd
wOk69RBcn9YNg6aV5bdC9WocDsACSxpQCBfoDqfhCWUTgEuJP3deXhARErhdHQp0
yW46mW3dPxEXANZW8n167jYqWThX+LeBR0zKtqEDrS7WQkIZywzkbf1nsjfunPKF
egB/STgKY0X9PcAqkXgPBQ+6yzo+uI96cgvdLJbT3ANeoSbTYwALBtO8wXpZZPW3
rhEJJfOuCm0e59skZHAEGRZw7esxklp+6pooP+ESKvhMMIvP3+eHuqziXq9e+D8h
oGkPgix7tqoNaCRiAhozv/68gYe80aDsSc6Qr6rJlgSBVhz4sJT4Mt7XiZgXFH50
XVHCwQ6+mGSTyHuMsNOqfgPczg9Ghgc+KIW9ae0agJB2JeO1A1k24r4ErJBYeCBm
BHt+0dqkWgxzQMO0hrOZWB5OuWynXNLNBov8yGJlEw4mLx+s9eOI5ZMOCMQKVEng
HhNk5JluGWn0ugu0y+VP9m4g392sZUPyNmnZZ4GsFvG3Xl+aQ0cOKWvNY0Kwm/JG
6svE17xrJC0/rWsjIpJq51+IhT/IssXWfp2T6vftnn9mQXdAnAF44E3/RK9Vnco4
kC0Jn3NBUZxKpYkppM8YWP3rLCm/86hZCQt/+qKCyHhLNfdULlmls0r33JLfANJa
wNRcCabB3Poreyq1c9x7ICLBFJILavoodbDLMHMBN9/5ta5+Dsidb3c07Gqgwaa/
uSdkA+vVQyD4217wlO5Qz7+P83MZhFJxAvDZYbK3cd3TQTsUch1kH8uKnBwOxlmi
tugT539CryPv+HX6SRfsNgUQ2ktOiqSFWYxDxQnR2DRUKPSUJO1ceClhAtkpW7nv
cadH0ZQAFORuii4lu8CzfajNS5pMPR6iyJzkJggwmKjcSeK5ocYHtpIvP1JDk+jm
jWRD/vAEpwYAAfMQBp8KDW8OWpBUPaC9hcky77YLeooALbt2qAI9fdI6pRWwvkRK
YWOsWxjTq1Tt97v+Vm+n7JABMkDqdcN2cP1moJOnx0uAZrLwBdeMRpuSUyY5DLnm
TmJ+uQlbIX0NZ5HimBoVl9c+Qh86sP4CHK/Ro38RsZcgdiQkyXDb/69n+UHvEg9N
hYcotmwY5kqT652O32IPlDA3NpUUWsYbdi5pCSiM2c7hHTMfXl0Hg/bxT4NiMSLd
swhILCmfzczcjxhLqAmmWqAmsQl1Yk6OM1kD7d86arrsTcfHkMjxhuSVFyoz6F/L
JwZODIWEfj3T/Ao+5VVwVWLPgzbDD5UUDHaQ/9Fh8jE8Pzv3PbZ1iSZv50Om9uhG
AfTkPXLbXEIzUgdLmLDrgr3tTx22T7SzxlIx73LsPJJ6mxgYGfswgJjrKMHURkfR
EFjIMv+/8PnblAO6Ey4JFt4iwKyKy4A1MndIUwjVOwbb6HMkNUW+xZMdxrWVE8/2
ByVeYDD04dCqZhO5p/VbU1bLVVLJoSMUcHUsl8DbrtNvrmjCabIWuO45VRZ30ABb
gcg8Ua+IiPQ6p215E7100LfvmbqpYtenfuEGudXJItYPOwmv3vHIsIfSL7yJDxRH
mIO66pp1sPYFRF3cX/cnXFQXkHa6en0vBkdsBUuyG3k02mi/fGvZsIq6JgziUeFq
jUBv3p4YyvWsG2t6V46PZkRbKoDjfoJMpqgSuyggUSts9ZLEQsumhvrV/C4Wyydv
CayMLkg8D0RRdBYAwfuLnF9rkJgjEPwyGHydeQeoWJ+3p/YdoQWnOxW+/PNHU64U
xO16kf0D5RpF7qVtpGZlzAlA85N5DWAnp+mRH96J96qR6VjIZFm3b0cbmtZ4ddWq
SARSV3CppZWOtpVS32rNqx8qalrGzd648nRJZ9jh5nVyRnqjk/tzPY0u9O13NIve
vllwpqHYc363paleNAXKu5RliRAGSgvrMGKs6eOLVpBgLCcCbUMfTZxuuS2Uu1gR
AvXfXkrmANrjtYEEaPIBzXcIlFY/PhgV/gwQY/zPqN6rZNV+WnlvTSJQsNS5hGBM
Ji1NWPXeSwMAw2c5ng64YCzHoOnw1Qh86eSvqqwXPTbLgC69oQfNlrTFhMQn6kbE
yvOqNbjJ3Px9+kjahtvNjiO5oQlG6A8AaMdkQ/klDZPGr+noQoYGC14Hk9Szw1zy
7PyZrrP9FtowUUVksYzv1ysx9RFMeAK/WV1Rq50qUGteWnq4/GIraTjQ99WRT6+u
C/kgLhljgrA8N5VF7m4rsKZYwgQuXnKoSBtaqfs3U/g6xQUehPgRwp5zQuvQgvGH
Q2TJKJmseler74KtRqE92aKdQkPuPbiM/Qw2Pw1tupK5/qXilx3Wzn5j/TPgk8Ii
udwkvtUpU3Mlr1l0+ZTHEqw8mzvnY9o8qa7hTDnwGmUdTumLcbkuvemzp4jOmDm0
Uq5fc/FrR1NnGmi98lZF8cfzSnBD//y7DcPKO4ksMNcUgop9wxqgcTPZmlXSPpew
wIxk1Kd/CJb8x/XYTEhTaPEYjo3RtSC3cCOvPSfKCoywWGi/b0P3rD4ivtMKrU1Z
jZITkxlskF76Hsc2yRiMzYE6YR9m4CvdUnJUUHIife/7pzCqjEFv69wYgglW6ZYP
xLubNTQ2ryVYsMyPBD6BQYqcOdL7gk9w2Hn5FrzGylBlBt4y35jzdni0o4zBwWoy
Q5NPXJY4YmaOJ9vcevhbAzpHnaA9K4rM/dRegs2Z16y0n1NB69EFXC1KUZiUcFEN
dbpw//4PxE4g13AwKLe7P0ajmM0eZ07kwou+kicc4qA=
`protect END_PROTECTED
