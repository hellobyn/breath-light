`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R/8rSLLhtrFESEYfwjytUhRD5cvCMSmyKHrkFKnpKgA8BfgSbomoZRvFSNAarUsV
z95CoAILhiY7omfHQjQs6+OFEyQOFHWoMiC9+oBCk4CS+/qFE4sCTdwlUrrJpkjj
SBDuCV//XIyoe73sWpEEFlZ712G7KYAXR0NyfbZuZ5wcZn8na9FaLX+K6UWq1BiP
lnez5ZqJsPSlOSTBOdPZnglltA9H7S4PKjfSxeh1UcfwjUswtQitUfR5HdK0oQsk
E3VVD6ecejjq1PX8Z6tye75fdg/gOjgcu/KG9vb9/Y0BtLuVtQqNEZFa06yfadPH
UNpMQk2CdJZg8gQashwm1uOIOLw9DJuMGmwYqAwoTWd72BZg2MDOtgxKJVJ6WcDh
`protect END_PROTECTED
