`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HavTW7ZTzkADYV743g+5htuOY1MNwv3FcMIr53w5CB3qQRJNlZYNfkGAVl0RPmTe
9S3XnKMpLAFeNyWfF82cdzTv+Ksy6CYoDqCy907HsWlFFQz71+GJo2+KQyxwJpEV
dRnNevAtgx4vLF2YWOwa/Ze3q75ZeypC5QFnCaqmgHdCwZoTd/mQYz+wu0baflLF
MVSI73dqcIZ9mePK8Pip+xsFegY/zrdI3iE+i7o62+m8xFbSKBvS3+GLQFkeweQz
b6tJmnuXri7aIGrLX9p2YeH+3aYOEOBnKCbfWVPtWZkQY8SWrxDiJv5/zGVdgcy8
XguLbXyGZnj8gOQS9K2obt5ialkS3HY0usH/5ZR/3GcSgaRjU8mqu4Tzrlwpvm7v
+I5Avwdzoi5J0U9+H9PUysJ3pFVbG5h5fyDuNtGbo/9K856garqyUkj5rgNVkkXK
JqqnJwdjN4VfxWaWuI58xJc1rDRHYIGYaJtaQl6eTdsS5d7ODw1j86dNIIGiaIBD
D1Cb1X0fjf2cgINi/J3yt46C7v6YQAObH62xSY52x9QewbyDeoeABfNb931K31H7
YqPNa8YjmaULbR/lxIC/rRvSKwSGTzjOGIlvoUuJC26UjrbdQ8qBOPykJ5vkafiG
w2tAUUxjkRExfZzZK+pLzG0MpVs2xoSdiIcLLbK4KjwJ/1cMNpW8WT5/kHv1MWSv
FdqglsRTOXl8c+NSiiL+qzZi3+MEypP5tYx8Cyo82a/+LGMa/CSu+gCjP1NXpHN3
Si/gm9QEKIJwz7dbETH0aW8YOt4Hirul1nD24ZScVxHfoi7LX/Yu6fFObXshqGwF
Y4a1EXLDUvMAg3a3i+D957EVVoamZtbEngenqALZOq4=
`protect END_PROTECTED
