`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gr5plOAUvWmAIHVGHBx7ojjFkvNOhYmVpPAdqmpwUMtdBrYyXR7DWN2DAI99vHN1
WMdkqclN/3Y0+GlOE3v80uKKb+T74CUrgmuJBeb1GinJTM5CJpQLM4b4KEg05L+K
TLUPPuWLpukpq+PnRYJLoQWpnLrd19i6OpzYuZ1fMyQwxN6YsowdUyZyoh1x9DKt
LwcQHxlmQ+bESqL0SUIvUcaJlhyaVha34bt0WfDhLOAVy1/5e5zu7gjMRjRrYxJB
dd+/1Q+WE0Nhng+oB4uMCgQec1ExoHTP6qKSTdwnL8bLH6SjOuHx8+570KTAwk5P
FOqeB31mNzdSmECZNOaeg/E2IUzfQSlGGzH3tM/2bjaBw7+qgn3fBQoSijJDsBGl
BvsUn+gFHOtH0dCXx4Ci8wetUtrqsHTOijEqdMNPXXVtV1v72amQze+G24wol2K9
jbtiZ5Ke0rpMNQCeNw7tGW41XfWnT5niTx0BYyQIKu/M2qt5Nai6lItP/9bsL8t9
IDpG2VZmwdhBtPpKwOId9+V0avBl7Q0XUdL+0o9SP+bF2mrjHGuZZsYdGrZy0Qcu
qvSgJgNqXgoE/3FG2G45AX9zjCdfKXW7AP4N7XucWSWmYR+HeiTiz1lLi3DaLS6u
fUHXDgJJzuh3gQrL7btJrElhfhUtZPNaGH8Cz1VixC0ZYRp8oHLdGKz0a6S2NsP9
dS3TgGxDpzXyM5oXU/Ds+w8b174dRHP0ZKMV6eLUTR1yjfjfYq4zFjoV63EmA1xC
ZDOuLmLTCRaI4KLRuT6eh4PjESt3wph5DU+zBHspzcnvdlniWu9eJn+ErC/96jjK
pqozrVM8sUhwUbq4XIWFDBDu9OIwqPMhphItqw0ofLUFjNE3WIWp1CmirZQZxchS
VqMF6MZgud+i0WOaY0aqwMnvYmKuGeBmn2K48Sw+vKuc3M1AUl8RBPjHRldf6HJJ
YWGLpKWg5+AJXyyF17y39Zv7ITBzMN4u4aFI0aRhFZY=
`protect END_PROTECTED
