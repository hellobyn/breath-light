`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aeiDujNR5XSGSlhj3DHFFM/gSBv8/s7n7aAfWdqDg9HNsNdtJoO6QAG6Cy/Ux7ZN
6mP7F8Oa5DN70dMtof0a0gH88zWwoIUpXBA5Y8wdsdUvE7R8Ya0LrqfhqiUxmhmd
LYQ3tbF7xX845LglU4BwMbVtZ+qLu/WEiKotRChOzjnaCQFhxiG/IwQNkv4EzPIY
JCXOaSMIhJuxkUuyP7uYfQg6jFN1JAX3pwsw+zVH1Vxw2SGJ/q/DmbFL1D71sQ1G
RWXdQcrPhZsb8h9HwLOmNRJWvCvdHfCkfixLIswkeaymz6bOkWk5kIx9WaEv5NWr
LSGrmZSTM7mnxzQ3kvQ1+R+UlTDksIxoK58nS9QuWGgfNnJAeVuRxaAqtKg2qyrH
`protect END_PROTECTED
