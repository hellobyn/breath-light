`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qyz43LrE4yyuh66SrillWRFB4DSEqjtlltkVGCebQ3LZvtBRd4UndCPjgfeu4Qj
85wHDCu3kqUF0hv7nurL5CgFWNkuHbd9xBDj8q9OiIALZz5rhimRxvwYAibMCDW2
0BxsmR/WJHJ4cvUHZdWgU1FlEN3OXlA4TXJer+plWpOMK56/MMldH5TLcRwKHLdu
mN5a3q9BqWyZLg0BWJVmktDhby09HY3vzGzwVamQ3XINKfSHxwDAWiMlDoO2CZ5E
bGqjCi9QhHHLTE1DQIPHatRvEwk8yMlEC9sxlaHuUVF1DPsRkBCEhx/ybaD0+XJD
JpV/db7E6aq1/atbxHK6xmqoUp1ansqpwIDAW9hcjWEv4cBlzjsbkTCibOsuwQ+Z
dxuvb0WGo4D5y2yqqTJmRTnKFjQ++bulyN2ABQN6D6cPCBywwsfRtijn1cJUeyTQ
aDiqcA/zzrxBH1ydMpexEIR9X1uPPnhcaBlldMpU7+3gFalepgR0OFBS+9eDpIW8
B1JUacPh1nfXaHIHW6CKDOrP/4aktMD3d8azbiGI+8iEdcFdraDJbNodaOjEOieA
SmwDh7YOqOVv17qBorefe09bt1w2JcZsVvPBCItFYLUWohohpbOJtglnvtb2ziif
ecl/UEbmVEGX7d4Fd2A7fQX4aa827q+qJyOunvS412j/fuI5HLdPEfXspruUtiIb
tKerOvx52VsF0psbMQ6LYCva0AwQoYedM1oU6Qx5fPuCJJUUccUe092R5QidQrD+
eEuP+zfbDT/BGB71EUcyq5ZnpFohP5FeWvA3Pi50QXAPf9Nxaj91PQbfSokNEgFE
HWzxsm+fsqYRgP/YCNOsQ/7rvOfbnWWLZrrYDILSQSaAbQa5ra/64MR4kwGGdFZO
9arhiCw36DYONeIldhrItA9QW1DNDYzYoKvpu9Rm0FOwxHf/qHMNikRjePKBD/rh
Qx5xjgaqmM1DDgADZOj8tEPzbhwn8sYLT0M/z6WGaclGLz6vklcU/+v6cbe47klk
oma6zvEaumT/DJ9bvWQzi6trfb+glSMHAqUJlhw7lZjyxT9AiZPI/iY7KHUbUa2B
cMcsKm4Gi1tomlsYrax1oxseZEnttS1xLqmC9MQd2555EgeJBjzwOo1cNO/QCci0
xK+uEOVTKhEsXsiWa25Wf8gP7BB78nSvGs+fahL7R4vjOp7EXfRPWEPbh78tZDGs
wJmR1TOAMZy/ebPaxMIs1s3P4dhASYpu1p8D3IEk8T3TMNkuFbaYn5tBHwsTQiQv
dhpcHEjtE9NeN07vEcDfCXg4e2Zn5BPJU2OMupbzviwKPFf+OOX7IRtCpXGweDNw
OpFka0aRsZ2ouXwMsG6GcVUAbzjuBF4n0eR+s6RC74e6budERpDz5j59/WbB0S7C
Q/HL8DaJ4PJx2+rv9VGiOgrbqNOhkH2rvumzx+sXvoHJbzTdnhvyslcwJgXtWVyA
1pU3q+a95VT5GvzvKerQIQHVcsnO9kD6hv3s/fKulKBjz5teaHMxKzgn+Z+Dj79N
wPq5rMyGCiXTXUCwJSPaF/F/xOQ2x4x3D7Po2p51iKgSISh0GU42NoYnUQnMMl/T
SJFJiVAgYI8YcokS32LpptBAG2Vm/H5X0/mrD4On92Jwb+0fygZ8Skpw+N912x73
fVsSmN18yuAkiGCEe+YCIaLKMj7Jhf7qEzpGMNzoIcgSKGm0YxKtA84o+RpZF9gY
VLYJRnWS167/QSs7gNnWIgLVI38YHx0FuHWUOybtaNrc+yEBgOe0/LZ4JsUg23dU
oNL7tt4ysJpBVyir8WYGeil7l5BE4ZO3XgAsba8rA0Ax/C83IXf+uZxdHWl68xM6
WTohelij0rPMR1177Rz3rwoVstLTD9knQma556bj81In8Ai3Jr/3UtLRfALO5zGE
M1nlEPABxK0KPgQw82zUIHM2o1UbdDUnGBuaufZqOJF60JaCUrdvlrOIGXl65XRG
oVsLbMLEkXKL6YJxNlNS7lrchdYmVC1nnkLO+75Qio9EBSSasayMberxBlBY5bIH
JpozsinWvUgDmemRlbThgD+xUvJKq9TqSjD4hBDfNYW1rOBzx6rvxic7E029DvHI
UnwTGOQku1q2uxszWPUUsjHoSVEXNk7Z7fOtF+T0rcf66k+rChwlskv0t7kpMH+e
WKz5MhLUMkrCBqli5FVovqPPqk6SysUjuCTSEho58TtQSxVvVI8khYVCk4z+gILy
JxsyPDbjOmo7fEcL2SoLvKIaE4Vwfl6IWTc3WzXPza56awpbzakNYz6pRkaeSrY/
g+dgE7vm97dhUD9N64fqii72qgDtebGov6Y2/PiVbnRP77qBplMk1FeZDF5WQOnd
O48tqlFQ5x2JarafOJ4Dlh1zKxRv/ua9TgO6Ydy+E3EBo3QwfG+lEmBoS1xY9Qbv
On0TDWkySxQSzfOnPNdIHARJ8kvPGsetyWWCx9OmGWQVNW0VRMuWqetSiK+bSLF7
Nao+3Rr1SWBiG2uCR8vdj7T0aLmU8X4Kg6IxYe0V0kPEbM+xvp7VybK5ZjkHZtxC
ScaexszzwyjxonZDuFsRS6nj6Ver2Och6CvrtMlrd5Uq6F5ynfDtEuSmrSom8sD8
Xul3xoTgDc0WfrBIc9tixn5TpqymmmBoPzNOBMbNob03bydWrvhA2ry91rjNLQ3w
SRvKKoilpgG/cgrCkewbHw==
`protect END_PROTECTED
