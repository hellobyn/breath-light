`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCVoDtBHD8LnBuqiLxIkzj98KsdV7RNSkWPnq8rzCrSOejXMNWNIhi7XaxLjKBq2
wk0jV746xKC7NcfB1yajoMJdYquj/w10zUlpko+yG5Uw1ESaI5CMaTjGB7ZwEg+l
7jwms2ozjfljQytWdxTVbRZ2r2PwpJjPhl0A/itu9xDcA3IcScw9XDzkm6ns/7Xa
eUdCxBRrIZI3vSvwiUJbShBLtfnuDSl2xyw0Jo9xFueAV0Gk2RpdmuEtb5udpEce
MnDJ8mQlLPgwJ5R0kRUBz9BbftlKWGg0zUqmNGLwSG66rPHthkT3vlI6Y/oxHG0k
wGsqcuv5M6O+18+q7XxaWjKuHv4uebJDfoagUlXNpJmrq+Vi6wAWxo0sewJSC2p5
ydEtoe9IgnogU33Ja/a6JmuBJeKBt8/M1rJrw1gM6F3ZQ8w6CexqY1kB3Gbj8xSk
GrXQ3MRo9xTcW8fsAST6kJfjopi1jFXtKN5BDKRE3lTzgUrSSAuH82ZR15OkVvwC
uX7uP1xpREvHrpuV6Yvh34z6hI4tEOfzh7LWFjnL7ksl5QkwGMSS0s/ZyKZs2kzI
aWfMKGABM6f9xjEhgyoFqmPHfND+TYc3zAiBByoyXxMeOyh7msZ3QF0dVjaoYoYA
ZqKO9hBWEgou8qn28HJ+7rzAy4+Lv7KC9OIzEbkKW0Q6V0oQ0NGLZdyBRZlyW3mr
0BhUSmxeL1Gtt3bVPl78PO21DFYFVELNMBbMvZcZjttbW/X3Dlrcu6heKTyZOy2R
HAjiAa9JM/1puagEQLLyszbWOFJ4ycrLTG32EIQreIJ+72n0NM0e9KizmAe9sJGC
BEw/6XhGgGF6ddMxRvvOpO4VG/zNoWjuHUllHNdkjBS+Rg4K0QN6CgV7ox1Jiit3
GJ6Mh8zZv8B4Kf7vHdJA9WltziVNqqTcj2qhb04Vorlh37sDFe7+t2XU6/UCuAof
r8CAWr9MIoWRKCJ5rFOBZOjFvBwH8bhHgFcbhG7HgRgDhfYHlLhP0RMFvpMbb5jU
k04r+du6tE8nZEg/l6EGGfvW7OhxrasPJKNl+3yJ4faNTMJaApx9kuvETeZrTDsT
ArdTk9HvGVbbBBrGwKZkIsvxM1+8ZJegq5bwi26Rzl69OlpLqFqAX+y05TgxGPgn
fXroutEGWYBNdJOHl5yY0rZqBJrDIsBSSNIUpJRtL8++wzhdGOw6vXwmxzXDwQLL
TcENRnisHHyPNjVLVn3V+Gv/EoPkIsJUXrK8yXl2G4M+JuNBFxoSbu07StT251mj
D0Uxpvakx0YTvMFOFOC1f3MgxMfFcDTLelzq5fBQvp0O1KfK+YaGfoixjy9dIsUu
k7KOeKhHcL+LRYRTZtkHwAV/W64nzlLcW3Dgr7XkdjsI919iDsytpb1cnVvSc5nG
j7g35aHpz7PEw/ffMOnRMArzjw+rkNrwvVoTqlQCInUiVnsduCCVRBzMi1kXjWb/
JvJyCnXEJ+P38OpTgzyZV9SQUAADRZdXY3WPNSTRy9urZwxyQusabevehKiPuPUB
H0ketls8GiAou40TjWjSvKEwBqKEpwV/H8a84FK694+nxxOppns/V7FX5uvOZoNO
TW8VlytOc73NGXugO/tN/QqArAWd7CaB/xpPg10ccYeFA/yG391ZmXjWUTJpB6J2
SQ8FmfZiDftjK5gou2j2XpNgk7TgmzFOcnqyF6UaDfijuQYJcn+XJHE2Fa65jTlE
WBQqiBMAGAI262Y1U0s3wfMWx8Y6jL7c88T8S996hwM7JBn5gP9r+qunDPbk4UFz
fR6WIRRdn9S6LQYmyKp1XQeImfAiBlnVUVCK2DdhYp8wNeqyPf5fkoL7u4/+xt7Q
vJAFTf5BIpgORjyUfVRmA8YsMbfQjcmSxrirVj0XQp7s2sZSL8I+af+Is+PbByfi
GPnLLku60vRZkDZdYTSLh+I0/87mlpDtaqIyz88BUAkth52iO++C+Os/Pzvwosar
eXyZftlT6L2d39WIx47HiXIsFDz86c5caGBL0MAPsWrUrMtk88kQulHL8lKd1hgF
h3n578PDqgHtz5BmKQ9O3rth5z2VLSrSXFA0EeupBfCRJmpnfox5Me90rmIZSWkM
LOj8+oCZzyVld2O/rrNLTzQkgwh8sw2RTb22+L2zqcOCSxRMx+4P3etfPTKz9XIj
AqS8g3igjyZaYqhGLLgmXXXXiPTBVS45B1mCRKF+j5Tia5qNqQc5X8OkmL7lddon
TozwI3leMDQc/YUcA9EQYHlaDxDl+HXQUsMvLBPXCH5Fp2QkNTz/1Jl4TZKnahLw
WcqExsdNzaQUxsqalDNGUleXtbnLg6sUS33J4/XqBqDjrhqpuYH3Fm7g7y4SE+6o
hcqEgSMVGCVg20VO8SyBDYvQZ2NyQkVRmllLbIqmqXQfPBEjJNTpRt4TYWvuFj56
wrWLN6ATX1I6hdGvh7FrPzGH/hIXWPEIszcSTVNKRHYRhL6S9nl6Nrxw2LKZm+pU
XMz7Um50CxqgP4IUCnjSkankhvnQ/R8TPkKt7vESUJsVGuCr9PaGoq9p83LoPrpH
nn0xqKWZCyv2cte35RfYzsNIDfhYqg80yqCeLplJsQrYdFHZU+EqsXzuBiOQvtrd
qJskoQlGJWF8bPyzl9QCqgc+jLBFRG09NbozGCvIPUx4n4r4YVp1u1bXqvF1Vu7H
oYDYH+m2z1XLQvqNLQzTL20Ahs8L15ifFO4u3lB/TyeUtNxj2s6Crc85/Me9PJi9
8t7Ugnk8A1hU0bJnOMItLCrG05cWAouBGmN4fgqXFheBNm1lirlu66Vdv5QHEu9x
oJICkS8l3oKTY4QL0gUMzqm2cZ9UxQhwbNNPuOP3vSLljCWatFniidZGKsEwscto
c5Dd/Jpdenqmp7wtFlfO3ExfjjwB4vSDcWHpqvCyQFbnHI2CQC9BIlGvdHqzFgIo
KVvl9mjGckYDeK4US0s+QInQmVcejnhwXiCVK3ie05sGLPeHCIJv6OZoYZNPbW8J
MsNlm63nlgtOhEyXWTkB5cIgNLLnJr4RZGzGExmB+Escel6B+unnlMWExLFU4zmW
CfZzSZ8k1Rm6SaLDFovP5985HJZrllYsB7+NSjZy7QN5aBG31pHH6h0l0MCrSarG
x1caB24hkJAsuh+vcoji9rHSbVgzBWhFtgKxRt2MFDFG8wBq3dRxYNRa/BB3VUIA
pUmVoIUV053PGQ5QMvGc2oEU7LO2SfrHTc1VnAcYLwXb5uYjXTcFkia709boeayQ
nhPY5P5C2vzumAqwTab0hezC/8v30yUX1InrXC6UPjOx2Tnex3M8YyUhrKwwULlX
UGmE6px2Kd947Zi24GomP9jjHLzXy/hfPI8rtmgJXbsZNTksZrEc97WsOwoN+iHs
5Ty/rTYRaxpHlk8MWm3Z7/YAA9ZwcuJPIburq1D63EPXm7ldKWQn6kmYj/lv9pT/
hRZpbc2J1zZn2XcY/lm+JyfWemy5UghnMaf7HuMMIuZCMX++SVBadw++pu/Ay5OX
A0sm4r62yvEJOLx7CxRpyWlGNgF9zG+qXJbJ1yTYUzJNNJ/PBL3B94J+t9w+9VlC
ITQ+xIaP5C2Ai5/tRfIBZ+G3XTLfwakSBnwZQ3BzAAuS4cB2yUh2Toy3ubmqk+0U
bxiQVRx3asTk9/mCLW2WXyEXI83j9zj4wA9nYARRM0Pl8uaJOXJw0r8MwYtrYMgC
54QQ51UiBqhPYCVMSZJXlwMhZRKPBG/KFqyjpE32vPDNa4quU17COHZGCDhP5xpL
fSxMsUNbuOoDZ6iHHNxqvxUhWqlZThjmxhmHXUMcmmdMevm4oqinXisLi9eCTSwN
RMNwVsI5zUaycXkMLZZH6qW7Q0VwHHOeA6TzomJ85prLgENSxy11fzbTVw2XWjFS
ofNK6zAfqM4/AOmckDt4k8sLvyXQVzTm4eICH9IZImQLcvvqqCRnLZ2XamAz0P3p
Dy56PU+ELFl/DFNz947dW6GWFqVyEwN/csfyKCUfXZZxlu50lSN8zoJvUZsDckox
czRFiT0FCw43gR0JkWZdA9dzz7v6EfN7x4Omp2SS8Ki0gmB1166DRsLAPBXO6+6M
3uhRPJ5kEozX4who3UGSjlZplnKcj+cxddsAIbekqhEZVe5KPGZmEPzggbcil4f0
ytq4xGCyDYmHSDBtz6bdylfpvo6TTH4NmuWGgwbCX/uo/43EVDPG/yZ/CbqS+V+q
USKrRXB4AQ7KVzBX/JrdYM2X0qvTmXlwfT3JX+MPXqIJdqQYLne2S2vqVdRyFRL5
c5EAo2hfDKw4sy7Qy2DX9+51+jhOvjadDpvk3QCqNYsbyz1pipsae9Vom6mX5J26
dhwqcNiZlhaTpxcl8+ErAs6t38UYnuBEgyCDE4Mx9s3HGknMbFMJFjE1RcPreyXU
e2y3hox5KqbO7y7pJhmuGibOu0Jvwqh7hqH2Tmvih33RM5a0ajCt4CMU+6p0o2VF
QWclaPBtbtIK4yln9pkj/ynWrOXFdsOQo/ODVb0vEN7NbJdlT2SG2gL8SpbOz3/8
aPg0oqHQmH0jT1LPyq1Eef+VW7U0ojm66sDthmArDoxUwdXBm+ciNZ0rmpioo4vZ
bDeKO3YKQbCxO7z8FyzX5CKGC5pX7q4SD+4eY7fOStWe6qFHU5pvd5C8Hh24oqH1
xVAL3yEZKQArDniR0Kj5JRKVfOi3NlcpWgmBhj28qsMELxjuJ8S4GghpHbS9Jd/A
/DLyoiOvmaDgXdqIOPB2lZI2kAdAXwIO/YfsCVOcFM56lxBHXaNdHx2XcdELymM1
WLYhqut2qH5wwfFa2cXhBiAHhT4CbQ9EPPSNDTHcoDSIGabrrag+bV5Q9RmY5Cv+
guKsOEChggfFwXMcktwVDpM9j8x3kzXXJ/uWBfGFxtza+iWk4nd7AIq6EWcLatqd
V0t6xlyZFD7fagIR1NoRnxvgeCrH7aCpZDTWwcOxWpqWkn8FeOGOE9TE+pvo9hgk
p3m5WD4P3vjsEAZxP8pUb7pfcuSkVzdFwgg+zXN7Hjc4sAwxTb9N+slu8YWd+Sjy
vK9Vs8Nsk2GQ9Ez9OXmZ/vpRcH+NlBgBG9kka6/FT1w8Fz/UOBaZHETLuII6yoya
1oUJqWt6uazbRgv5jZxsVAYNBC6l5cKTtIGqF9s5fYT7pNCLUPAfg0N1M1SZ2d4G
j0gHnzhk/0tjJ7eYLYXJgi/sb0akf6IMRMLlOsQd4ll446vM9vL88g43LjlzdXzr
yXIRnGoyFwS6i8VPtUqrf/B/AZO3hnJ7wrwkWLCxkcb+iL+sqI72hccw5mRBjxRU
oRgoXDZw3Mo4P9r2NyZALMabhtpNmoJ4k6tAO9JW3GjLj5ysVb0aBC9etUtGWJJ2
dTVYl40zYRDdm4RSpTqMnzOFNxYGEevLtcT+U/hzS5kPFCjdEuJrAefnMb1ecQ3K
Lgl2QxWiSYDdfbBcJ/xEmjEgQA++yQ1F6wTBAVyenBZKnhLKg/JNxwMicrRQ68Ru
gXj9pZw1Stf2BU01lrFzEM6jh5ZDsHDeQfobiS6P25xmK2zJTzadchyjJwKVFSeu
MmN0F3uSYBJJxuJQKbojtQCiYrzU59mfG5JT+vu/vBUk9yGA1prZY/w32+GxXk/s
Em2BSgz4/eM0g65hGY1kLv/CwyGH+sDMjGoPY4Stym5hk+lfDhrnYlY/53iAcJAX
RYRudLp9wTbSpdgOSTUOmQHEJ1Np2AvNNj7zQZBXTy3UL2LmjKmiTgK6apg6ZJes
rN/+5y7Ff3+tMc4v+X4EMhsqQHFZ+17EtfnL9AAVZT9uJCFZ9BXP77Q5RH1cCvGc
CZN5p+AcH4kjdH+TrJ1SaXHh8dY3KnFiAJNF5cDrM19Ab8UzditaUP8eePGDR5K4
Ta2i9kR+GK3UzGWT+gzOUcurRkxVDxA1xkAJ2uSpWnfpZaaRQ1BOxWobjuGcECg8
jT/oGnHe0vdAgbIjb3kmWO86LP/aGE4iCCKEVVrkpRYna3uaKRMEBccWzYAw6wvr
6VOkEOEqPj6qEW8/bldZ+6ema04OWa0A7FuM7WO8P2M+F/wivEHsCoqQEsvdxJEm
PoscEMGLOWQ4DgYCh8ILmDcbU1GcSaWFjyrY8vDnWAuD/tBwoX+SdlFSJfmWap0Z
CqATsY7AQ57D/f+5Madx5UgjuttDWGOIqT0sh9BR/k4eDcop0k+qnd9U3qsQwYEv
71oN0q9coHodIbQxj0BMAGbAyw3pI2ovZ2Yr2ggNtHL8ynXVEqMrxELFXiLIqbO3
8j+uLNDDzNkmF3x45bKILH0KR/9q2zQfb/ODMbQc8SGRoueERZJk0573lIV7MgsT
DwQFgA74obsR86BH69wvOYNCV/5PyjpDykGmWiXtBbh3YNr7ir7tD7n9py6GjifI
k3SelABlJp8Bj/3USpoTM0YQg2V36sW5BAWVE4Gi/LZIUQ1FHfbdLdeVG50Z4WZq
6vw5sQMNVXs52zer7w69Vs3CZldjSPHja/oFv71vNxGzARCR2mTx1Lp9KnZ8nNhG
RmHhO9XVnSsTyE56BS+nwnAX2vIzPkQyMa0DMuVNqjqlHu6i7lkkvfD+3xNmJWN6
akIucGCze4hDY88vMdsLcnTfHBQ2tUX68FvLCMhvSGiBhQsGPzBJKzvQuI22gQ0u
1Osf3pqMMy8VVsMkoYHe/paUYAGCMK/j3AOo0IiNRKacG74ACZquc3xAEBOfHzMi
BRWMLMcAoa9PIA+O031BIbZYJnU/bZAb4qrmTG5L43/XSmJS/+NoR9+ppOBhnoVI
pexLZTJfZ9am+9uZ6ewFpikdGucuHRZN6am+b5iGdoqCMFT3OiwHDgwlwOKwoKk7
40KGiv3A6u2wJ2lSFuofHOUwz7Fq0dMFocVKq68zfxIkL4hFpnM9zLQr9086WjKT
cf8rYDPrfQFJlkADQ7dLZ/82jCpAuwK9YlUIcAQJKaCt8jtPoIKWHmrS2zeZd6ys
6fTzqlNeXwzw2Sm9mmmM24J3GZk9lsi/VJw08JauQpPm4Lb1LFKs9d9Prl//ru4Z
dUjBE6KNHfVohWoe/XNG+VxFKr/rNfJ4LH6qF5uDD1Rvvy0+g21othFnC704ebeu
xX3l1pv6bF7iDiSTNhfr9jfHZscEvZSiu8a38STe6nOU0+uoZpEc7PEluCWflTnU
w3kEnRZdDBHwFVuaVrGepAjhhJNk4txzvSEnyK+LlQ39Yy4lKQ/QPe1ew9vqQ+dc
WlxmPZMSBjhL9JGXtXQ4RSN0J5zrBT/e6P2KVH6Hx5b3KraMF4wev24fDzCi0zdY
Mw+C6URAis3WRJekV3EILX1n8wYA7t04tsQKIp4qnhDYphQUcDTOuvLx06y5/99Z
XTF4nVtjYILMmKuYgDaNWMUzu2vCurjno/wpbtHb85C6lAFi0+fPNsTWF8KuH8Hi
JwYKEnj4wU2L040j+ssHqlEWM2Dr43HuiYjiBJsW+GoLmaakFlxvfmSPLSbGJJBG
OWK8vmr2CEOvfwB3v5OHvqB2Jh3Bn6X/bs3xHmzhU81Z4ICoWzHvCpy5AgNOuDvr
lGscCFB4AUsDWN0iG/3j6HXXasXwBPLcEpCXg+KKjFMAKJfQQ0Yr/5crgIOH0vlg
LarKB7aau0ArW7xTmxcWuLzr9M6UMAXrQcJOHhg/8CPbsnXBHDVQ3vM9fWvBDzf/
iGGgNPrqaWROMp0HspkXQ+PKaGD3Ban7xnZtDGlTdZaBGET83L44041QFzjkShCt
qmHvRoouEWI1PnSc5EkvFizA3kJF5CVVM41CNavosIEfpB7Q4TIkYR4MQdHWBHTD
IPGGH22V/wH7qe+XWTHThuAktFXMjTez6Dbcx1Ldbl0Nj3tABRYdq3Hl98k73c2N
7mBXyeh/LjMagM7fctW9GU4oVgeKeZ30QsLzDVN5Mo9Sv5hzBept4jqrRF24OdGY
s2QfyhAT69cD2QqtO8RNNKfcJVKlf3BD0gKEN8PR0jnOr8JxJkKLIQe3Pq7MKnG0
puZ0El0Y0udPFds2gXn7aXNy40fhujDIdmCivzeYhOk3xKMjCv2MMRHgfi+kzw77
ursWJmxXfFb8th/vF1ykza1s+voFeVMkUt74X1BRK9QP9NwVezcq36L4Jt0op3tU
1mYZyV1ZE2rcel6iXqi+E8luJ4/LcH3s19EL2//uqWM1GBGePEMV5HFGGSPZ8g/V
IQ2KJYQDMJ/h3d57wEmmi/CC2C+RFlmB7EeqR9qioIFuu0N5d0QgrF2+r9WXLGUU
f7IRu/54ZBC0StfsbCBf9c4y/W/eXM6ocPHUxX0W2uMYlTSgxPCVI8M7fssJW75Q
sjd2FwHRayOuYEQ/MJpPqLDL8jtCDBvPBF2fnLjC8VilKGbNVFZ6Hk2Zis9NB+Ym
t7YLyWPaDCtp3v+aUqUNhOiNSFMgDEko7L0SVtbn0MfoESrhtIxNEadmqgrC+mXW
rrVsw1cB43kTDsWuFORx6mFgiWxJ/BnFgfkdCQVvLHXKcVmMsUxXat0o/iFCEQVc
i3CMhZ+mET3tya8cbAoimVckksq2Mv6N5rMv/bmlm2PdCWPrVCjz9N240bUz58BY
v1HZrbE+nV6Lj/AR3U2+zLTcK/zcD6H9kKxudTq+X94C2fMjF49lXN6GdOwum5oG
rL5WEqVWyzcG6RVG73H397l5kbj1lnhntPERG37tSgh8w/QT6XRspX/bu3YzYyB5
cO6cpvcv1aJ7VMAj1K6nA1+vfLd4Jy8Jp5P1pjRxylS2b6j0OylKtvLTBtE0Lp4g
hfBsL+EaFSxe7jlVfZ2SIYNsPD7sTS+Ygunl4ngqP3p9LCOKyZcvkVkTpP11DBKk
YdMa3No/5jCLImfIlEig54X1fHd8ilZq31E0PUMZNKkyAG2ylTV+KS5jU/ViqUQu
0YjwFsgU0fe3EW0iUA8vbrue3NjEqdSA9YY976smxrzsMDgZawimuj2QX3bxHG+S
c33SgEQe1sAWyezzAm9UJIZ5ugTPXTNMb9TFmpuN/Zc9FrNOTkm7yhUGNKtovCn/
eOiPv6aly8FQeE+fLw/PWhSrbK7A+sdyYdrvcAegOWl3wT/B76u2Ug60WBZ3pfuf
AdGLAcZQaUcyNczjDSKkgc3B4hq7xGCwcYNPLM6svVbA0JeFqDIkq7Jj6lGNXy3p
LPW65tt/uBl3ay1DRTGq58g2V3rJg/5iLfS8Eba/BcdUD9N9o10nPXxGa3YxPKSH
lOHHuT0Vb88k0kfI4kW/GiulZvmWd663sBU5yBHxSVnJQ9s32oxXiZZe0vpF6AxA
JrjKU3GomOvtmwCUC7tTpIfHCIEO59rIqtzfGOvh/CDjOflEoPfnfqV66hCIrdKy
plrmqvMtqNDhs4qMvM/I6DA2Ujaj5Wl7wlIgRJQ71+CrsMLeUYfYOfObRJ/s1HNm
zPALCksEcxbpPAkj0DQTJMwOpurGp/MGlwC984ni4/MqEjIkK+JU5OD9y+xnfPVH
C8UaYyjMsFt5gjDqsk5vP9jzCDdfhfYNjWUzFQWfn3YY2J4dnt4bYXuiKPixiCSJ
DwnHrbHwWzm41keglahx2VQVOOuJY2fAwEe70xuEfWIfyIg5+CD0zJu9OwPwOnQ0
5jCT4zw123WlQ78qEUlXvkmZElFKVxAoZgwW2397mTjyZTLMStOf/6ztxlGterb/
klg5Nd3sQL+RciBPMP3Cg2Rxy5KUeGCZwtHta1mHD0s90A2dq76J+qXvnNEV+r1z
5TcjEa1zRxA4aXmHwShIsqLHKw1d2dx696C2R6T89zLvwmLnAls1YgpT26brA9Up
0MUMXAr75L8bzWP93dUoEuYRkh407HViRbnhOe3ZsnMS+Pjabx6Pr+21Y2DZp+v7
6cyGiEVgMQ+MzZFWQ9zqtQ0TTmtsMSl/70ChTAn7eSBnfSQ8dmSm5mojokVmWYo7
4aur4olEskc4BbQMTTyUJSq0CzSxUJ0uLBY4J/CsPPfxEIpEqErNLrfujFPhhgy/
eO/G0CyRQ5ezvk8iai3Ki4lDkPeA06uwx+hUwoXItg0ByrDI7athd8eFp56S/Ki8
/PktKRbD8WK0MDrs+AJiYm1s7f5nEtEfZRu6+tBjrXHEMwxsCA8yL1FyUtR/Fw8k
XwsGZ7omBLZqZl7p2Vz1Dvq2KJzeJ9CMk8zZNZI0d26grDwsGJ66U0q39egAeTMF
Wj+xBFzwK0oWy3OAfxUkJ3k5v2ZT/qT19MTmxHO89J1ecdu0g5KGYWcK85A45Trj
LkfobzdrkqGOC6sRN/qhE2i+Tpxjw8CYBfadnnFSI8QiF4ew89dWDJ2fHUsSmS4U
sUYbuCKroTbMo5UVOWu+blvocRNCz7luC2sqWISOn+NyxDfmg3IiiNyLvObq4jrs
Eex0C6d9MibOE/H31uGmsLWKf0ige5hdZyyXfH79WjbW1rakQE8KeL1iGOGiWJno
6vEODEeQfY3lykKJgAzkLyRs4iKgjxjX/WNK3jpTzDqhUNSsrFLwIKdRolONgKAz
Ql/eZqyAMNP7aGPOpgolAN31ZRADFdmkX8pQfw3cgTOhtTjoX6lwuhjwYwSZhU/u
uLq78ceEY14gNtfEuLUbEfJ4bGJ0/I+Z6J3Z8HjaR1E9gWSN0QodmZjasjuBNQ3B
tnLor8/J0DYI4fvhtIfOCCQWI+MBD6l+8VgtGpv6PE/a6j/lA3Gytvz4eZr+teTo
YTDL86ihadM4sLlGhY5ditxIQOgT2DEBZrlcnDboBRxMIUq5ybQM61aaSK7Tw2H6
QLiALOcfQuoKtFEzO8WGL/gI4jPEXiuKxM2lKiueFDspdloYrDbRZCHfqzUNKJpI
UpCgyQIPLHPyHa475NlIwtxEGFKedzs7pe4NQPWAFhiBooX9NGWGgl/o6kRs6q1t
qk4NQbfSQY7aob7eGEDy076DZ+SeGjxLjcqhFh0g95GBLkOqAAKUylenBNQUoXXD
sKqZlopsLYZCPI+fVYNpS4X/GZnMzHWhVH2gKYq3l/6qJSkbkdzyHTAtpAPexOLu
83suG7Oe/ALLpRAmzocv60XaVFD6Vn5nOY9YTtlwOXoEqkOipDVlva8owOA0hXpF
pup2MhUxaXZ8gU+ewg6YMMcwLGcY5rfnXjPVny1tB7Wq6INYBlKuh0LQrWOjZuaN
SE56v2m+TLdUM1LattJO2j5WAJ2IHwM66UDOXismeK+bAG2df37KBe8bn/2sARKW
X44/HyHrO85rFpUcmho4af/NVxfcj/1VQF/BKUfZsRPlDFQ4XgBJiiXIBjzjUawS
Exadv7T+cW3usdCn7lZUEuEZLrtZU8BB2tCyvbjz2+aBNjA6aze9Ba/OzQjSNLZ+
HkmCUS+oaDy82pGLc7eRE0ZVfkCuGwaegeYIuPPK+6xiWO6k4YjcoXONAGwmnErZ
HFwZ81d34f/r2X+4HbIJnKenQSe10xsyz+yTYJSqIALARvUHV2JhOxmfEBmEmvIp
pO/xLjIQ+RCHgqDMbk5n8sVeIwCAto/wze+YIYFZP2YoSDYfpmceAAFIcAKkJJz1
Er+9BvkHJHuiGUr54NocjhfihgQlnGpslk/CWIwGMvhAn14/qOcVZjQ0zPJtjhhl
lY0GiUST17sckUGK5Ph8QvGJeplS31DqKEVKHsfN1IM5Jr9OBMIBp1jSdX0dECUZ
ksmS/M1MGexp/8r0Q6r9VrxLMvQ1NoHqD70bP/Rb/zg+68NjzGnNgFE5yPhlsuTy
BPzHw/6MVCZuCdsAvMALkTizeExil8Zd0vQujSwhKQ48BrjFm+W3SzEwZcEuKcnU
Jk5gZWKcHlH++EhQRT8h697Xe495/8hJQM/nIW0/TtTa/6okMwHtipXTDciuILOg
hmc4Glq/ChuCUXVv/tnggS1Gyf30bGhuVaLXv05G4tNxkAh5ap1Ael+sg3lwIScG
0uh+5ljets5fM1hRdW1H3ModZn+5UTXHonk3+k+rmT8R8BiFEtrcCaADj27NWYsO
PR/9DeaCL+iwF7xKSPIOv26Wuv6xO81AY9GC9vgHXRpydXGM8NmUu2wDqcQfERFd
rUDgqr5ztfrraG6cU0hdzBtgW54GlEH/I/o+oFh0KA8z0HeGLXrjgRPUph0JMTi2
EqjSOFxRpA2KOIKv4Zz/2izAFgkqnurLK/6BJlbwIW92y9UoxviAw5RPAMs9f1+s
pIHJ7jipOWGxjyx6S5MxUP6S4q+PkZnVjffs/1ug9ftc4lx5KLINaXyisqvY35HG
gfwZheJJtJwPFrXPh9qX2jK5l7mQIXKNLLfCH+8QLY9b6vcOps4s4vaTkCJkFl8G
Am0j/YFrC/NJzB9BlB0KAlTHzozt0GcWwzo0OYtFpncAMwvty0YLRmdUMhX8OmcY
cEIbzqIfGDCgu//oGlKF/fOgQZ99GKyjES8t5GotGfxbUu8r7SxTQAoDEmLAfGnD
NiGFdh5hrbRBR30eJdZb1gwnLpBn8m12ISvAyWcSD9rrLJNEsEzaI6/LIOzyDstY
t0TyxFNxFII1LtgfO+Y+t7zivQfOTe1ltSfryjU9Y3vN/cXfncJ03HokX4RfdjlT
ycV6L9usWORJL778TIrNpKYTeXQ84A2RvdUfADMaX77Tu3nNAi+uQX3VUPiJtQyU
2r00uOiP3/uY8IGKkLOdJkPMlruoBENnHnO6ofAT/322CIY3b+45105uiPRLX7j/
nwHxZzUuAEzHoVpPIkrTE8wr40ryiy7dpvFg1I+BL6KJV0EJ28h2orf41DEJHXhj
8mLcfMZMD/WdBvS9RPu4LpzN7aOV+6QI9JVxjjCbpSkYopJaJLjbZ74+aRKZYe/1
oziLLVA6NyQfZ7VlVl8ckvtG+4ntQUho/p+4FbqYiiWbpoYu33YT8F7tX8hQBurr
+js4oIQvFvpXpO1CNeU4zr/zfy5WMrOhZ3zVYRDBjh/ultWKRfJV71RSmCvByGgR
vbOvVUDyEIHVbk/MIamE9DWOf5bTJcvbFSuusFZfRYhBBGUOlCeoNwig9zVDqf+m
mT1AtjpE2nR0CMbEjdxS9uc9pYVshX/Zp2eSx84LhfsxsRojsr5lm++yePC1pK0/
Hbqsnv3HRSgQWENkEJ+c7g2GWDrdcCzBpp8Z24HiAjFO/wezrctPruf0ol2kGWy+
ZxpxK0TFoD5yDfSmS8bKxTmn6TFqqRlxZ6JTneo8fJpjuu2EQqJ+SxoLxLEWDZW/
SZmyqXyZ6BqFUk8iRUNkO/0sCx3QwMOHyJrkdjghJEZ5kDIY/EjvbKGsxE/zbs3j
faYIvR6fHOil+9vzBRq558eIRK1PzeJF65IQ9g0P5X/c4xD3IkikLF2YZl3dfG4q
5eyfzyV+leNJFYSgWaL9MH8fMQPcsgimU+FSg8HiBX9lbaCkQIithK4FQ6hz79e+
yayoI6hFu64TZbSsajq8sPWjlc/4kvBkMed1jq2EaarlOF0nQ8ozcSoKVX9K7K/k
sSS0VLSTHh532nJTSPGasEVBOSytO2q6F4h2duRPadC/Vlihz8Q471Ph42BAN4BP
le1NRrRXgqWMWazZF8rVQS2orNmBKH+ZUE0YlsZqUk2y3kJvKdH20Ai/I31OkJkr
+U14jPbMdlM9HTPuF4+QANEIE9RfhDdPDbKgcAbgkNwud3H6btq1F4dhA7N+pK2+
4Vix8XbImBvANwyoDa8regNmyFA24NM9qiGUnMLJQgC+04nQdjxMAKAWUp6aOKmJ
qRz/HvCb6E6gjoeUh5RjQ9mVqs1TlhVXmLaOOSHkIhxLvqgAqRx9ihVuzlZeMVN4
ze2xMSc44Dw3lQ+lX+rrnoPF9dHwJ6phEBxDWbzzEJpJEwfU64hizIKNUBwy6kuT
LrDbC9x3A63pxPV8DZe3NM+Zq0Fzgxh4vmIt2nuoLGo9Ptl4cyZ5s3tLCDdP9O+I
o/Npwmy3Pk+bC9KXOtAPFolSzM51YWsXvWyK9vDnnn4f18zSgnLw2y7khONpms8a
2MN0TqAF3yHGJizEvsLLZ4rgYE/j9DAj5YTMjcW5rytJq+N5kWghR+tozCBfMRcp
+MSjthFEwdKAxM/dNFA4Uo2kSVsD0BiOd2JBz2FulGo/mGnUCDIAnL8ZwQ1LlwkD
+3GZ6EkTzx8YJ0L1/9hHEQOs4oSSiHHhb0sV+BCC2RaMsTdwMNlYGWFxMfyR9lAo
6tsl8OQll8xGaenHWTHUErsQ0XK26jYxukCDvPJozLnGTaLcd6OSrNagwa9l/fN+
f4SP1Tkb+bY/nci0sZqTX2ormTc97p8dsoXOE+gdqSOyLxnSkMR7Y1DXMtbPMCBP
XnLHwCZ+9F4Q6kpnb9ac2eSkRQD/3wC7cEYj5AizlFcof5A3uvipCFgBmocL6Gkf
Ig6xpRUubmlwWO1DRdENcLx2Rf7T6ZcT/Jk2twe1ZMfRBfUHhs1hhLzmk/NoxjFW
Cs/gYy0vFDQNqVshl3N+5IGXRn/q7/n71cpCCqLrEtKfVCda2VQMflFZvLZ28DE/
lQgsTR40i49/zwAMf5Uo4DYdYDKhOqrGdIXIbYBYFm25MItgBiucLlJ/U5l2SooC
Q+c2fvrmAuoezeOW2WBeEn7tW84Qfs5KMJNn1PCSR0p6ALnShszocmestl/RB7qx
h0mWCf+gxIhsR6vyKMPSAgMEjsXzA29NiIybwnwY06+ORAWSP1dWecR3kGg1/oet
Ij5Qba4rOiiMF8CPnCEl54Be7smuvCpfVhVMIoT2GUGR4mxWPfexzvdm8g97J+g7
bJuqE0NBRSMgrLp8x+LQxUH8fvRCA6Wquv1iQ2txJ9KCVpkA3kGi+I4Mzi9kKePK
MiSH9Y7H3Vxievc+T45CD+3RyV8sQpZ+6eyV155D05nE++RopyJil/tPBIhgiKRx
/hpwAWHGjyAvdTb9XSmHTGzwKoupAvUTQX/0TkQJKsRoSDoxzKi6LZ84ur6QUhN1
olsWHirpKL1b8ACaWQS8uspbuVqqK62m2R22hCxDsjUxPkG7bOOyLjMEFfUh48OU
zFrXFD2LUm/9jSaxvVMmhqQRuHfgqAvfl82OT7jBBHnZzJym/Wjmtqv1+kSGEmyc
MNHfYhvvflfHLjjedGHEAavE1IgCKrLgtOx+sdxnSwOQe2OcYau5Edp+TR5Z+bDk
9Wmuohb3wdnViCYt7wq06mtRLi58EaDM5XVEyBIbYxM/Ck8pc92FN+h1oWgDhsyf
xnEj9sVho6G/YBdEyuvX931oytEKYmSlI/MZym/T2VaQ7GU4W9Paypc3okEJBumR
5iifPcC9BSjUBg3sx1W66yWn1n6XuQIS0dTEwpZEI61+PhuFHtEbjSz8PvqgPSgw
CmkB3QOz5jH4/0toxtVSMe2Zm/Zh812i9kOR3iJUN11LuiSt1HBLMV6bV4Bpf1qU
ZglBg3ITg/pM7awWO08MZzlUsMnNcl8MN7TqlX3mdT0sHjwoVH/y/26nR7RzOBME
DPbKLyaeTGYw5wsrGWEkWMvZixOGDS0Ym8RjmsFihRTco5BzO1ypp4sakK1FYKXJ
jaTZ6JJf6ILkXoQb+kRH4SB8xexT+BAEjLdwTb88OhdyHjiZRSftC4kdIE9XhgpC
uFJu9UH9Rs/bDwT8xRr53lt1az8Ah6VbHBK4x5+8Jwrd9mERWOFmDC4ZqjZIyCf6
6PjK7fccAOzbkuD/vmLSPKGGcJ6gQ4LYW917ZIfXPImV2xrlcIRFvJqusRUdcHaY
/oUEx+bujAS93ek8crHwwlxqkrpcaMXevYdJnIWwmrJ6I3PR9ZXSebhfU1kfiKCZ
RVHnvV0vULXkc0ylHELnMlxA7nonr0GQdSsuHt4o34umwt/kZkYE3A/AIKZhx/Kq
zZlZ45wpRzhlpxKEJH6N0JboXEVMGJtLKVp1u91SfLkwqd0DuUu15B+IGJHvaZmX
SmmrWIVKFaFjhdxyTLTgX7ONGa9x8FJQLNrMRe18KBMvjNQFoV5OXDCj4FmcJ8Bt
IHttZ8R3xPTpWGX3lqF0DOYns1lVfPl80HEcXSAb2DrBm5ZQsY9wEjOZMb7EOwq4
HdJxlmbhJ62e+IwaLivLPGrgCORkMUekmEVRVNoh1aPLfAWSsjEd+N+xGJPqCBO8
Ydy/sfKZ0vLVhp3fNiurlBeeFy7CwwPbEAAdSWLEP/lBnp1lw/XGgTHY4KF+vX6R
eMER0jHybMrW3mgwYcCNTMjIrTp/gyZ3z3O+MP0paEcqukVRJt5pmbviRNKsFtiY
H4buXAnvPONGtxA0HKry1k9EUFY0fnzl/1r2I1oeiZ1CHnZN2+p4vE2qoIF+6GOa
mQsAaWiITyMyfL4xnRZrr+ytKV9o8OCW/EPrfqR7m0MPa01/vbl+jmgJ5ZGvVR8b
eYayZg9jGTgAD0wse1fF++E2tqc/6AGN5b7/NAz+7J9/wW2rbm6fwmApMhJCU5Ax
WKGH3HKtOCeNXdwlAKz1+TPVSJXmfGW+kiZKGhpE65WDXLCodgkr8um3e2EXsa3t
MLsGTefORkhJU0yMWmR4fQ6W4q7rgF/2YvFajvjWENtRtlur20A0TkUxSm/a9Ao2
x6AS9EFu+jtvf2310rWHE7fQLWE0dTLt51ULIYbNLOJ2l/S6YydH0RhFZ8gPyz0j
39wowViO962j41Z269H/kiDeggtbdhhc/J50WVvEG1h24l+GEzWiJAIkNJn/XWXx
a4aTU8GHMGCqviENdTtLM2q2FiOiHEfOO8zfWlBbuueb+5oqzrI+tOK+dXvpyXbW
79nNTYaiptQriUio7Xdk2zC84yY8EbrzSe3EQY3/gyBpw1CzBX2+9xbIbFhAu3p6
XIxsXAw49rmWN191XKElsFbJlHjguWdGRuzBhBZJqw6m1oPo3i68nzwkfxnuFKJ+
1ltuPX1YJXV5m4mJNa3zr2bXvnR12ktFH6XKaP5J7YMb+IzCHsAAEG8FrJCz4U+3
RbZdiVe/TEqFqrAuh66swhA9kwlCiuXUr7+2AOJbA7+RIio2vOxOCwlJKTXiv7IN
U5ZFgw5Rn9YZfewL5kOiEG0yIdVOQLc57IgENmmXrskh0T3uGfizCHN6MKEJMibP
pqi99VVVBCxSePfrUNhmXVa8BAEPyKGdmwupl+dDtXzkBywfj4s53WLgVACXLpIS
fUCHvi2N9Se2Vg75ZV6nUYoIAyM11VjuB9smnoPNs/1IaJyng2ed0I7LlfTCpzf8
gEyCCg3CPclWoSNKi/pHIdv9opEeSw4ajVLK2YOYU53O2LJ+P9BAm0G80Q6MQ8X8
e6s9zhq1lZzqu70zhdM9jPX5QsYYp9U53zWCgIl75CxTq5FzkuuDTNcgUGTmUzyB
K+gPHVDKTMRBvdk7aE+ESQQsZXQ8ffGCRU2NiIp0czbRj2GIa09seTSMAKFnKYwe
dcGgTM2BURnmVwUlmEmytm9e/KpNo19e7quBESCsQWR/CQFC0IwhlkQb1TNglluX
y6euToXDrwKPHCjjJNU0tfW4wD9AKV5b9UFWYwrkElcHWlgZL7rzCyj10mQhNovk
gObzRcFa5x3oO+mPvIbUXlofCqJAaVB604tYznO6XuluX5T9FN1KmUECcjUPRa7P
gOT/iXtL26jX/xLAu+sP53656/I+IVotzsnE8J8Dj0kS8UQcivOkSSaIXdshnczW
QI1IkIBOWSnl+nG8GK61CIXCwgvyru8Oz72bjxRBX1wEwfAUUo6S9223cUzAK4eH
YJfh/o78OQYSHGZRTmOIVyE8v8pKzMoxH9BNvVzBgaE+XChmU/Y8BlOVQeJXqIiu
+WhcnQX00XKpn8erPYJhiIs79sVPvAYvRW9LMjAzUrguJjDCQ37HYWoR0eWchuRF
J76p8j7jyfiOAoZDir8WfOpX8lDVC4OD7Q+uiL1Pt3GdWpo0u39Qd4KEj2LykJxL
t6Y5hXWp+jWqWM63nHqIovZqxrhULrX+xEhPPC3AD5ZJGJfKX9jrS568LYalbM3x
fc7ah/kxFaucuO7UH0FIO9cyLJ4E1S8f1CaRiOncpUh2ef59+FDxiE/dpFJEI+4a
A4ezF//ZmnZJyCvdP1YxxMXqMoaI01qe4zcBJPTKklKH1Y+Oex3TJ/p74PNxxpEn
lIFiAkJTwoif0zFIv/iio4bfqJvWXBH/r8gDNFVRNjdkGrTPsPG0iHHIPzeaX8u4
tiKne1XU31NjJvO9jfB1B+gi6wiFGtuDnLGl+DW6pK3kmsJxpMiQ+5oJIdk4u2Tj
yNoUFAxexyEp7SfB9Ya8TRGQGOyR790k0YS3CBHkI5RZUhnn3XiOTqGx06YXnqt7
05a0iozkq55RcLm+dot0klyPz61WK9LfGPw0lM4zuaJXortt4lcP4eX+uajssOsK
8qQQXdwGSiQmLE76DqyvAIs4f5xoO6QC2YXL6dS9hjuvBP3KqEI7lLicFALihW1O
Nwk+dxf5OaFBFReunDo/NN+vIVHUQiQe1VjkDwASMsIT9qUX9BRqhcwGWTpQkkv0
IOCbZbV3+1P5It5G4M6eWk+LjbxcRnPCmPR5iLMvFosvEQ12awccy123Cd3u+/Tw
vIdxBcNEoXZy6thYzyRnq8/sCafTfGGWNFPQb45TTrZoPFiff/wS03ze0V8Yy6ST
S8VISNN2Va+o1vje/ltmTPWlyFZKNm5g+4T2nSEJhoL/l3jQ1/yKbOSt/nIvdKuy
J6+FKu9vMZAtqel7PNl7N7Iq2Zmq6cO77o2YTDDyiL09RKmwgUG+goQf1dvcRC7b
mgT743U/un6qYd8Pvb92RmGM87nwfXSwbmoVWsYnMmj/ocwCKWDEU9t/wKzkWDoD
bLI/0U4RLu4B+No++wHmLg47CQZYFu3NS+EtlQIbZXuXgBwcHBBCt+vw4H/35Ebc
FO6q5sxN8WnVaxAYz1y5Rq4WOgC3Q5rWLDgu2e27gUfa2CGFMSwmc5w/pcIdBGEy
GVdsJRrKlZLk9efEhoCsM4fMPc94JZuZHrdMBSKvmPlPJlpqwO5Vr6CmjLEleePQ
EafYC215I2rVf9a3XLm/N/r42RVxKyjpvka/YH/ndkwRVM0Gi05prmqaKcoK1e1L
rTrGF1ChCoiGLG9vIyyTFyslck8+egcrjjyO0PK2D3wn9sP+NRKxj97UxiRwQ8GQ
+hECgRrihIObMuxoq4M0JGsF1HiOfiiU5lngFiSSSb2pJ9Krl4mpj9+nPL3cBGc4
rLhO/WuoqpfTDF+Vkdvug0YM2tEiaBaGX7Pd4IUTj5+k2RLi8dNthloJOtP49oil
kSJzVPn7YEJwBhdrYjRS4zeWF0ZA2iMgXpKJ/dIwNT0dMva2RH93q3yAN+UvS/Lt
Ls7jsiw4FXhzZ/ZeEVa5mjQM42ySCvYaupgSYKEo8/RnFebM+6QOq+zs7AmP7oKa
lOkX51R3p73PROmWutAkFsX+Y3zBCn9UP6LuHwUMVD7nFLCqhJfZ6T+U2d19oP3o
fuziX8M/LmlPLgmEQB5Kd5FRjMr0a2U2NyqCZ9omoN4x8QG6LROXlUbOCZgw5mU6
WRGiwRHifeYv9wz/p2J1lhNl9zL8tfQhI1LWVGtMegY1fLbwdJXQ9fixD4PWIwSd
cZXdnC3oy3iFaV1VVGieEDuAEZGKPodUZ6UvAJ1wNqP3tz4jJ0oJQnHK4HktQQPk
kxqMrPFhbFQXqS3Qxa0C+9i6nEEMGxx0M1bt1v5dDv5p1QCoHxF0JrYqGfUpnFoC
JeMHXmEXs9Of76K/KaqXrOgIn1Wli3LN/aMjLlj7uHGVdt9Buc520zSPVnlfrgV9
Zath/uROGIKKaEheoPvcaACQix5AkW6M4uBly1PavOsVoXuJAaOsG16/s0v9MoTY
Ir6+3nvVUEYCbFF8vUDo/dx7Lt2kIvWcCOcHdwHr5VuBJESBHhuykvY+LhmD1Jvj
6XfQSTjI5MmkkxHlZjBUoLbcPoHac0YC6xYwZrjGbMVMfuZmyBt060METa9BHazV
KyC1jPG5kB7NiGeQ9P+xoBT8guXyqm91Lau2DrSodv/yuOlg2v9MEaq+E4h6DRME
OZEEJwHYA/LG1WG0Q7fPyC+aRmNjMLfbSYtqQtLu4DgvFMIQUsDONCvRoDFtg1ud
IqBf0aDQKE+I+DW8nPq7qaA4IOE/cRFqd/+ub4qbJZRRhBAzb/pbN/FQCt/WRYUQ
HJfZHmGCCuTP7PokWBcRUsmERt07avbdm9qmv5B1MAqeanwAxm8mKACJ8gd+xEQ7
byiOU6DAa4/ZehMYmHuNkMEPqJczZTeJ+KTjob7Xya9rPXxzXjsf/ZrgNoHUURc2
n9QU9kGEb0s0rIwfEtv4C1h4DDTNSBGClTfffSuabcJwQu/MPtDFCcCAvjyGFoGb
761JQhVrCYXa/V5aSSTRtaKgjYbQBs0OaWBrT9R5vTIDLrSgPeMpRF/UlPW5xX0E
DNjotT7SGEIzXGxEsyZN/X7Fhr+jS8yn4nrJOomszmoVkYZ53eDr6UM9QneBX7y5
IyApyufckidjrJhFtm1JCl9GKdZh6IAHt6nxvjPX96VKUSgtgtNqYo8JdCJL3IvW
R9bgTYxVXKH03D69DqdB9avQDidOvfQgPu1+c2kZfDC5BIV1+ArO6FooxYh5tLBx
6OF1KayizsDiZ+sWbhgLp1TE+DaLAlB+1QRBvXicjUTUEoLRDgX2y8BRj+iTQOXU
ncTkNKkzbZW2wo4F8ER+rd597lLwK1/lxRIN7llH1AwykXhGoRuQaLEd2A/V4OpE
XlUhz7Gyy5bqyoGvSCfaqrEK6IRiDAwxCL/HcSStGx0JYU6ngfWJvgIMoCdBaFAQ
IWpf8LoFiNjEFnOeCghRJy+cHix42PoQH/s5w6hkBDmVB6yEC2Yw9cqfKeRaT21d
Yeh6g7mvZsgJvbvydFdpmqRUYmwWeH3V+3ordmxR9qfoQnD+lBw6spQ0zGfluQX9
bgn3vB3UdgSo+O6OHJOXu4i6q8xUQJmdI4btNeMMgukG+5q7T7dBCpzKU32F7rBg
/g617GB72pXmjzTMV1ciO4nsDs3PmyUV4OScV7Cv7AtKIYlA3OTc1+GywdGbmPsh
BPfrt7UlA4Xjl24UTsi14Br7uo2IhoJoltbZ5pxnQ9vmVB8eVz3r5kEwAVATgrM2
JfMlE+qw9pegtURBJFMPteHBClFn43FnIltN80agnIWLVVGTR9DqLfxNZwRhizNQ
BTagYhMKXqQPUwnWeP79g3oLscfa9xLvbEpW6R9kZ39a9Rk7v58gONPnTWeTdr2a
UsQX92Ci6BdTUMg9WVgTvkILhrsItYoMU1bXBi+kJ3b6K3rQrzlVeM6RD5YR/n2n
AZgSZEkutyYpyLu7ZfXGhnPQ35mCv6ehYXGBzZgE+J184LMzqHpG5O6cg8qCsaYd
G+GO3Ae0lM3zU9O/NsYIPG0K6zvMCNCYbLCsWJPkgewxyeaTZNQD9m9aVFNYBb7V
He2E2SIiodJM9uZHDzgg2ZSoX2oh/yH/NeWU6qS9KeZ/ySCDj8p4Tdo1TV7yYubf
ffJUNvtlIOp5PDKidp+QEnv8SvxjOXmOvq22SKSSDDbRzUNengKOk4kPZyY7kW+O
SZPx0xu87SL8m5S3t2Okk9uZdgcijzftMQXJoGJinefHEeoOY0XvoJZuiuRQgDvo
bARSYDt8L3EU+QcpZ4ZvfJ6JPo70ODAp0M70Clzqo/3CDZYoiqdVrPUB1Nz1cfQO
1Gn1/8C7FnORx3nbiFGiBGVdkx7ww8wH2Ih8onbcbaxzNcwvLL3RQeVnSLoJrHus
Xdv7YDCAulBoOh/OmYhm6rPpD3wYCgylAN9yGY2ncADR4dxCgAe/6ceA6nQpv6Ym
AxrYUNYDdHrzIl4zbdAWnRZloTAe0jGKzCGxWM8NjSoV4+6stuA+AxUTwF0S8EV9
giX39w8kyFNicU3IJQQLCKcZKYh3WnIbdEuIgXFEBkUEwA6m2BWF+TCUAOV9e4xh
g3cQL62ExzCzqUKdwO6ZjSscXPJ53XHs/H8BJf1Fck+w7k5Kwpwylyusz+s5kIXp
5OYesVhjS4sHNsnYxuSksDA+Q2WJd4YiKJOkgyPcMzybInZESbAL/1LXSGq/NUcB
xxBhv9QgZPbHgMDyohE6KgIhnnBMi5w77z7D7LCAHxSW8JO6gUtBy4NTWzv+XD16
RSyNUrD1VsFehg2DoGOOYQ8Q0gAjTQ3HjJL3sNNrM/EjJPWpd1NJgCbcXgOLWcNF
00hR4rnvsU1kw1Aam83wArUAtzuX5xrFyh1M0LVPwbrf6oiiHQHGvn8EXfqhRiPU
hhF2wULdGkHDjUFkti+9tg3MRpUW+oam+WAe9GbeIBQlP9/2Tp/greDlZdNlucb4
w2XGn6ruPTV02adlCQJHGnutLJbTeU4Z/RdGRj1aj8seY7aWeZ8LvJNTOzf1YGSB
ocvxaTG3RrwBR7sEOj9VrJ6c+ObuU5YDYsar85TIq5d7px8UkZQa8GS1PS5baRrx
EN1rqnHzaJZeOGqyJ1YsgHhdmJ9XSjlh5m2fTumelKzj4cKglA17/j+xLCpVZDH7
GtV26yHQlMI+Kyt/X125BaJpUy4Y50ivNnd1lgx8WrBCOLFNAM9C92nsn5IXOPJ4
JgTEHrBYjeR5GoT1orsnzCchvkB0H2LQbIq/67tqNwZveyrxAkE8MC/uKKF5cOO1
rlBbedrI5FyyjWof8gwHcgOhFFw8D5I3wM2/X1f7vNiEFxxaXWIO9wLt9AwrJyl2
ge2OXG+jXQSH8k4hEp0o9s3H3yy+QWBvrePYUpdl+j6QYE2jDU6DSaC3PAUSL2BU
CdngPP/RmV5phMhu5WlIqzo8Cllb5JA7fuHp4BpJFgoun5OWhuvhn3zw128n05mt
jhBAyLbbazoxnPEEcY319Rv5zfYkvhTS8Sjpb9IcA/+FlYqbDP+T74zw8JcebYFo
fTC4TucTFCRmnKhEPHwXjMgv3Pi0iBpAmIDsHhDTyTDY4R7adViFhAtwooG6BU5Z
NBS/ujZam0x4AazZhGwxrPyBwwUvUMtVwhKcJ1gfKGVS2bg3Lv34UvcxtsWfdlC3
+OTBpvkJuOAP9GB8e46QRg+PIkoNIbNhV/vDfLfkgzmh+w1iQDQCCuI2tlO0Hwoy
cWNABwMdqwPGbTSN0dU1kWCifH6sskuTqB3Y0m6IlMQzqz9Omuyc4qraTK6r5TbY
e4yOQRW/w0hcZnnPLrS3a6+TNLTewTHRgnaru8yzR9WRU+faRtyGDg0on3nAcjwR
wW8R8hjSfRytpoMsXgTbd375gTbYfqugTA2hpkYtFlaVNpvts5rCbT9gWpXTa4uM
5xApcxXSdmyW1fZV//jFYBjS0p4p0swXj+pr96uBjJ/iB5orrEd8u4KxvnurSRzP
i47Ldd751tZ3ph6TqBiYGvsvf8DqxhCVGrEXwlxqSj1Es6dLBlROJ8Bg6f62sYi4
JfxzSJLt64DV3ZQVuZ500j6lPaNJFZsQA8qrgCKcFzek6GWdSrupn0hb1rMj9PXb
tKMK7HIGkacdI9FbP45wKIhc7HgsOV2jtgUlWdBq92RawycKceMJjDF4SKcY0ZQo
qjk8bHSdyhKmNZHjWWC9oG2Zv/EyT5fI7li1YL8AK9wrq/bPnVB9eQlnTI2TJCtw
suvyQIFCgwK5HLuV9wepGErTUdZqBynWNTMC0l7d0OKN0i854jH9U8CuMKTcwRbb
irZC0Z++lXKCmp7Yi6doTAaA4CUH76WOWOeepfsPQWt+gVTkPny2d27I3HmPUXb3
Fd8m2bjqr0aUlTn005M/vmTI0vlX1KPeC/J1iS8ehOzgO5eShCR24rtlTHm6EN+L
6INv3egxZ/LvuwOnI+f+o6BcenrvoHwzfNK2JXiBWUbivm1s8/td/GvS3XIJWTB/
ZBV9vmJnu27n1bTNC8rcpuc6++G8dDejTS2ZclnKzoiTbMd6+XN22J5MsCJZxTVB
Bs2Dv7V7vHHOfcJG/3y6SeGOaORTIq5Q/uRogQ0h5YT7FSVyPeDHyaNbQUMR9IMo
XmKyIk4ENMOqwkrQUoGnMW2VB6ND8+qx28l3Swy+S9MXPp4Ju8ZJ5Mgn7rwhJMGV
PeWsiyqjLPxydWg25cPrkrLz4tRECbqYI+xhsTamLRoEWD+ioAAfqOMbvQB3u2OY
AUEwuRHrzHoLO78VIGBFHUUhYXBIkQNpZG+WuRKoSkcG8pbufY3k7bT6ngV6jVYJ
VUxnck9kQ96OkKBTFUpJmtykoUhipyV0VNUwxarfPwTg2wsyhUQ3Ot5+PGST+jqG
drsbFJi7OoWq+XJS0f44CsdIn6NnOFwH5tT1Ey7Tyb5+CvXEbV8bCZCUcip6ek9M
MT/RADXPdJ61y5sF/aHF9qPB1EnHUjahNjsDSns3HCY1utuoa9IppeFrpPJAYEVz
zeVftjeYMdjn+FjdxUrJPiPAkSZISlYNSM/9gtKt4319+RgYJroEvmxEsBUep2J0
LE9j0X7UXQn1oII2d5JnUCvxywxRrr66CgP7OGS8xjnmlMMpCPnfRv4KqbiBB/OK
n104vh6hyzAczuhlJLHBXDecqU4i7chcL8BcgdVzXMPymHSLs7BVhwZeMdyk9psN
IHfoIOza8+Eu32j+lvYZsZiH2vPx1yl+de+ipWzAbYYMOXfuion34/ChK54Q9JJF
J9HD6xsjzs+h0yaCec5ohb8XOj7atGv9xmcD72zXs89/bg1hqPs5LSB47lYBSbAu
QpG1FmfFaIy77dWHLSEqYlEknUa13BmwxWsMDEhj1mEBG1O9ge1RwlpRBd7FhWzq
TNYhbHM2JbdjlfLjlhRm1rARbPnz/YThv83AKkvGi2Gy2fcqkvsQZb10U3Tp/1n/
zN0K/ndFBc5IOLhvXzqnOujCg455oxLVPjxuLf7yEs6jOeGFqocZ+Yw1oVsmJ/eS
jyFfnxT5mlgEQud0xfJCUX8Pt20eoWOyZPcTFNzQ4zbWfGhMmFX/DFhezFfTeBXb
f58XzoPYBIyQMQhnEAcgvkF8RWdehzFl4NdCPCMbsxprD26vYMHWGG7xj5PQdKNs
mnJ2O615ZaoJb8diAHCj77sNjTG2HoqOf6WcxBupVrlUEgV+/P7ETDv8OlEk8a2t
4qdOXaXcN8bV2jRVOabB1XzC2ZqKBy0VYPu3TJNLUqozvPRew+2QMt9BslNIkHIX
+mbYUx+TuhjECOdwMYyEvAj2SLKZvOLKysNY/XNUF83A1CxOllJzHEZhKul3s/Fm
xw2YYE6+BTzvm91PqNB5n5giD6/UEkkaekFgEcW36bsGlFSwFschkIEEb3aNmgNW
j6xpTF7rFgUddHJxCBjHqKWsigb3zAYxxW3XytthMVDi52PzjtUIoo0eRJnHJf76
rH5ot9lriXskAr0Ct+dt7jKIqyHHXjf2RCYTxJK74MRwjM3KhDgmJ7KkmNJzKqXj
pRaS9AmZpBngNC7RnF9FYl4YFFyr7y7jzGqF7sOkJsHnCWdrBfpnNUyH/DPzsDZ9
LidSa9ov1KBQqbOuX/HIk8waTBhbVy4pWQpMu+znhW/nlO1nZK4bQjqvq8nCWa6O
epNk9VC1Pe/799jOkBc4k3NTAtzvjLTwuk79sCrXVkEyOtlXv8cIDa+SP0wFTHcR
bintcakz9y8/KH5JMwT/MiOweFVgI8a4x/THHRYu8+PVfWIaYvq6RLfk1VnQWrzv
HC3q6yjgkN0Lis5RLxd82MuyaWk5dYwALjisB6kFrHoYfOVCukune5r+lYBo0CVL
GWnOFUmJcmhh8Fu3Nr8ht4p3lkT0GLNLI5uB5dw0rLqwoJC1ZOpqo9/dK6L7dp3u
lun+KiW7nT1B4voJ0Ur/JUAVLsHVjQXBuEUs/NgpYr2Og1bpm0CFcJjb4S4emjOl
IRjh4tLierQtzA9QAKb6sp9imREGYjSPz0oITpEA1CgdMS/yVG1K/HffeIAlOfWK
/RMqEk6UI5IABKvNckcBiftM8halFaL9vx9RhdCaV6b6qVaSYQpGVvNTf4QgSfSE
YDS49Cq3ZG9JZs1ysdQ7uwLRoHA+fEVqsZtgjSr6Z5jc9TeapnFw2bpeTasV+aOA
rUnM0RN/hkqynq4YQXQlNcZ6I3VzBT5Q0uLJDcWZ/ycc0E6dwAtKIS8I9R/BkUbU
OFZTJvjEaBSlJdhT9DKeLM1OO9fpNVFF72mO4+8hTtwraqYRLQjr2eaV5Y1eN70S
5HQKGOtZNAPDanmcAJ/uq6kYozHJgofHuWClYID/d/9eYJRCy5WSoz28osf4VSr5
qegzljmxg0iaHmCeqEfLV1NykB1jlVCE4MZEUboWg+2KzQ+OFghvs9XUee9cYZHP
DqYXej/LMQ00UqWjJ4BXX7qMsRUgMGYuDmRKn+idH2QcMy8Jmy9UdYQ3uy5i1CFN
fcaBYQs4qLaHBUQtATHIDVpzZlXew8PV1RvHIOvzLbbrY5iYymsvmkxIrcd1Gqq8
hbg3YZ+/3WeRFhAzS5coSxCl23CPi//nxiMp2jZzvkHX1lqNbY098T47KlT75J0P
RvzZQphojoXMPY2OKUk0gsJl7kpTGfM6grgTDegYIDt2usUuh0J+WXW+1zw0kDkg
rKaN47SyqvNCiTk1dvu1dEdzJkEfnSI6lC+m2OXdO4mxMW3kYW+68M3srxNa+34z
Kicras/8EKTuQoqJfeXhZpospocco4bBWE/k19A9hzQjv+4zDV/1rqvkcryLfBxd
0ZbO95jtaKrpFxZkIMq4cLrRBlFDPpXPBeKjF+5ZXbYgK4B4bDF5OXRa1PMwD0h2
pSJytvPWIUhxDzmxVVlxiLd92i8C+LdCfAclpZfHbPRBQJkqqOWNSWHkBMYb4EmB
1ZQb3ERuRxIBziud9H03qE6n/5QKMBoBpbGkf4gwBa+CO/6oVgVzi2h8We/q03Po
1CWHDZ1olxUCARsaK+a3e4LsBxAD6pP8DgoZrmJIqcWW4X0GEAgIuTAuD1+kj2gk
FwYj5Q55bTqBaaKf02BLqmAAHNZHPDIdlU35tpMzR/Hud+yQ0C7a/7YF3BESIQ3j
vmK6gey7g3Ic6jQy+CMoy+hg/VYzh85kfwLhAZmo8r9vAN4VA/rXCqVVCRGebHOO
JkiFAwYLqvNQz9P6UJOXhos/frENe+wjuvs6YptclLqOHg++IT+48l2MTx0LjV0i
tEK/rEdAzWkVslsZOKBGGT/fVRhD5bU9+maj83VL2LKNS4W8JHog1Hgeh1TceDEw
NQZUQTRMypOqwkKZsQRyGjYrllLormT1YapyCI5rsI+TvvApPb6w4N0V0eHzGCVc
jkwkqwo3mnebhZpXBoRvk78oYNMxQLKn+lKaOkBZ+H5C47TMKIeVlcz/TSPo56cl
BRATKjisSUZs3hh1g64bAkg+8h5jlem1DbNZJItts0bz2SKfRGT5/ip37UlQHo3w
LBvmNkdX2WYQ650u9gCXSHXs+NobvGvCcUH8GoKS8HkOZxyL1Q2xRGQM5XV+4s5y
4860hD9touZiE3ghxcHs2JdXEnKbfYO6HeqI1IxYDNz5BiH5z+JXJCosGx1ufFCs
QBzBIkl6nG6YJrK08UK85uYZCu3ele166Ho3rUfT7wCECIPdU6ZCUO+X0NEU4qP8
auVZX5g5+OdpEBzV2ezOxla+2/Koa1WSt6rx1K9q6+7njti6z4g8YHkCkTi1Wz2d
i23tuEa0aVTg9hYE68NCKWTLDd3P1EkgadaUSZvr6ZyyOqbqZitRZUT45jdcY4ga
xHXCHttkcIIc+sujYflruv4FxKuzucJuB2a6oetmW9aDicEA9bPJBkoGSG20GYe5
V6njKHUaq89mwFcJctAHq1mWtMs0fhGugbenzNWqOF/IFTtuTvFM+sw7RKoHNw2V
RUOejOHiaU1Gft61Nb50tdnlcuimORVAcmh1NeM4+pa7Ns+IktSLyQlXqTKmB+N/
XGScRWCeALwCqnLSrjpszilNy0HDf3mI9kqB/IcPdxk7BM6k629qhwNHuSEPLCXg
fg6wjTxAhcG54s4h9nak5YMmDmxTZ57kvSV1kjp1W8OBN9skKJBeV+vtzdCfYzab
sTbmvrdY81PB9gKYrFb3Uc8t5g7kGXnHnQbsrRGugfjbW7hUbbu0PdhXtmkYJlIR
4JYnxSByXTamzJc+6J0gfgYHOb0rL/yy5QzYTWNS3dAVr7FigOmI7jyX4CUbVOCB
ImkpbTRlRnh5xFFUlGFpRegyW1sP4FcodVMzsGywRPqRfbrU9Qo/D0B4daYbYxkS
OqLraH7BAV+n6Xeia7FknnCSB6Y1V9uekJ9+w5Pgk8Y4S1XfVBgWG0Q3Dbpi47CB
I6rQ4ZeJhzKRlxAZHNnmHgYyh6OModQTln61kaB8FN6rduXCmaWnOqvF9xP5F6mw
y4B5aRGSCYuHl/rES6IxpFlwnuH7UIF6BakAqwfFbK/CmNtJ6xV/Xj/pflerTEmr
Hb43WNTQnbWqpI3lqgEJVBcyVaJ3O/bHSFvOlRg/2I0uz1pkq4J3BIv9Fhlsvtws
UJYRQAVkMGzLTafwMOuwmU7DQ1OCJmKQaVMyAIMvuWshKhF1a37/JQVcKop8Zr4M
o8DoAt70zt+Az+CTpwhUUDgzCx3sjgx0KkhgTEiriXcuCUM8ExYVlOkap2FyEB7B
uyKyiq+R5Aq1YoqTGo1U86uBjekuQnOu1CalF/7frU6l+Sva6RuWWu18tknj++ay
H1OB/ufokUL5Qe2i9jqyId0KydglYdSEUo/6o9BqqE+eVAAgPX19n0vzlHWDj7bp
1bt1AatOW55LqI6XOO7r4hTMFIlB0QOs+YNnvLjf1KjBSsn1+8Xtw9ui+UFrn3MD
6DqgSsH+rRIwqDTOLWfMMQDAr9vWRdtP7Kzhnes5Dd2tNLWKl1F2iykpN10H63oY
hurKA9W5VsX3CJgm7EvznqVNe3J1sTvf5gcAuqFBlMkOnPbI2rrLU4OCZqr9U9ig
0fUhCsgwqECv0YiXIrSTju72ILYgD9/yNqopAP5gpaPD6qCZc9v0bAmvlEfXAlSW
+4c1ALVuNWTWLrgFY2rgTtoMmq+OIScVSbMw0+6k97Gv9oCfZxCO1QODuLqr2s/u
clQNUf9ryKQI/lmlsdhZd0/VmvURx9jXAHuZXHyhYEbT7QEJADIkPsiDJqhEER5S
uznuEXiXpTzIDVMkXQM8whLe34JkiSi8VeTSOIE9lacnuyL9rgzOGoWEYfwOM578
HD4xXJPJfeeaGwVUF5pnGZOTB7czWSYwQcFIFY+B0IYn6Z/XUTgABDGF1m/efu8a
B3LlrQJ5IHxMC5ta3a5gdsYparRnLwJ1OoM3ceCixvHhM1dEQhWWxlcOkcPhBc9H
DRrQLzfq+G97NFEMUHbLNnlDufL/L+oNUZ6zxM/7sKD9qurA0proDl8PtQhVyWYz
k3zI0n95Jee5h4DERYufnFnmWRctXQm8lJYmwDyZv9SGwm/3PeAV0m2RQzObuauK
n4uURuJaOvOPxEzD8kOK5VDR9mZzSmoCtKKhmePZVd4jJu8qisWtcgK+GNlH8bAI
FsRyBWMF53yvqxt16nxhac4zLEGWyCWAVEYenXkOzWfBznPc1dBFl2PXSPUok8G6
LGonWZc2BsSkax1UGCk72UPPRy+8t8uPvutm0i3z5i8sqD/2VwX8h6O7TKVQrx9r
hPE2QTgCRzengYvGuyaHKCVcTo3XRw6jEtwS2aYNKMyP+Uwopv3qTUb1nvf/+/HH
vAS1bIBVPMIhDlZNaudVMkK6xmxnM7si8738w2JuOy7PlD7RzTnXAWXCgyrPrphX
k+idc7LSDrDTdGm7Y/e9k1xZGzgvEGdxWboOb+WzWbu9TQxuPnRGTNbMq4AIji8q
qF4M6af+BuFOk9mJKQ6E8jGCUi61UhTMrRD3mq0fn0uR4SM9ilNnpG51OWbaXmt3
RUxGSOLF5PIAhZS4j8/IYBzqf6TCUww9cnMguk6B7rG2qasRBfZjrcG4IsfcS/fB
AYhTrv03K1bHONFp7OCu3aewAfuoakOSA66Ehf0lk5W8K8pNYUGUVJUQ3olxrgct
9nIoT56HAjQR37j9cj7pGTEwN5wQa4N+pwD/XDFzDW3IPviDgW7rTSDyep84XJ8R
pby/wjjQWj/ewcb02uiR6Q3/lzp6IpU0lNovSaa6sOFv2INrI1kYKKPiOh23COvK
VKQvzcaNQnT25UmbmQKCcQfJZ90UcOKID5bGamXooNS4it4ZASjccZHzwfu9Bka9
oGjMol2AcaD1S2knk2+RlcFfsTKUGHHOkpYQUAuN6lLcKsWBa6a9ZLkyJE+lU9PU
jE/+kNlSus1N8hZtpVA8WHsqmEq+VtoxXAF6TViqjjY1s0xd/fa+D74TjLdPxxEK
Tslr0LUn4YCWg9TdlI6iqRnBcS6f5XH6annArpc1lv+Dpsg0K0mVcNvWJ8z/BAuu
YF+8AILTP0m7v1YiyvmyFDwpW3q7UBym82qgoSd1Gx7YiL+ga29oUmerUcVXA96Y
FUa9cVXBD7abXgxK6ZhZr0KJDv6JZ96ZFoUgViX2U4XHNJmMfmJNJTU2lb0JuPOZ
v/1lJmfLNAxDzbewTWrgUKbufh/P8f1UF8ApZsHquAgxXMBPfN1gBFJWZ2VIsrQy
jfofhk0ESgXX4okIImsriiR2Sa193zVGxQWAu8h6+25XYX1xKYCtzzSAm6QuVBh3
aQFOIgOq6c/7XC52heCrb2sod7g3UEJlwh9GBwjYdy2qYG/hPyEF9nYBcLeedV5A
ph6U9iyabGiSCQYKY6LkZdU4XFw4ueOKXZMQwk02Zc8hhj/jxGw/CSnZgNuyZYYH
gBsHODy3fTRBRMmg4V+v7B1/RDyyqIbdOLHUQwaZJPJpaKJrPaFL0jSoZVItNwGO
R7R2mo33l4SMUYQrDF3mPVjT1ZQgtRQdfdwRQAHF5jHjfjhIJn82D2ATPnxW9BjB
K8itXWyEL8hbLeD/ZplUA2bUNjgpARnO6iYMjyCNGSWNFpXXstwXlbQmccYZxqCR
V1CuJ9XBKbzPU9NBM/UiSkVvPZ3g58Ip1+TlkvK9WFzUoLaAz4Cdsw+miUVIPdPR
K5PjCElLVuK1l6KURgKi353AWew1V0CibDMLsTONmIvOcwxgXWLZ+Ema5yCPIaUA
1zRTArMyi+/Ku0a1fZzgf77+DsMJLtzxmipTpdcuCtBdyDI2xdk29YESyjnfZj8N
JIQig78V5P2b+CNKvQlUkQvZBgTP8KeGeEmB7NNw1YnalXyEq5FJuxmc+w6isWSk
5qdpTUwqiMcug2tcyxQBCPHo3P8yvUWZ37anc5uJ2RN4JbENm5xtCVznCwJBTjTe
2yBVhFnPIp+YefFWMTcj0r76m2xnsW7ykjngjO8q1XD295yhsDgAq7vYU601l3iS
oKIqpvfdk6OYZYVF366xBKmdP2JhVLuOo1oSeGcnevIglSyqKEQyKNdSsnckSaZE
+X2h4vSIw1+z3KE3o2NZb5DP6dORORJSrZmo/2hocqMx+0KNMUvCOYA6nCeAzVcA
EB+WxkfjknWsss7gVAasEN/74HtwB4vONShq+bDk8+sqXSAjoyaqYAFvwqm/Kb8h
buAhW1l1jYwsyT1h/W74AwrdcnhJC5YPmeW2mdlqH1aBoGrPyfHhJ5GSaCBSrXbd
rY7lE+Mm3++3KFuVr4W9LzxP75iL8O2a7kysh1/GhshwN1mIbxMdOlWG1MjXBQsp
h/6iyKqOKeiK4WH2la3QPtAB6sihwqRuPgSMfRQ5OP76wTLP6+sg8wwIfqBcuJZn
r4f55CDdNRdU9K04N+iFcKYYdKIMI5V5skb/RUov1DrJjF9UsvSKs7tZFKAaj7wA
onex3hkXJcqBr0NU8w01/aBKCKSMTVzcAdj8vfENWMpX8Jbel4BoVMym4vtrfV+s
VN0c/2ko1+FSo2fgDx7bDIiiAVIHFRmmsE4x79P3zpxo+ph8w7LpD+Rk4hBPYlID
XdUON5E2Z68QQHBLRR0pbapdrA9ytJ4dqKqGNh0esMufgztRAJ80Sji643bpdYzy
0fjGT9cqk0PeTsCl7w9h8aRTCvdS1ScsZsH9crG6GiV5Tq4My3bUWFCBP7eT/5Rr
2M6nutdA65FfQK7GOr7UIrAxMK1om/3FcAkK+IOINKCeoEBBfgQ9EUwSBxRWxGj7
w3AtPHp5Z8xQEncXdFbLc9tkq0hAkmoZF/lInYhqX28P1YPOT36K9W3wBCgU8MHX
lvMraoaKiA0AhhBKAzLGpXXkkXaC2JWSuq7OSFQmRRhudOnRfdTR/U+cC4YpvfV/
CJuuLM4Xp5rlTtj43Cf9+0w0Es+WGiijCcVmYj292VuWvfIk0zAtso1d63eFDIfK
Zrq06Cp3ACQs4ZXdvOmaeQqbvlx8IzNHfI7Ww1gw61Vp+Jzl+rNz0w7CTsBiCFi4
YIN3HNK7+mZmJKofm4PEA1zGDUlem3gGK2xVuNfZEyT09goF546qtyP8+Z8RDBJk
NHXx1xGrhBx/WNGBhHzuovKck1/v1qgczl47GUSQnobjMDEd+9R1a6cAwZn9kODG
dBQ+ZddaRIOIvQ44n+z1wQRrEebYBkp+kQMXtmPhwDegBfipr1bNCdyAeSPjfOsf
gg23P08MTdr2E0OI/AJtH9s0Zjo7cUMKM2+vNuQ70BPwszsHp6ULa2lXkGMiv5bE
7Q0eYSpWS95a4WSU7ZDiBhxzbfB//qzX4Yj7kTMZvsEsQtLM3YB+aeQqjyAU/gCE
d/hhUKBiug0sM4D+kHaYd5juhaKxr42vfO8l7YCEF+l2ncUHk2FoPVYuoiv5zt5R
0OJNOjWpJtm4i2OJzduYg1VCa82BuE+4iQbhzcuCGs+Ptmu3Cax1lzF4o1yfa1Ip
ciLZ1HanfwzeJa8mFPDQTtKaPNNI3f7fg0XU8x+JDmylh4Qv1YtX84TMFs47kZ1G
EOdK/0HSVS5i2577oVWtlqXUP+hj5HGK5p/XvzKfkQuJN4ytvXNIqLRdRnTXh7wG
GPrk69Ah5qmwuILA9iFHcb/0QPvKkhTagjB9mWAnEbeS5qtb5P7ZsTSNbTX275U0
2sOiYOxgr/JRTUK/xAUYFqy7Coqs6TLf3Z+nKbmSw/aqxpfy1QBmfhz0xaWw2Bx6
/TxXitn7WhcEHFeCxDc/4b1GL4FEbhhH/4act//IfSKrcTRwTqyPKx5uDy02Yq6L
nJtBHH7BXZcFhFJsXD4HnVEYh+rK78Nzj/CrIwB5JVLRm6nA+AaivorHO9If0L9q
jw9aXiCseRnRrMMWlVpJ06T2kalI2VTsEEe1MvyZma+8nr9BDwVFb/yHp/F39Wsh
Vys0mOobsvluZWVQ7JtBqZJw0/vfGK3EBeW/1YvcWihe0jL8JT7ilW1kCm3i2PLb
XeCENgssnZPMKfBcDnbAKo/h1lp+AjxIgctdh+hLYTiDNI17LK+7Gk3xS7FT0tLG
g4c3kfoUkjfXvPR8oqaCwnhqfE23wg0Rs/281JCUO35wLkHCwSa4zTDfq/ZYjlpR
0tOTBK+McgHFDtI9qwaPeK0sNOigm4SQ8TRkFltjYR7mPydhl4oQGXYgJPwvbrhv
CFJDYQ8alnv8i8hgABjukQPpXS1rkNn4/WouRe2We/Hmee6IY0tgTUjdBfPYJ0ij
zDGO1hPUBQvHRaMmELRm/t/V+J7kZywMbyF+KIcuqgTeVlSSp0ugX2UVxwutek4b
0jsfSOoHFfASvixDNTafRXXMcPeMDdimLU5k86XEEm6N4kXwslXxhIMlFbsrGciv
tp3Sh5ziSzyYqRZvtUSi1RFCXC0bj/t3j4KzyDL9FR/KCYRtklujYw5O0sXQAlPB
2Y4OiBpZ3Efi05ZJoDqVo0gOfOykBrtlGKto3srI2blG+ZQ2PxLTrNkULYMR1qrz
fdoyrjS31KPa9GYagfF7Fq3+jY4bqB8Et3+uRKpZh/mbZUewqSMkHzYbmWwonj76
qlw/BniqSnlCU2pdD0Fkmcv5UZsKD+T6zktxOjur0+84bdmudNdffbe5OLypID6E
zHpJAU508RB3663rUDKsDWClJQLBt5XquXSdzapbW8yVX9A2pfZIaeaOcvuhZBwS
YA28RjIfi363/CnveEGZ0bj1qRJ/I3/xqdaMpnYkjCkPw2Xxf4cxrO9XbTXnfemm
NwhXrz6xVZP50Thi4cVBKj5XetdS8RsLiE0BsFif3CId00BC4D5W4tNvq5Ev1nED
TMSDayM8ox41KpL2Bb3YtKlqeJuUiKSpVkhb66q4epu1p57y6HfpbXQV45iOcu1a
64r08eWiJqvZoxGlzqho2DhXBexBJUwKOxsT9Ty5vTjfyG94pOmkj+2d3feHFkFC
oxLXM6wTXvde/Y9cXy+3kifbpJQAbX/uV9Wt7tL+o3zyeSRPNNmXaBDjPboCfaYA
okjjc+Ost73ouU7fa9HwzcIvqvJ0+ms8Bjwr6uELjdekCedEPj5onl1HlRyLsqns
Va79C5EtXAe9hAajiQf8JfYsl21ZGjFfbnwq27ZOacrycvfnDfKN1dByzfheCbbL
3dgMmI3K9DXMXxIqaU+AfUGS91lN9l1K0cLPtFkAY8/jPxodjeCGGO9/ukeWYF7l
6UZJhRjXhAevhrT+8+ijeZkzhs+CtF5VzwN4M9rWIc3WhL0xwGu2GgWl4A+EF3dO
AxyImXyCujh8fykwOcD86p6uH5CYbtX69mo8CSwLPkr0YOIVme349Tx7kjhRCBUO
1ERJtpU47QBTHdFdbob+ixhquUjiRyc+xHlCJkXNkylP/I+moynCATK+fUEk18Jt
XZjQ6iQc8uXkaCOTIV3IEPz3/MLEWKGai4UsYg/CNsa3iRU6crBRtqDzu77EmGl5
3a8SpAh2btOw+3jmOk64y7cgYj0lEqmz7JJhJOBpWzg1POzK3Hsorx/j6/RzEHet
AYB8Y1IMlxdTR8HR05aCIquepW+PglHxdNktDAQSjYf0wnLwTOCaVAVhyu2jbYiM
yDLQ/6OtbQSulfiIJ2dlxDmnBu6zPpmSNWWunBXgDTLPlbNHLzHI1YLNBiktStbm
WQzGH3NSt221n0BQO2TsSSgMD1Y0d1L9lcHfpN9F3neLWd/WNJ/pgkEY39aJpVXh
U6goxYCBelS8hrO3wNWvJmtin0RgeEIe96M9VJCIVwSYhTnBrey8x+xpRiyPwLyh
+5rZ7DXskw8sR9STBuzILWtPN+EMnGF6dmTN1ytOnoHJlU8vXuPTBRVOyPWeOLWQ
KOkzHvHt/T36yaoDJmocpSojkpcLO+YHBWWlUao3+oMWfL76FK4vMBxdLuf+1Vgj
zA+iixcD3Ohd4Tc4y6W2q9JVrBKyCNEJEN6ZV9smAqTW8rau7r5BqZb8JSaVKchr
xtrtc+LVn/1Q0PAimBI2QXPslnkZFJPuGLLV6Hz9RkKv2bV0ZNL8HjwTuBe3oiqV
ilpKiCHi3HI6v4Iwy/OZ5Hr3CuruQaD1fakLIPqC9zBrJ5h/3J0oCEhdBqVXS027
hHDYjJeFlfQawKUoYVyRhH5hlFrYD0edsDPD4PC6hIv5UUBbRyxi8cL2FMUnIQUv
JuFjEeXwGsJe3rzD0+bAk4+oA3VtA+3dO6+Syed8D9QXDBq+SiWH84Ofg/ROWgNg
eqRnEq46qAORk2EFPgtqGiQt/SvvBG/kS8z4A0GnwKxl3efdbSUJ2sicOGtrqPr7
tD0UixYmoSD6/fd329QM3amZsjrVqYKRZpIzDlFXHxTrDLla8iLG2rb+OEca4KZb
cY1yWxZPecswB7rKfto5/0RJzOhVJ7oBjIBzNTWrvJGQ+GQMKvMN0HWg9phq+Dnn
5vX/JWJloVgbPVuZsUfSu6Cm4jXvjx1FP7O07+lqp5Uk9AApMUHHOod8Ogtw/Eq9
fUCbm/vKJF4/c51JzW0cc007upVdHle2jFjoZpC1vaeLlv7gEK12ih9iL1V5c4Lp
ZJRe1hmo93Psy6q8yv1r3E8dIUoIvoeR6AZgnI8+fwCsEavcllQsDqUrCofndBSw
v0meZaiuDA8Wbg7aCbn9Bf3YaaHDxXI/TL060JwLVRw4kDwRFWf462LhALGXVd15
AI1vzeBZXkyw6TjFXkaBC7kxL/oROYE/S3sVZOgBa+dBBjY5H98R3GJYjESkdVeF
dOc0Mb+Vi9dU7bwOqpwp6XFleJVwxu5qcfSggGU/mWSs6GWya1Pe8z27qbxicmDi
zY7Ira2yoAP3iJ9FHn28wCgnk7VgiHCeo+dmh4lOQfxSXRCdlY0s65BPDzaYD1SF
5PqVbqI051tGNoXG/Tj7lNdA2J35zmWhInLROdFzhuTaWCcL0vIGSnl51w69/u6n
Z1uB2z10e078vkr3OI21/1Hhc5kxNIfZh6DxTbtn8cPwWxlewg8dv2xupiILPflG
W36qRgpjqDfsw/gIqGRKnf1h8C2GSf6gp9gF3xsdgABZI4pWE409ejMUjuVfCg0N
JOAsBKUyRJHMCrXOfLOyhYzb7tyKqhaHknCdy+rbh6rEZhdxMBJOCywlFsQVYmqF
QH936mrrl2jFZ5WqIZM5wZDvAZ472wCKbqwN5M3nFuXSb2d/NgK3QFmqChv/rZoI
7a6qvfj4Tbwgq7IZZIuSOWA0irHlhw/oWktymuJSufg0208EZFm5+33gPbMUXY3L
LJdYJQNTGABhlHvr4kWUBMOBgSa9Rmb9ZKkwkhJO+CEi6oAQECdPplCsV8wa1skT
6Gd731eBqgPJ2boVt3UvJ5rL13I+rGfk5yZ4VDcBc4D1XpNEpAbwnhaNcJCmcPrg
tYWgkarKOhSIbPO89aMi3w95oaBjh5QE5x36vd/QmQs4lJOaMOO0vVbteV5Aa8qf
YdKVQlF+jdHoBBzXZkKL5mtOabZldNj6NslCI1t3aeavabgEkmthhuO+fOSmmUe4
bhlQkUnKMyq2CctSo2u0WoI3rPDLSuvMJ4tnhRL9K3SDKb1fERJPlZEM1gzrC8HD
tjCqQ++rvWwLRU/FCeP2cDyA3i6L40dHxcIO6aCXVcc8B1UekGKIN3WL6d1ifPto
OiKYs1shfMHPgVt5lE8AfC77T4JkNIZunhBZjZWTspBc5WmZJ0XDEHa7K/+z0eBc
FDsiqoGPojFQ7lSY/j6KVoxrlh3xeNiSffjHOiQ6RKDugVjxx9BWFzsjWTh9c0ig
euBudOLxr+MURQGZDM2QLjvJY0cv+ru2foa4VASpoL4xF5I29OvsD2dk5IE5FZ9H
G21gzrK//hAkR5e0u8ybJmX65SfLeJcPEtPHgiyRVnksdztMVNEtC4i3lchv19YV
SpLOyhslFCbHpRHHqJOP2C6JSGTroezONYTsP9nIMWo+zfe43K7AiBhyZlujit4l
aoh18HHxScJuQYgDksoMnjmrMK376VW6VIaKnpmQErCaZA8Pd5OS5Sp+fN6pDOa4
AYZ4JmF3pJQewiOQw/d5IGxGeeY4KXpJ7ZlevuqaWEzjfZO+w7pqHSdNDzBPrJuT
8lNC2dRVr01m0RyU2BlwNT3wsIkSvEq9fLNna6/hgSbjnSuKdcWY/F752ozLcHie
MU4hZyKUVj0L9cmfPp9Tiavkct+kZNyJlYXtkeZii8LGh+pfscMSr2sGM+B3obBv
M0RnAp+5UGd/bM2vyTQ8r4hbjVl0vp8u0UTm6GyEg2n3sPX7Js2nnw+q05hyyynb
iQozsFXaZZIUj1k1phK9SoavCHFqy85ZcV07YcdG0Aa3fbZKiq2FsIaxzrIcNo60
RaMl9hibQik4RxfHoT3N+0wiXY/OfwUlVusNXUCfyU4yyPFRCU4/XVk+MBUCHK2d
cYZ6/GSFwTc0uv3O3f2ZAtZDKC8U6pZMtEeMyB7FTPcCQFvHGGFbAf4UR1S4FW9h
6yVkM7cwi1fSk8T9Pty5PS9u5JDu7K9jNuT9zqQSDs+8mZUKiIZONRK1QbDaFkjR
hJpNdGyUKX86nCIfdsVSyRJGrIkkJAqR4rokTHKANbOjkwfN6PGQqR14dVnkNqhr
uC8wdEMCUDSjVfxB9eL2ZxLkibps5MJoa8Ftaj4VjQ7N3GVo5pClhk+WfJdIyYDG
+C1Yv3AX7sXD7nKSXm4U4zpGf2ilNXdje9J08tFk4qjaDiI2GV/cf8xMijPqXVy0
JXJSGQirqJg+10iIIrnzOk/5byum58+1B2qaWE5xAwpY9xGzcVmciKvs/j3F4F+T
VuRY8ohIa1S0ZRWwqGpHcBeCUBXfFiJn8xo58vZr4lwDXruF0QzAs7LjImxWffTD
y2ZByCd7Isp/HFVMdW4KPAbWLniLVtXWnETQGqC8EAQR6MfYk5fXFKPr748iNvo4
ZwmikMB2Dq1QLn6aZff5ahMm74eQYtkerctoDJbRhepQFX0pKrnHRtCVzbKi3KkG
zGlsGWfZUSWeezZmKlWjv30OXuLNmprKsmHg+yMmm/W98X/0TRrG7+q9qAwUMJaE
oY71umlyLVli1iFZ/QOoUnxS/vj/fJPEiBU/jIFgBGW3dKBMquWu5hHQ5VIF7p4W
iwg2+vUSd9zYzfpxNTRn0M4/BxHw2f+5MDrh9+VsysBIiYTqTk/Vm8txwlIxuApo
0HSPIsjm9cqsTJhjmw/wPOUchycPV88Rgb4Ao/ToTb8yGcKfvCGNviQaDahSA95C
eqjSd8WgbtR0oOu+F0n9oJ/ireMB5da0TOnv2UfF7/Y/vmojXzjADAAmwatb59Gm
aQEijcuqDUl+TLhkX3pNQK4uV4Y2CuXbcJ7rnWXipI1aCYNLnpEDTM5toX/vx6GL
PkaXBdaMGhmxPH5/CFkCxB7eaNorumn7z+qkyOGzZKRGiZAMSKnF2vlB3/EnuCmp
7FO5lmQ6sACu6QIZKSsripjndEcykc6bjq7ejQJt39+gMyZNRMntGGnJMUuAgazq
YDAc2LcAP/ClCRf7H5wkLZVCcyoLVCv95lXbS6vqn0QFcivkYzLRHH52zOduSS92
Y/veSVfPowSD4SZNL29DcosY8j+cETpF6fNaNhLgkvN+molWia2Ws8/vhwY9YrEt
5Js1lGw64/gzyxmazz5q36Iw0Z1GUKnTcPLyuFoYy9+HqYsUR/jA6AwwnZTQTkIW
mdt2laXUMjs3y9Ow6tp5Xv9nrdGVdCz8qURbrIaL8TDpEMPQuDWj23ScunDCjI3O
zU2pFtTeVLyLNIMWkPLKzHN5D7wqKl/JrJBFMFN9A16vBE0qaPV45uXA5reug/cr
GO6QbOerF19Sq8sFtI7kLRTTnHMZLLdbJU7zsecCw2IiZlguKnfiZPMq+ZybEM/u
/JIlw9ZwVMDqzS5FCThWh/wDpS3E5O+1AG0ticzhRRWtqw1vIZ3HoiQ8OsXLNeFP
gBNGs4YYq1aOs72yU3/4hTI4VRQm4M1F5RXZRaSws2CMoSef11NKrjLBvZc8M3fm
szt+zKT/kLtuUBBxl2NsRkGkjpP1ExnJvqlypJkX0OAkhlohnJAv92OEWxuRMKhd
6PXSVRRLr3RhebQs9XVJwcIAauYqeSkSiPOn12Gqaqvcrjh+AUk/GyCirKU7EJ48
XFL04VH7IOb2NwzIrttuAC6sTfh+fEUvBintV2XjxxyOwRMT0ia43NA29vY8/WDr
K9V60qZ6QkWbRE5NlDVnY6NkCATmWwUYUasDbu7wK2K6uIdXqAnMSva+nxeWpxrP
Z3KVL3qXFsCmdHzMjlllvR0JoQnmJjBo+4vzk23s7wxEv7tZWzRJG/WAq7OW619I
0fHsvEAH2cxrbqUEPxJYZggHqberoSXFac6XeeaU9l8OSdDRSDBeTjZKrKkwjagZ
/hWok9vRWIMXxVISpo1CM+42CVVmIqILnWDSS2D4IYvVKEuNYWMTmFlvu2DT3a6f
eGTSZwlnqed944eCzSXsnXVWc+heXXcak/ZhmOMu1G6o2ND4yn8n8UIZIScTIaza
Gr0FZIgqh8QntmDU/MC8MRTEqmcqZhhDH72aZDgi3XeNTs2Yv4KxtmdyFUrmtZDQ
JlSMZOEe8HtOzC41CDnZM81/IAdQaC0G5hMR82FbZVzotCUftivlnhp08CDQfQKk
3lhp2ZJ1pDvDXnyyi4gTOMsFgfRLAMPcskwiU7BW2O0kIAW7mJrxJnZ0wQTQAYLt
30G+wH2e8F54w718egntETeD+M10Tf1N52ufx8uRSPQW1ETkmYulvjmnV1HaqXBG
uJZhj2ODNb/dACn5Pj+ErcLIBAbRzFAFzAoFdZL4X+1vrZ/3QI0Aki/HHzYlJW/g
/vPwOBK2RagmpVAILqvcZtIZuaMXJr66DSZK72erc9dvL0X4Xo67XvA6yMLHqqCX
6YM5UkmQuQLDUCHZBtSNaY7azFbf2Pyhumn2v0v8ve4UYsZJKu5Prdu8fwX2wkpz
C/gNgHRp2YWQjahg6R0DRJkaTDCnwbXpueXf9ZhRQyDBZ0yVcojz+5TumE7GrNug
/peBdcarfIrFwdC7CtsF/QqwheQu0OWDrzKUiFBlI7RHmkhwk+Ul8EK+BrT9xLtm
16g1AKiJ4W8EGXOiJc5FGIOJNFjEKVsn27uUkwm8Y8ZwBOQRoX3PgZVHvUrCPq4H
t/yQfBjGG+FbTYC52/PBY5SFqtkW3fYtdDhgZvPTvT2MIrzPwuA+47u0ZQDeWNzX
aGP4NF14bJ/mVbhg3E7NSr/uj5otwdKIzcxyPLoRmkiChBwbMNQMpQ+hCvLfsam1
1eeDS8MflhH1iUYMVWtBe+ISjjW8Q8w3pWC0iYmeSsGRcMW7o6D+upMU69QIzk0p
dU+UA6MqzU21ELo+vebW7MfAP7biaZZT24bEFxtUaUDqt4yWJLAe/ghc6ZOVefUU
hGDAsj4tSsScaeylMdSW44L58+Ca8RdhY6pcfotxiOVjhClngg4F1neFardw40T/
lICffCr8x1zRpIlcJk4hXRuC7OLRZM/d/dTsg+s2FD3KIyso2wA74Rw053zsJNFl
mfd4C9yX61k7+dyKJyoEEDJay1dfhIEndURTW3ymybZV0y7BLgm+tljwnMTeuW6g
WbqeDlEfCCePNwbJR1t8fC2/j0YP01rjc/MhKjThb73EbAe75zmnVkPL4pkhV6k5
Oib6GWtdFFe2pf/9OenZEDYGvS/N2J5jhDT2Te2fapNSywTgw9S6k/h6MA5DCklq
1c6OFfVRSMzU8dKEZ3Rfevxr2LmZacxRHp6vxZ+0OaFnCijS0RFHBOyjL8Hbeig8
LIeHOcqOOgS8BJQzxVWPH0zRw3I8dg/xnre2LLJoE6KxjORQJzH0isYb4iGDWVQ/
ZfQC6FSUbcYumTQBxh1i0qvIn0YRHQcHTIpamarBuTgJ67W9ZbMgmFegwXvS2pHg
WHhLhG/S522a0zfXAuULRSR8p363KNzn/NpQwUwvAPYJ2WZ4tBdSVLX7ahLa8QjJ
ahAkHo7cbPUXvgJzI9oypGJ7C6Ctp+QRxRXm44EH6f9M8NrhKg0BqEpNvHqvLkVW
6PivOK+dPCbPDyCAsN+mV4FijvhAGskzH6GnTaXHiN/HriOaj0/kNefiBxqH2XqG
UnOUmEhUDuSLPwq/WLrvKe5a///Z9K4MEDCiBIl1UGQv2VGNNcjsRKvtOV4gVZP9
czlX52wQnsxZ1E6XeqOzVAelv3me1XBOU3bw3xzE/o+GWESQnVyR2g2qChYNt97N
G0Rg4XRjtahPpOflIA3q4CZIqj1lt0xRNY59nLpgIO/0JJGZqa1JCZDRUqXco5Um
aLu6tE7CP6uVc/5yZqsAGvLfmCkWF50G5F1ObBj+zBvge55TQJGbnsBC0LUHDeVJ
CY0znxwyDmmO0XuYl22W4SaAYfYfBBLf4X7Daw0SOJMxW4QHvmM98rvGT9kb8IJQ
5G5p4HLdw5tD2iEAp/L4eSw1IpQr1s7+1LM+INJYwzOFPew7KtnEY0elKF9wAyxF
3BfQFhpkC/fV754uynNU07zEOmbRlgwMqcbs4El4B0dHRoRJNUPN7l+yhgoNOqNg
64s3Km3DAi8URlxfaHB1PjohkK8gP7DxrxDmu/swUwr0zrQKBVqeY5E6ROFxftx/
zeLmj8YlVuoyvaRH9zWpmTcvzTjecgOsPNjNT6DK0VhZTXh0wJ1HA4D16DtfrFBA
iZ/f/MM3mJUOkyMu0V5X0VG7RLgfPY8R6mF22O60AyTsmU5g650vw9HS5eruNWtx
PHeKpSv5M3Xw8UusIoawSkd1BMqd+EdV56w/g3+H8G7tar4sG5tnd9Y7t5VRAwVi
TdiTv7DNqKOotpcaeTFz1KC7XMq3oS69kVLCwf61llhKKzmx/PU6g14eO9bP4nfx
NFJitdufU9rJNaZr3M8VqKS+eSbPS+lrwWIKAdU8lij1PLIixwizbDgDqUnuH27z
iaV8jLPZSl1SovUTCQFvONG1Z9e4z3WUKd5nUOrmjE/zNU3Z7A7BYed9cnCgX5bX
mZPE9diIF6WRcwYkDti6RPoVFddRyiRtg0izumdpUDsAVdAAuwPe+JBY7sRcSdVR
tYkhPAq8kUyskRObJVMJNlr8g7eH3kSRrV2+6RnBDeLbI/MeronMc5vFijDtb8K0
QPyphhkxZzDHGBEH9+bvZ5z5OSzJqnAtCUktuoiSEin0qzjYhdJkPh9ONefux1Eo
bXn+jPKNuYmcMRom4i2tfxBsYp+lbSjB4VqhhQX7kGaFrQNnYpFcrk+ClZYzTOTQ
upfDWGn32CPOUBuvT4Gr0qNf3e9VHc7ZfkfxPGrTjDNXt/Q8x3bSFKtQnY4bMsh5
LSTnp5ZUBB7rW/r7BKhh/wGBHdEMfSXIrnaGI2gOyLqTOASiB0r2Ya1GFEB9O/Ys
1/96bzRFU+s289N45MvURPsBgGPrBqgwIbDk+MX+ImgWuT1WVJwDAm6AsVeaGEdU
j4AMz10vbrXQqLEGt0FTVVX1lslLitLRwRCspL8oMU5Uo5vPFPycY7Frk27WsMyD
hh07kvwpymLARFb0EoSThfbEQ4cjU0Y+fOhXgVeWuq/E1cwjM2nEoK23UAP/9eHR
mGjKH81ExtCI3qI0Aub+3cCJyLA9FzUjy2dVKl6uUe55S8Irvpz/iS7lqU3+wrzr
6pHxRtEIH0612EP5sdeLRD7SF9SWKaqEZgiLnD27SG4nzQfbNR513NglQLhYCdFE
Ec8G75wu6IrUyqQ9kFi83QqdOidyhTOHnTnU2UmXOtbyL0a3Gpgb0Htj4If6ZovI
GAtmifcCY7bKcJmrGe20vvHX+yQAqhhna+fi6JjVB16e21OGdA0czgJ1cSjmad5S
TTG/5CNNvv4xErrFx8i9VyQxG3vrhgHzGl3f1tOb1cdsXVWP/ARHTcI978XxKSnO
NGSb2u5mOHZGebFBjy6s58zj0BaccTFPiXTbNyWk9R6r9F5u6r9MyQMAchYBF/5s
TPoPEhwnL5DY5fn+0b/zkt3VFCkJIWH9lDbtnxPwvRp5z2dgltOtJt66tz4oWByP
nfY3iz25n9aqOIRaHYDgrOtUoy0ABkMDr7Ac+bntoz1ppbFH9NBJE4UVUAac37c2
JuuKhZqLxlgTYC+4rwxsmhets+j+1Wbfk527yTvFrfbAwIxgl9YFArGsqzDuOPLu
m4DD83CLvCaJSlqnA37CJUmzLwF4wezQYUIV50cxvr/SM11TvZBwtToo9IWxIJNR
N4P2yehc8rYfp5e7b1vxfky6CNIif6kFTiZ5mG3c07b27LsBN7cA+L9E/+ckUrQf
QTpbmEiPPzk/8zxUJRMdvO93SXMI/XcMK8XoaEJmrG7xMV2yIsT5EjyE5fcGJSSN
tZ4Oxxgm/jOv7PW9H7Ov4/Q3CRoH6jUGr8BWeCijGdaBppYwX5LLYtVssBKH451h
Mn2XVcygu3jsw1R3kCgEpUZjRlM+1U05zbdRY59GZj5XIhKQq0owsTgxmBsCOLdk
8HrcXx/aJFbDwotpZdnNyArCeSTRFHbyAsPVKdyjHHoDddbfnawJ/l+pMk1nJ+ub
HXCwcd8ugeKdnYXYl+BU0fnyJxIaTZvay5PXUcx/liPQrTyFOkLl0G699PPpdRPT
omV+LuvXUUzAbsbPoWSBclq99g8ePlFh7mdbbE2p0lLnIAEWqvEDSZh7XGPZ9/cZ
jiyHkGyx8aTYPr504GaskL2kYU3cuAn1jMeLp1Pc/txcr1FTI5tZnkOw2TcYaCic
vmTcn6h83jolyMNF3DSWe+UcK3pTGuAzwPqEVoBzO4FieAZEKIzWAOyeh58F/pLP
REbUruoedvwWe8omiTDZCTp6oh+3UAy/o0tHYuWxk8ZWe9NjUTfu0GNgZBQy9b6R
HBOT0q0If4jgSf4L0kwAL1QmWAAIO05c/IDL5t/CObSVY3K7E8f3eYnHQa9uux1W
qkSv6GcbIMQGt6kaowjSZalm61yEzds1wE5Djax2loEjrGNeZeIga3kirGtPJe0M
E4eotTeXUjcfqtmcXZ9HErHaKa58C0RfIXffAgPdHZFK+I4IlcEW+oJaV4Yk+reg
8KMrGQdubNKnKxK0f5K0a9MeI60HGtyUXoYCuOXGdrR9P/XbAn90G5BW3VRes6BR
RCUohiUe51c6eZ0a9Pe8CI7cF5lwJlAxAn0NC6fEa1uhKnqV6zP5VHArBgk2HNkf
NWA3i1TJeJNWFf906qkoJX/vNdArM0jv1MTMXNf8vuJqC4TN1O0LMLmbFE00/0Kb
R39vZ+TJ0pzhdeeDqNK03azhph1F+EIxbDFX3Xk+MWlYkMDphIyiHuhzRL49gcGD
yjabQW1RUCF6JdYIv7JfeX2A0nEavaZIbSiJbpzLMSFVEtWfuImPIaV951EtSXpy
pLrSpcc3Sv/R21bJQgli+yAAbQirWr5fQHZf3OOP73fWxGezI6SKqddgkwt21oHI
ruUrlhLCAxeKUOuxHb6avahfk4b3rY/IBFpWZ9hJdG6GGY19UNc++CrWAE+l/EzT
WmjGSgi76GMKmh7ETd2NZVCairYfMEYTveMKCpQrHUTdGgWC06UpS8x69lzU8lVp
MUGd0gZvpjIFQgNEF59GylJTLbtgRC8/KXw0KthJEQ7yRCluTvLr220LSLTSkDmv
Az7jd0uS4t6rVeKSQXV4IlfSHmIcJtwi4E2Sx1TDV+aC+rMaPE7pIcNc3Pl294X+
K0F2hKFq0kFepitP200Yis7ri6VmY78A04WdtNe/iIanek3HFBQVgbTthlKX+pZh
tr0UAUqTtUR2Y0EA4SAKPAAhplsnWnXvf4Yeos3C5zJoVKDbq5C4swANexfVe79s
BvGiDVlJvYn2BygYeEWXXXDO9ntq9KJiNsRMTqq6jrQ9CHFNFVjHZZxZGpf1Wd8d
OXbnjYlw+ulhvr+17nKJCsnohFhWBvifzETNXIPkTx/KDISLIjpXCqy7VN0OjLc7
1kOaFp+ajGZBdjBsi3iUj67fQrVgL1SucZ+5lGETLRXLxtReYVm6X/odhr/shD3d
q0gIU2P4ERYuPZJkV7ALcFn+S6jZhT7KEyjNqzrIrZNUQvK5iMQ7dMPTsd8IoVsp
1bqwCU+MIY/AFgmq8w3cpf7o6ag+09Fm1L5AqqlzB5kgdiyntJgUzc+xLespBDSY
z3UXKRxpOwrz053iHymsafhI+1ChLEy1kl3xFXdAPZQdkmsM/rhjK5mBKhzj4HTv
M+YmwpMyJ58RVnO7sb0ncqHJ5mHxvIPLWpZHTPuzzfQhg8Scl7+d+ep1o0Mb4+iL
0/B3THCGulVir1F3chgo+4VkfPmW3wfedS2Bhjv+9p+OxCPPXjlLY+vo9oTV7B/L
ufofGuaAbRmvlIdhapi9IgNVovmhhwlQCKxgW1CqzPmt/S5z+S/BKqyv1b0Bm0Vm
gb6MqVTAxkVV66143L+t/qhY65WFstklcutgeF5UQCD2dkK2QKfAR/qLK+3KfTkh
F0777A/pc9NcxlHup+LfU1lBaHZiaLEL5XSpjYkB42sz4uwHvPukoiGVI4cHXnOz
FjUw6QqkEr4soV8ciZ0id3qDUykSq2xL5IE8BxYDTHjwzVqkHJCCd6PV0towDpRV
u07HYdL0pyab9lAbSsA0hsWgfqV0jtVP+n8tmi6PzhLVYofesDb3lm+rDdovY22s
gnvYWW4v2a6ZK6LGT9qZUQb0lAxk6RvRoQJb3m5xrxEme94DKhoWJj9/jX3Idvjv
Ps74EXW3p8uFfp/gulDcaU8NDGS2xr5T+zIy+6isYrETD13ZLHgxXikhY5Md+zrn
roa68SRH6r3r3afnDBMwRx92kSvtt5JKjnP6aKsZdTPD6AHplykaL4SRZY3SwbdM
W5UKAsY/g3AuaDbY56dvnvLu6zOe6pXWKSjrVqCJCk7nrByM1sOQFvzh6AixyqDa
UOOPtc5xndWF2fvoNW0aNwfk0XWtyzikQ9gb1imw/OcYZUgCZdNvJI1UvqPYWYJm
SBb3xuGJFdnlqVh+zKCOBG/wHM6QpncNMA8exzpm1F48PeUdRKD8ukmpKdD5HmSi
ZjbO2BqLZcI9/WuVxJnMRiY5wVPEOSQkuC35+GI1sSXzjy7vS4WpzxCTuD9EsYe8
e+ns3UZBoaK5bZAjyo2/6tmK+JprnbdYX+lmeqsbVZ62NNjT3gA/ytg1TFhEg/8F
qW640MFmzqHYjY3yWYWDl9VYhdNr1LAFntL5UutaSIQMnDaj2QugDKtI/5ujRIGv
aE08G2uEYe7AmwWbBapcAO6YgazcBlkf23CAamSu49x6OTQFAQ6MLYdZ5HR8e2Pk
sdlm5HFWd6WXuwq8RVJa/YafwLIxWfKEkDHo3+F2dFNe7eWCZlysrTlhgNasrxpb
dJNeB7His/jIBejxwLy7wz02Iba1NTsoZylNzy8x4qUnwyiToxh0NLxJTqiHt+ns
KsuqJLXenNIwQYq/3odMg6zsw0cZsrAhpXi4FDCzrMtVzdUOgecIsUvwJhmNLAJp
PcMX88kxdn+auZAZCcbNnD8IabM8I3xh76ODrngZ0S5O1hCzhIZXlr2PFnU3O0Ao
WOy/TPquUlbCrApqBdA4BNdrjSip4yUnAwauQv9YEKDNcb11w+J4C+O2HiMe9ZPg
f4vQGVE/sxeUVIk/NTIUbaoM4AyNBdvcLOLptVptTAqS2FnhDZOAnq5X6RzbN2JL
xN5U6vUrG0+o9r3oAmWs29UmkJoO3uHsDBtGF7Zd/CIn3V1htLC1xjcyrq6lepSI
b+qlConv0SBDciDzrTy3xot4Yej65rWKmAoXoTsghWM/+e51ACcGSb7IOjtFmcj7
kfHmNCQs5rTMqHthIaTWOvllLjXr6p83LIeLz5R0aW8gSg1nATkGmRcSQdPbPWrZ
HW42FXgt6oDTHnsybOOTt6Hba5s3XhWBh8DU0xof3H0d0rUX95XSxKJ2wRJPniII
qpTphtLXt9BB2fM+w3aG184CHwOp3F4EmiBmWWNrUXOGZ0QdRTocdUWu+gxSXbG6
/+pwFj4oMwc3OXfolddTpOvXDaF34QPMZBE9tIuVjELEbfsRLdB5FbZiZ+vEudo+
nI/xwyXTOo+h7OGF5fYzgExaKwfzgM1kaTzwXH8a0bi/+aUnF2wa0YmAI5JZi0WM
nIBV+SkkfPUOTh5IxDO0HJUQpDVXtlr5pwBUR0LHmIeWoUM6Dj9cYoLBoVjqjr43
KqUgiExsJAAAm325KO6vdEdPnd5G+6cAMeDClOiTc0H+yl9mvb4OPPXiEuIbBB3k
YxsdJOcwDJbTMCJlOsAVbfA7wBbj6MPMIRPmdFQa/MVYiJ5TzUi4JzcNY3YwsC1r
CpXhByFuufKpb5L1ois6m5jPAndnseuKdaZ1Sn403KmxzWiGXtlkX9qg3dkLKW9q
Y5ncd2sUnpOlLwXm5fa2UYOmJL8s9iaIxNNgAethcMj5MVltCVIpH31mfRxZQdWU
8QtsAOvuxiJVuzL0EgXkRyhw/4UA+CKFreSQw89sB2XK4ZXFpfNIIKDGroLPD7AN
jsE8mvteuOPBe5ysZ4Mlam+21qXPqrzsg2r2tG/aMMk0W/Y/R+sDJaus0IxHd0RV
TmV0lvvV/t8oYDmBq8+jNhj8ZVhxMG4M05sLfSyxOA6yl6fPojvtwBrFZ74PtDYh
l0lHNL7a2U6XFtoG6V5V8X3n3TbLfhAVn1f3TEIA7rbTrPjKuyrkC1jsrM2kiN7l
RveCJ9CtEupdIlr5449Yun99uIz5/VaC4GQfyqBE+sl5NbIVHNHPyhNW2CXUqIbu
rCF1lzFcj7z39XQHWza9RIJ1CyiroyQwDPvBwWs3zCkVjaJIGVsWWXYEHeQOtORZ
7E3FRQroLmUX/F04PPrV0bYzkFAogHXK/Uvp4p1XEkcgJ+d8FMIWiNcLL1a/8pRw
t8BaMLerQ9dzxG6xjmGMscROECEjjaY+QHOIiYIJbZG2AZpOP5p5lqfRSP5b5A/s
jiu1KD33oIiMcc1TMneL3/j/JS/IK4aZ6FDtocgm/y6YpWW9ZbIxn/v0+2baqUcq
vW/bgPWN5G8/j7XQdJ6x+tHZnVUQVKqvAkGB3BubA2o3mkZzwPh1ktIixPlLXLuU
e5HtcqJwKj+pAN7bYGGSt5tVXU66vbTI7B7WDHjmMRKYKWXgp/T9PccPpPgoyudM
tKP4HKpcbJrqjlcnhaafWNX71udSLH0XsQiLKHFSPWytZvbpI8llBi+7xW2718kC
ltTgLeYf/dG8lxkDqQ/5PvG3MDIYhOT1BHBIBbd0D2f+e6369yBIZnaJm0LxnxjB
x64sHH8mPCSFfjtmY4WG9WgrlGPn+jaW7I5QDCiOgMlmUq7/9O7zM7gC41n0KaUu
v5T1ERlTGJzRRYfjNGgBqEs/sIdMJmhhGym9qd2fMjiZSeMvgvhkwlm7+Ti7MBWx
Y/dBjO0xjaLKmTMFSO84iT01/k2i1qBGafceGr1D4Z6Q00rdn1nV6VIBnvO2Pp42
Y48+mFLW0PfMcP3wC2d35qjW6244tq5QOKnV/pVN658PeBxMrmEUHzP+/kWUDCL4
NpfJ3BiKll5vtzNtKbmgI82i7WJ0M/gQlG+TT5Z2x2zGHCYeERjLuJlRXnU2WDEj
1qE8dM0+JaimT7Ni9o1XemnhubNzHPhB/yluFsCCw3xc3447J7d+qOxMHnCH3kVw
jCV2CTeUPMEFXnrcsDkCDdu8JyH5KBiXpy1X2XMEWYVaVwCCGLG1Ii3OY6ZX8K46
ruZEirtP+Pn2d5bCVdhFk6s7ap5X0kt/FBb37ZbSCHUKp0oieDYrAoa5MGHBM+0d
5FmSHyX1M+OGPqyb4eshjJk7c16KTA8x19e1cMZGBprEPhca9kll9v+T5+iG4JmD
iYTPQlqiziUBeHokjgnVA197ejKy9STIop/YFmQQyzhbf/lOQaxrMBTKyCoflK+6
vrGeoqEXhjYivh72i+ZdxjiMERK1lLxsUX6kEUwhxKlJK++ulD9m3adZwGx2X5X+
wiQs17BQ1L4jbMvKp2o7UnWZpIT0q3BEuYYK8G4ZrCgdzcQ75UZUB1LuimVqSNPv
SVGoi4+gZQRAXAnJZniTlIA+PXKf1Y4X3lVwQfovzERKjxjGax1KhTJqM3pk9ebx
g+9SoJPiaCQn5HieI2ET+FIFn+2csDq+FooNmDJcySexezdaGKx8igeBxjmtX7Gl
7/xd4wPc3UrtkOGRlZgz5lL4vo9ivzq6yOHVYeoUMKh4fNj6CCZyBWN8wPuVIv23
jQex6lFulUrti270EC7Tes+OolWzoamoEo99MjDX6+OVJipNWXJS7GQEl87i12au
yxO5XpkzMM2tUqPbuN/a45uwq3UciRcek4r7Fp/BZiZUOD3jq/sJjm20mhjp6zeA
jzmLIuCidNwnm8XEbj11M/xrt6tCkhtMEKtPYDXmbCXqkw9/bbfonvcgcLURzh5B
cRG/UO5rRujKwRsizjroxUlfjPQBGlMh+j8GvSK4rC0nfc6qvxJtoEkkj+otSifc
+ERll0joCzOXFodgl1HSBSNy/a1E6LFE34zFuhnluPZ6Qn8IJcrisohDwQSkR1I9
5si+CK4pYvvrpo0P72WUEEzslDcVFPcgMvHDTYyww1QonNnprNmhJyVl+mjIGlIl
wf6ItYEvdlF9EUDl9YE4HTNjkJmvCJzsA5ksXJLieJduxlrCJOOSPLSiPW3x6Xzp
Ku6T1MQnZY69TI+Zd70bDVlYXCyZX9cPbDWwzGWxbKhgS+ZQU11F5FDjckWLVJ82
n4Or5wvDZ0mkm7pjKxJ7U1Ol/VK8tnBUGfbJuo/uY7I52lSJlKaGyzlo6UctM5DS
aF5I+YehWJ9Vx2WGVzoTKVAOngCqJ9soMpr2eOk9wDS/gn8zupSnf1w+wg+AhaA1
1Z85XURRAlFEpMXavfhj9BjwUfsjrB0gnGUE5ha/M6rKiuHyAUgyvHTMLgG4lP27
uyvLbH5s8aUAfm/OwAy4wewIZvnSmKCH4Cx9IvqJXEnh44xEjvyoxORxOoOFXk3y
I5Un6KLho5HzpaZS4+gSKUUWDKxIMUaKFLbKcsR+2kwwpXtZr0NSJHZF2wrGjAlS
EaecTY4SQXhbaWCHGPsgOi+BWAtjZVzy3BWYtHi4r6NrQLL7qrzpjoG7ZNaSQAvN
WzO1pg/GdYUMn/X9aRTYQXGIgiZ0sGSxFE0IEpIWaqyxBDb7SzEVkqMcTKcsf6gU
gqnAVBD0dqbhcT2GkKPRcNWJgMDVZ8yKlvI2mUvJNI8fOM1R3CiJfPuZBSbXoVUq
ADbrwLS+ytSCq7e5MVdTd+Olljq7MIHzNQfV/08GT92sXM33d/HHTDKkaR1pI/2V
gazrPDvzBmPp4T0K8QWbhTyJIerJoM5P+9CFmLXHZoIKIDvBMpRLcOBiQBNBEBlY
iY1svETLHwvv8MChKrA7jk+9HGpFJvp+a6MJkfQ06DeO0IHPSo89x992wd/AKZNb
t0HdFZnRpBDF48LyLx0i1WmpfHZaAdOt1gCzJA51yRRAa6d2DCTZvfsmOX9u5IWi
cSTmXpWN72hpvm6Gcx3vuaomrdSAuFD+ul71NCoc5e+dgBOwCA4Dm1+E71lzoOOW
Gj0RQBOVRxdbJHDmU2L0Ikq6olsYi/sAYygQ5iq9cgEIDDg6uNlLmwT8Q3RBT8yP
4auwJQTAPTFuZB0YDJrhYP19pWTz91t44CCwHSTs5X9EOaQmzPHEUWI9aW85OFd6
mD8DJWG3sjpi7H7VlKB7Wr80vG/z8boTesIf10ehObQeREg0/EV7RiMggaFQWEn3
v4SFaw+IoETCj56nNBbJAdHArUVTxvfHRZnVnp4UuTjBtO6NPONWWe0eYVh1PGkP
EWqN1qns6sHPi3NDmCGFNjLuJPviHpByRdDTiw471icEAblxYDjebRQJ9moFwQeR
azaKMpSKUXGwShzXckYTKc08rP3X4qUYklmQuTNk4U+N6NqDS1cWEiYzAkWXQrQ8
UN5mJ2Vr3Hilw/IJ+8+VnoM5atvYWCjACQ1JsrJnaul4rb2Ejwt2DdM1ccEzy5Zh
m6uFGuzJ5jfm9Rg6DEZRcNu5Q2a3LaeyiGSK/DIXFv3icyukGG5hJPoVJw19M9RW
1CMTmstHa6JZegGdVVYwclGc0JMZm8cpHAG1iq7J+mi2LgrDgrSEPNnbfLh+po1h
Oy2Pcf/JBKpg72mahgcgd4c7YIu9c3Yum6yLHyt3TOYKM5GFxBdN9zo/8NW8nNaW
BI3k2gYkISd9tpDtJJGII7l7qinOe+7hMF+xZJeH1QJtOR26WeC8x7YkgIpbEvbJ
hEfOalZHenxFMNC6AVAIYISyillZo+9FYsvI56sVTd9WxRuwD/vfQBB7Z0TUYZux
vHnSohUrSF6yH0he5rwaMZHnbKXzF+LJj4hSVoryWDZPcfZh5Z2ahXpwDTR1sQ7g
Ioauj4OHjMcT24G9iHp6sWX0M4sXZK+c4YDs8zt+CKaenitPLGNmqW1AoW6M59kr
18jvCDV3MiKlf8HdEV42F7MqtIa6AZA4nu/co3IDmJi97qOLJQ5VnJN/JUAw5fFa
5VLfw9DBFr/y2p3HnAZb4Vqa+0PjMFxSbBMpjJ/xCMGDqe23h85jcxbtUMgseZSc
Rl3shqM4FFTE/UasEqlIakymMWmFYomyIhxCJuW8uf15lU9Naa368d8Dyp1CQFcY
ian2G1rCjn68keLW6yaEANhPpAjTFjgPchTYIOlk+CJySk2/jB12UQQptbFvQeQI
T45+mH+KOhlv1gMJGewEazkiAldYP99wlMk3AfGr03qrGB3IothjVchWBIljRCnA
vwcTe/2gz4P0wvPA0rhwCFQND1+0H1HKiLMRNZXSOEX6CD0OnDZi1lrpa8lntBcr
Pah5GkX1yeUSeGg45SV5SJ3z4O7CoUAymcJCd5avLci3dof4N8QWqzIJRkYFv+YV
3xpE42jW/kyXb0m+yImj4i23iby4jOei3GJ+Inj+bC4EP9BbIpaydi0THVixC0w0
XQotNDlSWXXgfw7nbklWYLbEeb4B8jLnMSkEPvl86lJQQks146irCGmnOk2lHV3K
RNQdb0Qv7meR8n64fCE4h4/7E1hl8psH32akiSPdZqKKts7NQFNanV5xdYnGFgQN
PHpcMr69rmKoFwcU9CT4O0LCl/l+AMYLqeuyK/F3S1vOKbgKf4KFrwRSlx/9vcF5
J/YbJQOILNVaBLsXPR5EOJSSU0bHjA4Up10cGZyxgmlSfvp5kqMRYOChIcu1rRnw
0Aqtk4jtNwIXhsRuEgO+m2ya9Ip+qV9ITRG6FJ6Nvh8l37HJBCnu7Vz1JG7gJejC
a8WzRGKuiwdIAI0cTHCnuvqqxp1PE6G4pFCHd9UMU8rZJ/v1AWnSjAY5zo7mByqS
jNX563rLDahTsgaZcA0HGfZXJAucmjCnlBgoZuhlMSkko7ES+LCLGnomP4onEiB7
ycOGye12xhXfOuUc7txXFkt8EyTm7oTz9/+MFXz3rZFbO+FCFNDIKVDSxvn3pqJO
CymzybcV0COxQ3djdn1u2e/RqPO18cPB8jon348VnvoPUwNYAz93F/ToZtF7ziNg
JR3e6po8zk4Uent16UeC+EkBxPoLabIvNkfCioWXYfcDVIDHOtg8XaZyJuZGEyKV
5q/qG8DWkKPwHoaduxqxkU3jZ5zwBJQzCCtlVtEuKYbF2OTZ27/9N7RBbpbpAKLw
vcSJ0gKoFTJcmvSFTsV+TaPic1hneThHGqwpXl2BAAJxKXNZWYD5lKeeRiRXU0AQ
WhpwWA2fshyzdWS5K/PMlM9+xYGb04MXnGodJ4JWOLbFEooT9pumo11UJ7rF+cM+
2lNVUMO62zVPd44ALrG3X7YM3pP0Qpb64Fn/c3svM1ePmu0nGJ1bGG58Lm78A4F4
Ma58oJ9Vne65Q+sZOO3pSoVRLOPTs/akBjHF4b/OkkDpum2hJbHiXTTXj5pCwapd
dL499smF/RK1yUyDGwAlVJARcssMwHyDkVTuvVzjQxAPFVVdD+CKj8kdqiONnUQY
OoPQYRdl18pdik7n3bVq/d9QJg4NpE6o16DZrN/ZRscMMmYHpCrG9GjywLKaAPBw
D4pnWlPoEJO3gAJ02WqItFQQ2GYNH2lmWMmQkp8DTbQ2eE4504u9zXoeopArZTVe
rfUtWVfRs1MY86GW3mx9fYX8WaIOBN3eqyYYgv89KySqqszKZl4S1sPQtv8YLFR2
+XRVXtwvQ5g8uuddGbfEWkA1XPx5zP0pKjhvyCWNvzzUpVUdyIjhz4wtneFFTWV2
W9AWzKdCuNcFAaYD3PvsZbgPaC0jcd2Ins962wpVnmZ/aX4qQEXrmPte9LGwmm70
4nKK7VYgiQS9UuuctR1agSmRSnbnai6apXkiPady+zWZq1+EteuV+R2CNIcudnc9
x3alGx5XVDInznqqlRD+tq1R8LRiaOenAHVuyTpZpTdgENhpXN+ufWwWYPfoyddZ
Sdk6u0rdIRFEabwsfxNpf41sEIM0gbRXac6mMHQk8lGsD2J4euNj7PdqLOYuXx1a
rBmbj2Z9CRMWiz/k2jHEj0NyaHbri2nMXrMSjBd7rYDNXWUI4LbDy8H5YfUGflHH
1NbBrM9UQsRFK3EVDR+P9XBq5kstmd2+Fm9d7ujd32N0BIa+YetRfAc1AwLkwuNV
CgYZIOdg+YZHNUwUSW5df3nsIBQ0ohEBDpCdw+U5g5MrD5QgyXQBjYSb+AJAdfd+
HqqIbFGQeRTEiqrbiZuVUG8ClNVoGlNp9b0zu2Cw2r+cUf9uq2Bvi/QxZF61IPpP
wQxHIX7iYgRtxqdhOXgDC6QgaS0/NstZeBFCqIGRRKSXAQOqzffadrYKTb0sgiF9
RFwJGSZ57ujLIXt9GB3gNop0qZ2jG+Z6+W/LyYZ+hHTFCwlQ+R6nJb4fAlIVdc22
93WybIT4fPX+VIIKRf8wq+YVLnTqlzWqL0V3TQxd4DlFY/QSPmQiUn9QGxtuzIZy
nblkDWmldnLLYzRtsPROq9x3yjnBiFBsvmvXLzNOsDQ42nBwH7xSeKj4szGqTgGT
wxU+scDJo96tVBGiyHh2+TIW9gCTaPch+D1jje9rFpPGL+58yF58AGtD0pWqaqLE
rmv7Sglv5VmV8DPH8YcgUr7VMsrLgXi00IXIgk4mreTc0c5NhMO8F1h+kYp+DZEJ
3fq19r1jmjNZhc96qho0BXtWKLkJU39VkDK/xVmJBK8T9H1jYnwiUtSMBvR39/0b
BEb572RcfS0hZMWLNwU6U9eVY6nZzyLld4uGV/6QPYWUWHZq78+enEqObuiFYk2m
YRlWRuuAgsAPXFI8zeN6ceRtPNp8wM09S0e9D4b7yY3dJr2eGr159dXgJmhvCCWP
mywrvPIFUsT6BGcua7rICx/fULpYVAhND8knZhmXPmw9klkxxtrSd/zXppKeRnOv
hcUOQSOqB1t40ZkkXQOvic3RPfxJql28y3Drr0zOEIgdnpUKMbetQVACu6wYG66o
jEu8Z4A8Q/YdFZJzn9YPXHmUUHK0OrvCQH4TaeYxoE0O6GXNPVcKl7zayKFnRbWt
YyXKuwILZI99oK7QH3bjV1gii/hYPvWLmYtGGc9z7Bqb3SATHnUJuC2Uv+Vd/65J
5qAIJUDfmPbU4Q5kVL8TKvDnqbw+F/te9FFfUv61M3lthS0wczRcUBllTVRZ9L8u
t+1189zA1rDkSdE2ivA53HyXee5gMSnJuyS+7kQFcjNy1Om691PG6YQ/xZW04LWd
bP0YRPEnwcf2ErX985oP+xDPhBggu8R6Zgo7buH0huC/7VoUB9l3onTR0XW8ScIc
q75VmKRsf2ZDTjqSwUNrEGFGq+WDSFxqZACIIa8P1HpjnAlWWinkb2/HS10CYJ6L
hfiQn4GK60p+uh+wop/fmEOfjSJRzAB1IWwc8Fkk4GqmvzTfRYjSse7GxBkdNMhi
JvrJkhIb+6Rsm37jCSqAXT36/H0OnyIw3YLB0FR5pa7ACcW6ZEgZXpXFzpJsWbWl
bAR0P0/TKyuurQXcA2QVv3PRtE3OVShOfDD7jnp4iDZv6A/17I6D7F6OQ/aCuYsp
LoP/g0YdnsypSiTgqQCIHNHFtMDA1oaFrNxYlalvqka8QpRHI/RbdgLbOgjoPK4q
rdZNig9/EfDPosguUJOR1vcno5N2QdYhjfZQbuLN1bcJLEX0P4ZIjW66M+sxUh9s
5JtfEUt1Wg/wX28PctvZ6L0ZGTuvOhYVcjOrVKb0tQz3ltvGMRwEH8FWngPkBPcR
QIY6FvbPG4TOFDuWnT2NSnBLBWpBkodM4dfxgZ63wiZ7tyONNiBJ85AKkg5+tIjE
UGpweFHNk5ipP8jWkqsZx79V6pcYecE7/PJCiISL8L2fJsq1mWEsLrGMAOViSxZ7
0o+M0IcTjMxE/HPBzk9CNTpEH5sarADNLHD8XpfDm8yffB1VDBSMy7E0NPXfS8dH
umjAnN3pL0nKABfUo+t8W7vSsn8L5pNJh+/nOr/MlnABozTBq+5Hx2yHXwy4kVA+
mPUYxiVilIWloPaeEbBBn6kZFEYOOqYECUEPVjlIYumTxPS9bahLuUclW8vCAVgm
24yUZ46Z6waQd0uHNQS1qRZTNFIVnzKs+JZOfILtP4IkVuSk+homnuwVGgi4im4t
ovQvME9u3npKg5JBCWzta3WtmEFHntQNJvVQ2litjEA7SG+FIp2nYkgp2BYc4tmA
b+PFrgO6sGkPwUv2RTexfSwFueIze1tuNCtJFxtFHq+cgUmVlj3GigzQJ1Aoe8nZ
icWGDNZr7wLMR8SS5bat5hpVPjfkAlYZgykVd1EvLORpPkTkuIJJRdnCgNmEDc82
KiCUDMZ+LzA402bJcYyc1UxgZXGeAXFrBlWVqFlqj8AWUn9FozE2UbDfadt6rt9Y
O1s/qJyOU+ptGjy82MMdBbErGl124RKE0PwxU4on1K2IEyF3+2vLvKWZfSJIupsC
1saej7+XBSxTw0wKcRGVeV+LdpLhLolhTv11GII3I7Q73u60Uf8pzoHKVUosG77C
tSTcPWrTrn8kEShDjtaDvev2JtngcAXG/Hv/B2eWvEZ67q9aksPnR++9C++XqQ/n
0fJYs+gg0dyh8TRYF1w7M9oH19ug5AljdcF+VS9vBvc2fyAdENabmeA790g5bZVG
YpgnC7x0gOF3NXmSUmT/3W6os5379IquNV+mN6EkxJ9d42I5NR3g9opq1vhCRk/g
DXqyeia4Q2YibRxkDtkOdqLL5DygfY3edst9IRE7Zs4vNM2By4LK7FipD+Tir3AS
6+PEl86IMfjzFDjZC5gN5rFtBztWB2K6lwQxa5Byg5v1BXbCZqqsPBNzCDFqwMuC
BongpQxYFfnRUfPLqvpaEvlMLi3vLKgxEU+LbbYiGOBJ55gqGLtqtNJ3sbgfSCsM
ybZ+3n0kbVkPJkLhtRx9bBH7l0OQ316/yItidq+ixqT0ehGe+9kw580CU9OG4j8Y
sSma4SFLF5qAi84F7V9FmLhyaLweFGf51H3jAKL3PGHOy28Ru7siOicof2AIfJBR
ymY3KCKEMKjO1WkdoFfIn6D2aHKqDcco/P7KwzUpPVo4uYM0smVh7yfUvvLE1Pp7
0Xz3SwQB2/WPtDfw/nd1B6lc481yLrFT4wUe6Sqd4RzT1KEWvs6FDl6J975hdGxM
a3Ob3IMKttasfVfNSY7Na9L4dEUk/8ECmZ5dWSYd8H5qz3nz21Wc45wwXz5TjAlH
VkXa0Km+fuADaesciFPAPYEjW1D4GINo+cfSOoX2Tywx0cprmI/ZJsCtdQ6AioXr
BpwlhT+oc7f9q8JhaGuUNEL8+mNxSDxVru7PhNkcTMobjbm5wIwYLElIsxXIWvBf
2xhvV3e18SbXR/E+ohYsFrsABmnDwICxjluUWSW+DQIIxOsmY8V5lYCVL9rsUAiw
Eq1WDEyn2pptT8huqUcfuA6C30Yjn6DHYCHe+DjKUl2VrJJX9L0e0kqa/hWxhLUP
3i3fWqt8pZdpP6kSuET7m1Kg+CE80QVFnrbygkrNHqzvtNR1UziiRZfx7kIAb1Zc
WwlvLdG3Gb6+qEIVPttyIr5RNVcY2CYqZOE5o97gX8/gEICSxbFee1xZ0XQg374y
BIpNVnlQA2J4ieFZG9fDVZlSUV3mKuJ4VO3AjCPqdq23qhlXgTfxdfnIf7zWLMyN
urfU1NtnBwntsqtY4yfWDSMZ/tND2bVFVhrZXil+LG9Cqrwrm4yPjzqgd7K/6cMl
v/NlgxIu+p48AkHzuSVtE124fOrIf1qFLimVEXs1xSYir9ibyKE9ggPZKVTjKE3o
UGM6GekzAFWf73Jj9uRCaVnkUlKWWqNakNm1eAlCykAmDYO9nDWrxBJGC13+vBAB
jjYmXVD0jDpL7aSt/C+WM2imiGT5FA6VIgApW0nWxDsRlW0Bh+NKsPXAbBPKTWxF
exBBC8A/ufRDFyZWjhF/yzY/TOKXrCnWtKFlMnofaZQoZsp9qfUoHHn5sQWcumN5
EW9W6KT34b4DUSOsmb1cXiHuSa4ZfQ7GCM8HUNzZzPEHZOUad7bIMvUMs2/Hp0dF
Z3IcP2lIxgWCzCgOYViwLh7pVhpg7lEMawXlwv9DXqfOLA8qF6KI7/X3xKCzLUcL
G266wEsKiCpygN+xsq8fTA9ITHRTkRv+LjnYa012DFX0teTVJA8t6TjuaFqbl20k
kPaLfk4STRliO+nF8uyLbRLG9MG6PiujM7fONokmgEZrNeXi8eM3sLR2p2cbbST9
Ojd+pvQLhh7UJYdFntrrDzSU8Y5XhyWtUnLewaZMDI8GrOjCmhSEtNWEuSFQgdfb
xPq+/ByGmZGyt/lIanji3wk/DujSz5d8fX2NvcKxuG7Fe1oBcDpUqJRExnoxQG+5
SGODoS7su0gBbrRN6Gm7Cuz3lR3/jBgHb0PZkfRO5AcGAmdoqHG6FDCTCvO0m93g
wy3I1pW6DDm+doGk/VfkxOzRLWBZ/pBtiijmg7+7Ch8ellEUOD8MRiWRp5qOvZfK
Oq+I5JgaZhSUO9b51EgiAG+gdILfpZ2Zl/cePDCvyr08Od41MeRQg2L48RNdmXqs
rGDbrUg1CLhpLrCM6bsuZqi4pXapvRi7mKjN1Uo1O/YOOQjYjvpuRUcoOgfi0Kqk
nORxf8IQU083Hau5iTe7hG6158z3sqQxnD8GW5Exig02E5R493V0wOeAem9vpQJ2
AskjRHf71k7OXjAAEzlKoc4tOrtci8bgmsjWUAvJOzxwfvcEfT9j7xrqhuSuXG67
BEs72ENNwVjHRZMiibicBKpe0mrXdE3LLJkQZkolMpphPjD+nGpqgIf9NE1NCfR3
4R05PTnjSkfNkOxvWtkYpRpu8TrtQoHzzYvI7NFT63Q/OrO4wPfyAn8FHFFCRhHS
B+Lpp4Q9/0OB1u/uepX1QwML/SJOQZnQj5RjY3Gfi0HK0Tk7iqJYUz3PTrrZJ0qO
ozhOr64S2q/z7LrQutftLxvKAmM/zUzfgjd1GvsLyTxBLqVVVVfVmz66yfZlMsCY
wbsZgLI9PPNT/9tERSG8R7AB9DSwK6RcbSo26MQQWOi/RtUu8/HcatX046Rnr51v
vN71s+k72i7ZnxfU6kcH4awjKlz7Glr2Ql1ZLLxslGzKaqW2VfTxg0uFJ7gprfRb
98mgIHNPAfNVU6pjmwBuT4B9s+2OM7X+GyFS3ZKhtNyHPUxoO+VGugwETNn7rDhq
2mI5FT7t0kXRGbwrApWIRo3VVQE5AubGT1bJzCznsG8UvDj+wjyAp0ufGXjC2AeQ
OWmwo5mjRR6SzHpRBcyLmHAIPotVRrywy74+CDw6gzcjF6jugnMQUMT5pqjClaER
aK1ZuQOWJAnKJbSExWsg1CnpJuD2RBW5c4geU7qOddoBkLzHKdvXq2cfZ8R7berM
pUdR0KEonWEwizopyQjUq4cxXw9XRHxZgINWwQBVM6jqmGRDCedR1Xf2fwAzOagu
kSTEJiC31dS0b+V5JWJ/bgdaCL2au/VrrUqYs9wMe9ML5rjlK8gzCYOSH7IXCu48
BG77n7eTMprAp2FZUalf+yRJPv47ScxBIZehYnteInN6pYV1nfc77/PxsgVHKmAH
W7Dsf3oD0vQAmb7LEpUJW6owyWOkS/q2nSEHBrMsFPq6XNe8xHQBOemrLSVaf26g
UInJJzMABvVAddSZ8NtaVhZN1W0d/6XU9XeQMH8jLugINP+bPh5fgmdoFKlRsrbW
nb0Nyyhnr4/PmeJWxCbTqRgLioOAgfB1Vl2doAp9wQ80jI1CsVfUT4mdRRqoVZ3M
64qR405fETpgR5KKOazMrVPvUhytaH4AtdPBzQq0IKv5Hhs4z/18Zdy1xQhipmkw
pouWkhp3yqET/1JfnAnWOPKJYPGizjkqLa98OZnswaGyNXyABvQLvHXXC8kVYfap
yk+jOShXhK0958S5qblvXBjav1GajVrIMb5/+Bwy6oR5d5HZH2eURkS+ajraJzsX
JVRqDIA6d7qy1xdd51dqe+TZaC1oZ61cZ2ityojR9vg56RhjvTMkVTrSiaUjgb/d
fm9dVj5rtwExCl+iWyX19oa7UKMC3mpBdYKvv3D0Fhh8V4BTAdJ3tViG3G5AkZ+x
Jj62N4agIGa/gZ/Bz4Bi4Luu9BafIyeHo5dHyL30HMB/4qzxKedeYHBDydsGVBiC
hqG+o68iLMbIvcmiQa2WhsYDneFXoxhucem64oHE508IY3gXA9lVBzmyUxxOyrGk
4Hvd2TcB+zXrypueJybGGlQj0056O4k4pw3/EtEPSSHXtZDqYFEDVFeAsnsiGoMf
VwvPSQlL9PgdUqbQQgPe7lbHizWziqWY32Z7RdAThC+USdnUgsjENp3xlzaAdlfe
dVavlMqGZXBG6Op8L5PtNqmFT7+859ietIwmOAd6Qw9CFND2aLIKIZ8al5UPf2sF
9mFlR3evOzgt0W5jhC2/McLxn53fb0AsHo5BUS2NwZXgaitn7BI4gOyxo/19OoIz
7+y/0K0eeYv5bXhJaNoQKC01h8miLlCchAkzw0Nyv70tUy25n9AQFbN2qcmlXxbF
JrYKEeaBZdv4RZ7SpvytNK0jy4oBLuQFMWTS2aKPyMmG2vxqDU1asjSeIk1625ei
OqhLG/H00d/QLrVtVSy3p4++SWjdF8SPldxyH5sFqIxlaUfYK5jj8m0eosBOas1A
vXbA3RvVHvCXL4fW8O/EWgSs7Lc7AYebkSTNxTU+Vba3Piz+n8Z4DiDhUAVs/Y3U
P5q1iuZhR8iQPU8cySs3aOEVAJZVK0NQAyHFNq8m8EuLnmb/dtST1iBIzJXFZ5aM
AkxOJLlmQML0EekmfCT3E8zoW4THaF3u0dNQnvUZB/RmAkIf5T30g9SnHshi8UYd
7Qlfm1chUdQ00j9RO8jYftURtZYw+TPN/IVyzDFysH3SRLDzOB6TpJyDYPgIOYXX
xLOQDNbUrybxtw5iyrz0NoWWXaxKhp/rkv77v7j4ClofjUJPDLbp8yr1kjb3RTq5
mZoukSm9ldatmgHybO5msog18EzZ6gNevKmUynRvMA1F+R6U/Q7iBSICecYnitW2
k+KnCKE+Vg/jcdXe6V7ciqU+VH1zzoCmC0GYyCY+L3TsDCO4GhtG8tvtpsGw9xLO
/1S3Wac5ITIGpiVMvaqtIFrUX86HUGl7vkLtIqa/7GF1lWQzpnky9838I7LsAhvm
rNF0/0q+BTeAnn+M0BaPiw0sMj5n2Ug7wBCBCN9GcvsuOMgUcmH6mYu7JA3Oe7OD
iQhvgVTcXvYnbYlEOYjgdOzllbv+1E52/Sp3ZKZLtkYdrP4qE5U8GZbzYF7onuMc
WDcZBrZUL9ZYRfTIAZL+N/RRcRmtwxSnCh5hPMW4PAU16tlVF2YiTOa5xCCwrZ+S
StraGAoSk+p+fuG3t+/vcGG8flBpUT9e8yBPzS9oCFkEDXr4Mf5sCeSrPQUaCqDT
/pqLrtxDKez/jxbUtUbmDkET5xi5cYpNYRmU6GQyBnmC8nUfltgVz7TAIRD1q/2x
bIztpCN5vrzMxFRVh6eCWU4lJI0yF2iLEZPCNZC8aamSBb9q+nt3EAskBwcSWkbh
sSsnmsXKO1H6maH/Tgu1pW8UhKuWABCZ+tdCEdkK9EhQvKzGDyrPl0olmaHh5Z8k
Xp3DTtNeE03ORD/OQ29Bs9Or7oonQWtt6cG2ZsMHY4R9JF+ChV8X8B4lVI8YeQws
iVPnOoEfAN4Kvb7g7DMqSa5+PlW5ipCnxMAanvjpGyHLdNhkwykyqMZY+kE8G/L2
/G4VNfng/m0V+I417cywLSQvmR489k5uaMDLnlHdseRZC0rRCAQLDbeBaJTawOPh
FLG7FLLqYWtTFkPgT70nUFRf+MnEhTCiYO3OOJc5SnW5vb2U2DCO6cn6evivtZ4S
cY2dyTVEKrh+xoM283d5r4iwxF3Gm6HhNFZY2JmDnEXuThCwi5xCkon/lMpqFktb
VghRVR3y2GVZraXUnNpBWmjEa0d7mYkrgIvG9diT+fKhfh8tu3wXilQGB94A8len
WHwvuNcODC+cR+lrRbqKvvKHT0PPG94sHzrVXhVBRvn9mKrdgcDhU1hBDZ7+Fhdy
2mi8QgpTX7chIxzF+J3xttlcB5RMHa3yOZ5BZaGNp0NLOY5Sb8UP4060PutXI9Ak
etMedXKKXBQZ5gBAmRUfVD149ypekYuEckNVUtWNaKGooRCiUEmAx+7Md8sNQLFT
PXa6qJKaFFKj+J6ZMZ2DJaHOiiUI/2xw6LhqIzpLQKihZ5hx11LVBfDfAc8mmz2x
5zAr7+7WU/44C66Ty3PGm9kV8cRMk4ZuAeL9yB358OD8k2nCgfXDivcND+EjHPvu
IgwD+mz9v8pxbtm4iOtB2bm8/D2rxarFOUzsgjiBDSenbzrObifPd51PD6+Qk5/t
yRJmRq6WFOfbB0dt3P7WP76kc3rXpg2EE7HvQna1EtVAvIAJeRkOlU9ZqfwzIxSc
/FShkzp7HTp8nXlujF379hP17mA0keEcqIEj9zBJh0DMJyaahTV2tNIxC/ypyOqh
3SzlMGnfyMp/2k9GS1Upxg2s4UIa80TjPmp6jlPgpD3/vInR5Po1VCwUWwGy5T2x
T19F8MuIL3FT6pWXlbCsbLIdCRcxSToji3axH9WN8BCkPQnuvITtTAKj/cJgrc0n
g/eYPO0YpT7obuCpg6gCq5kWrfPM9U3XszWAsxaZqaJjCgbvZebX2Y3MkxRFREam
/sgdUqhXQ0hm1Mww3VbcQBrRHvrQVLDH5P07FixRqSCd61w6FuE56RMZfiP8BZkE
b8EiYHZ5qiJQFA/EtMogYHaYun3I0hMZLu1ihjJBCyVAjQLKffNf3f3yGDhIcmhO
6WQ4eT6QQM3A3vSTW+bJ5kDOM6IwwrD8fgSQ7QpxhK4/LtXWLnp237uPkp7Ldch0
FQl2DbTxseNLD4nzcEkTbWaeiWRHwLFw5+zI8d0F0kZBZpvGoQpfW+VXGun+i7Fc
mG/VvYFUyy52SkyJRSSM06O1fIYreWyzgQDZt99z5o9wJn6HoEIO1Xqd96PwglGP
00/4xnLbWgQQJsXGmXfRvrvY+/k9bnjPejwWp6O6jfpQIWQhoMpzATjNwI3OqOLi
aPmQ4C4vjYzIjPakSvrr22jPRjfTNWezbIKZsoxBrPU35UdNFJg/QKZNl1hVwHRX
mXgJMY41Al6BTrI4s3tXCY1iQnRsnfaHsq8hlrtbAdU7D1lh21cYNiIfwVcldAZW
MvpoAaF//644nm7Og1LVkKP3X00EA9p7EJqA8ZwxP374v8N6TIIZ4hhbbwIFol7o
XNGB9rV7GQCaqLB575dDb+dCOfxE+uaUBduE3jA6afHSwxF9Y+h8VwfM3hEpI1+U
dQh1spQmtBQ/mRe88G5ws/z7J5FXpGEddq/w05uLhcLHOUnoFz/eLc/js7JeEpSx
bx4yNw0YcAZYZ2OWBHjjaskcUcwNCuDpBx+eQAbaeQ1F3Zk89xsV5NAvVvK+5Hv7
EOPbNbpjtyR2nl1embrb93A+w18fK9mByEXG3kua38u1HnOdt1Iux6gFdO8oN6Xt
ULdNk0H9ff2hfsZKx5R9tr6iZBcra/OPc0t3tGV6F5hvxCdYZxVZ9LN0EmtU6S/k
ZQ88lwU6fU4i9jjivVMgRd+J6vhBu5yLtBTp/SB6ggDi3CVTJeeBIWmPvql9MAKf
qI8San91Bv0WELlq9NXnkv1jmnUqXXOdHEWJ/vusZ0PUD6FP4v3xwV/AfFJejCa3
3GBHbscKj+JZwT3gQZO7PZnZ1p78vT0iKCAZZPdhPuhdaxx/SkcBY9Uqp0xlSF2R
ePltKX7Zx2sz4BInaVov7VdYLnlxED4ZhD83cYA6E8Xj/7KpqPknY5RQrjlUWEYv
fT7SA+fjKyrB3il0BLTplLJZwCNyQ8uSupcuYYTy9j6aEDyDG4f/mEWmm0uFll7A
gPQVs4zZmhJ2IeuBN8mrGTWu0LAoO2MjIAHZswRUj2G9LwArfqHEPk/M1+H8c155
k9cmcmIzvnhQx3wawP31WbvwVlkKksOF/nlGs8fulE3DS3rNVX8B8HPtJsKAdVX8
wNk4nFFGNvOnZqqaP3oPFwhyCvi/q53Jc4ldppcdCQ60YTHsy/ZuncBia0hGfdxP
VnPM6TwvRcC+7qI+GWL5QJ8WNutPsGVKdzQUVMAndZf5MkbZMsS6M2RDSw1Rpeio
fSgQwLbvKbLF0YjnYnBUlyA0XdhOc9Yk6L16cGyaxQb8XClxJBl/NuMKDrw4Tudf
lxAHsqYNG6hr3J4VZ2X2O99qk/oUy7Iig2UiP+PiNiT4NXVZ7Sm1Ib2nkRLi/MZi
lywNr9thQH4BtCEOWuAka7tddVUpzIsViybaCy8AUf2DI1/WEzbCoNANFAHHXa1y
nrVQmSPTSxZubphFqcWMT4zW3LMCjdJhJ2STMnnmW8rlURtdpNC+DOK2bssklmRk
4MUoMl360TLYIaw/gjB3Ev8Afcs5XedWKKbiJKQtFvQHH00nK1eVOCMfWc3SL9tA
WYwpELJcGKMkJwz9FLmW1IrmPT3dY5l96IbSGy4045or1TsTCxFCw1qAio7x25Ag
mrNX6S6C30otguwEPqMc4lhpG6S1Pgk2+8+otZt/H9EZUfAcCyWJP8kDg/G3dZ6+
vtMp5PV8iuumWU6tpnrIbCiWPx+ZPcNh3b5z/f8LPdQ4NQClmrQT9bMYuPW8RvPT
OUErU6mI2X2OfahYABlfdcvqp0XH7qTbj3nXmZwsthgB089cM+qA0sKiA6g3dHTA
Uni7fJyPaITQRu81h+q0m0SFX3IXvL/82zOHTZr1zLF90hiFRJ8CwGOxaqH15gyd
v+CvdO/uPpD3cD5tq9lPBjdEycxvxmLmDnVOuN2D19nr/dzAjutucoaupYF7d3xA
5aC8a5pXo+WCirF8woiojapaIhmdo4xFI2+7VbhE2Lf7jHVzk14T0zB3PSLMZqRw
gr0Mh2vAgXZ5A/93EzFfS7JadAasMrTn/uq4WHPmThClnVa/3ZzY4p7M70rXw0wI
3u+jpKJRZxEJGDZK7gULOdeVv7p6j6jvafyT4GUomrpRj90mLTaeSRLdHk+Mnbi7
oEkpQE2LL1ohaQO+gtWL0mYhhu8FtUc2dhwnnqlK3mGxnOUYFWrTmfqeFmYtKQzb
9MzGz2OEe5Vi5qvJIxMZtUimUr23UCuxoAq+87T/SHGmsP9I9ZlazXmUQRqY1EA5
uiEMGIqDZF7ea17kmdcP3Q6oYxCNAzaBVV3F1JcLC/HQ0XyXpVftNMQL3RMy+Z2q
2+5erdMyXBLmNK2wrGj2zj1YrOaqxmPbGNV/YwpGn9SulYcSWi6tcCynKLJhuLOi
MajBYvRG8mWxcDXxtpWMFL96uL/q9qPNtTMpy8Moyzq43fkDzuh534gJsnW8j2w1
758EXbN2owjpK3SVn+yCrGcPjEMEXA4OAiqpaf0KQ6EFIH1mozPRpupel3Ik44Zo
Ud1xBX+LR/Gno8LrFuTMQAnIucGvkMlok7+4+FHlv17j4bxAbOGmgmhK0fjFgK63
4QBXdyNiMpA4DZxAVgVKxyx6UtOi88FAjdKy2lk7uiOKqKtdeg4pDbZJossVok9g
7n3eNtlbw8ng882rwnlJMLLSx84DWesTzmzU71sHoDkdXIPs21IH6XdeyY5P0rOs
DavDvqZU0gy0LDThCJzn7htJvSYAcX6EjR5QNTxjWrhYo8wsG36OpgDqktqm96jK
uiONrOkvHscB9tZv9S9ES3AW1gnUjF47eo8dPg/ibDSZH4luuwgJoejz6j9j+Vi0
8nBXRQYDaLnYiUEBBXviY+jlQR99xvLJ6Vm7zRMsVYaDUKVa3Cn2SmN8uW1eT2Pz
wniK9A+xyYW7Nvdiwy3cY4BhaGWOhaZZC5/dKilcjS/OWSWMc9vzd0JaerVDwlwE
WjXXO/IGuo7qnXiwBKhkIM2uUvRcgGdF+80m1l+9QuMh6lF670hfHrkPm7aL+AH5
arQrpJ0z/ZeVdjjwhkiRWajJLZRQTy19haFUCAfXOlZlbTZoZFuEB9W2GIsfd6q+
mRpL/6eJm2KGEt4MMfFcZfHv5APRha1X1lHyEcXMGhK+xn+8VOingwA9lfWprxex
mo/0zl2I4hb/MsyOOyzDe8E6XV14Xd1IEfxaXaYwLYB/gdWPCVEyo9ijvebZG3uR
y4YgJzJZ9txBpWuhLQDPOqsxVwnaAMC86R3hrbpcrFPAbf5AZjmGSrB++UiSzAS5
h0UNs2LYFbOaBsICYScu7QntZt3l1u8UwAINu6ks4jqEZoSC0p81gyMqJ6MX67Lc
LTR8+DmjZ0TA/DQBqet/ryfwhfuY6jnJpbfchICHkibx0AT4CdsMDS5DgN+Axx6h
c4KZ5IgekgNS0dojtXUAF09HZg4NHBDhhBFQ/gn4Rj+nY1kOE3JP8ZKnG53Z23Vd
oBmahUMiGI+XGf8EdvpyABb6WbmHLwS8ukzAJhZ3kbcX1fryDy+QmheZ7leaDnSl
9d8Sj72vpSHfJb2FllQ00y/ILX6ohdQbkk49WR7jYOQcU5r9GcM1KJAtTCaMUG5I
o//ErM0soLm7yXdTSt9hUxn5jf7EnyMxBRGPMBLAAEagmlq/fx44WDCVTLIvaUMU
oPChfx3C0HAZCzNzTS9z3BG/Vrq5zq9OENT2KQyGcL5RGlPelcCeiCE0I/6J/gip
BMobOR0ag62FJzUUTy2/8rlJRJVwOk97on2WZXLXmA3umC1uq2S7cv8BT9RjntXI
pb/75Fk/A3NWnFp1k+DagB2jpLgZYYpl/b0WgDXom4dK5EeJLrcCyuFiHaWvKKAx
XUAhrLccqH5pyHzx1NG7qxYWAULPpXNiiY540Bmk3oQWU/ImT1DjdwCNu8LB0FKX
tDmqTRSK97YVyncjHtvtp+rDBpg7qYyKxhuAfPK8YKW89Cixg91SHeQlGVyBfFj0
BKBtXSS8l+zVZjYuD8PSUfc6k4+pXzuCRlfu3p+ucZ9GZYUN0hCN/8Ss8GVaYrv0
k+txorf986iD1/n7oij7VgIMj/epaAArRIM+FcfW5mFlq8PcO2H9WToZxK6lp/OL
hGBNnOGwlxVMq1DViTGbVswZ31IXGqODuheXQnN/NmmhT6aJ93il556SVK0tzaEM
xECWomZ6+pl1djgGxE9+lxE7eAkqsblAjOteaZZ/6qSGHFt2p1niLrrlPCG0lO++
w/7JLKF3jT2uPicHZo3vhLJP4gBJXJK8V/I7pt02gVUgYvxzZ/zh1wbc2YBweBht
F53+Qg3szDN1I3qxa1pd/0tAkNmKKR5B6GSETKWgWhR2nVo7IEJwqsxUCcCCec6U
6QS0CFs9J0isedZTI7vEhpOMRTMttvkmRe6Hg5XPrgejJnOQPiSHtfKS2Dc/U5l2
rsxSAAw4RywD30R8sW+uWeRtuaKS9hS5fSf5UPWK1o31403nMybk96ypb1iaStV2
Bjc0OYkgNQE66iXgrZqEVWnP3DT28mJIstXKCs8/xLZ4sutlyXS/C7n4BO5noZt/
ds18oaHwvav5D7rPYctQCmnQyZn1KA41uVG6wUGN8yF3pKsS1oXFs5jfpLM/ylET
PeWGAZHFQl670Lj2jDZKtE+EotRf8ZAMsZGIZuMwzqeBSWcb4YrYvYYfIiTn9Ioo
ElIBsTeUrgm0JMTeOLQhC0Eb0ybV0HuEdOkDUhAUfMk3JKY7EcpCHPncaGSBhJpj
w1HasuaWsjEHqr5ExYvCpz2wv6Oc1ZhUGx7QpjKHp47DkZEazJ7gCHcBYIAMFwca
KuEzBmsiwPyw42BipylCTgo3IXLHm9IkB8jOaLsjYfxi7FyT8vMbRRdoPdzyB2bI
utXv/F3mj9siMfJ7UxYkil3anhqhtY7kwT0TPnIV+IthIraF1DUsvhIWHVPHkYQi
NJnI0biZ+eoHvUoJ/ylyE4egX16naU5T9whyjIOJZqxvi15MxuYJ+rRE67H9HaEt
xWQSm1+gU0Ex5xGssRyduCSZ9ZPnQbEyL8lEkRIC1MZlkAurwH/e6BT8E/SPIPDj
Tc1cX9R0lt3pMWAATVpRicnqZmaE5RG/0RuPEE/53GIaf7Ky8B3JpPabqYuiTxlg
2gJgYp74Ldlbalx0L7LSOtVRTGAw4UL6dtHBd9EFFgKX3tST4p+SK0wK4ntpTSZR
rE/7YU68sTRIjFKxn5ovJPsp+eJYOtSz/MFACsw+rPaWjV86258vcgNcjALX5lfX
OCjBlUMmOU25uFEc3jWjb8w6cEELVT8JY6V7YqshTXLo6RShsMmy60LoegEJVnHx
xxWk4HcKJI6s3Oh6X9C4zfft1WLHYoSZZbVRz+kScmL5mr2yp0g+DLcYWOTdxRld
AqGL/LUya8M1eZ5tH0+/3JegQtsB2qVXfEQeIIFiSpSz3X6C9oI5v1/s7gN7+Ro6
Wc55dN0Nh2fdLUBmNNmXhthv5gTY3nlAeXWWthvaLo/BViPDnkq1J12mpm2CuxX/
wJwR8uyMalwA4yqTr70YoIN3HJjvZqPu0gT4CqwtFxN1eg/m7SQfXNKJaDdfnM2i
LQluj7k08X5vnbDhkXAk7vtNn/S8iKuS08YtWAqJIYpnpR8Lk88U5H5NIxEhgrnh
64ZG6lcAen6Ueo79xWsNiHTcxVSFzF86mVTSKAizbOHTdGpG3D+RthR6JZJsl/RR
zLSTSSfbT0rWwzt3aTjV5GRPWYA9i5yOHw597yY89vl4jd2wUYiyCEzhxOUWRMJT
GLCPvBGFMarkixA0vTPhQ9s8YCTsmr3qDjm0TqiHisYM33RGt6gRAHPouIlfEcYj
O4gemp7JPiYA2otfHuvzQeLFPNsxWAcrAQx0H63dDn4S23PYnA+GlUF0GECdag3E
zcWLzFqAFraJOXKIDKnCWTqDfYpOKjLoljbx8iAAYdzXxZ0G+4RY6WuFwEdLyunA
0hENzt+3uyb8AmlaGK2Y48pCNSqHFM/0FMhVMYRXpuKdwNNAfdShqWgSa4SVEkig
hkNMccPaI/XKS3JzFrlgntuZIH1fwcv5ZGyvx7ASmPuVd7S45B16ynSbu/OztXgW
EUxN3C/NHewqI/loRi52cY/MmTueWIOpyAFOlIzX3zSbP+gsCJtkY86Pm+6xSBiT
B9OvgnK4q+k+2jKzo8XpmXp0ESXY6ZLEzETdzIj3G4ZK3TVIUtjQ9YP/QVGaEnZK
ITZ51u6iEyeMr+0MaJ68jEwzyQ6uv5qmqozGAbNXrsGsn8cbU3AD1Ke8ljpRI+ov
sTdMJyznVqYB/tCt4ttMThNG93UwZTy0LDCNVJ68ajYJ6nHy/8FdI1Bg2rJflk8+
HWwvgbN5PJobdqG/h6WG9G0m7gdYlMphbi7tubPvJ0paPVkBNJFlM7zsQjuGbRI7
eH9wEMRjXOV7esguv82OmDp5Qx5JvnbJsJMf6EWsRnLppNp10JuU6n8nyYqilSE2
KLOmXyJhNeXJqedqfpHroTnpKadCRU/Z7NBDXQaZAnfoqnSHsadju1aDMYvVdXru
WqfsP+AYxuRoaGQQnqOY0NkO1x6dr1FQLwaCmpl8WK81E5A//S6HYIhcAVWygnG4
Rb0czB3AWjFeMrYeP+3KqCT6Gs52pw4yl1DJkR9UzrUO0CeJ08IZvc3iUmrkzjLk
tYyqRW854QdREHSK7h2AcDvXV66YKnCS7vYvyihbhFnJgYpW2kIxxdNUxtfWgrzO
Ss0nOCIlZoShwQ3uzd1S990cAc7p1/jM/oMWZes4xgexPdcTdHwsf8Rr7BZU/ih2
x+GqF5uuCAXJpsLz7FE1MaSn8ew9yh369qSByvdR5XaLEvDqEiV76BF7SqxlITD7
7Km6iZmQZo0aa+e/SVZFFLvaZoYJ2KPvsWsVlUJAUZNyg8WJmZddC9JA/G5ECoCP
HAPUyu2qY3NsOuDMJXVyNLpS537q2Bl5KnSjWhso2ELipAWEkepb6lg+VIzf4dMy
lziZIrdUn9ek3RMAlsDdbUHdDvoH3SaN+PAcZzH2/PG5HizfgbV5OW/yKaszlU43
RkG02v6TjlqvUyyCK46OLsIBMNd4QvYDpeSrBA1xVYJAv73t/DOTERKym7Ec0gZv
2OLkCJL7juiZ4ok+1q5nTBx20kpx7mys5DdY37PQUnnfHthYqzzdcvXc3VIZxdiX
t4mRtVbHVXGdKZHkmUk55pvjF5tiq9zpZOmFB4rNT9An2EQs/Qo4D/+Mit0NsOeV
39d68XD4ulKACD7KfmoX+aoG9sHRCzS1xduYwtavozBr6q/18DnUQpTmctE8llWQ
7/bPzhZUtAXOqNQLM+uvXWgQHUjkMWZ0nceh6czK/N2SAOkyNs0AgGVvDTRc2TSv
VuSzwK3TCZZZxxD+BKBRzjy1XzGizEL7kJpOPnyDJ2LP4+OBjDg1pm9uEqakssin
j8z//VaOYELmbRxkdkVEwkzgTTUAoBlYfplAb5DikDSE3D/OkXF+FHCIidgW0Pd7
OguGc+VVAeuF/rrhgGAE7elrzdCfwCCjoQg5MjfPeM8x9eVe6fe0HF3aYGWWMD65
0OYaq90NEtIheA3dysRJS2hiQJ5b+RfFicsM/uPZRiS2OU6p5sCaogZVsLnWb5ZQ
jT9SIGYc2NYuM31shrAmyLulEtoEnOjP0/eqPuSGqrP7VpBGOANt5MI4h8BKTWuX
LMl4Yi0gupXmh3fwK4V71YE1UaUePwhCxmt3LcVmlLNsHqNOfAz6UVS8BmmAEVak
lWcCsZq9cPHXGCo3T0He+3dEA15Vixf0iNtuGVXxSNJFAffdW0sBQpuv2+epekXZ
pAc7uvoWWZUhyWSuBJGAK3L9io5Cw8WuALbSH04xaNj289rtvSe56NV950wDO/gc
P4/NhxknmEHbr/CEVo+cOpdZeOOF4dLXhpZXjVCUrmgzRqRgVB8lmmjbpzc7CSzl
uXDWKR2IC+s2GgUvCIM3VUFb0pJMx4w7f6qAJ0jVvbXyZ/3lel1xrZlcrYbQELVn
wOlVwKWKQ5G9+qtoE/cD+/ggRsYXBEbBe3YXaGBLgLgI5jYUNjnU+pMBJAe7bNVc
zk7VPoxwzKyDm5z3RLZH8UkJdWM3dds0ZN4DlGtSPVCyvPMhoPCOqdyC5l4/0bEp
36ySjv/WzN1nU796N8aCsSejOQzsOneDzWMUCEmYhaUEzE37NTOR8fPvGBzOAqR8
hxhYG+a3aUbsmiAMveKSYTJx/LJXO5O3d7bk1NmNNyYaHC8GGdpB18AXHhXgc1UI
ZlJVj0y8yIFIgIHFi8xK2vrwnaGUl5p3WNqKAE7R97oKrxRFjvUkqoAmhdeVSt0U
rEC0y61Ibma43G6ajMsQk3CX+FzCiAOgp78XQs3KqcfaD1l0kUkfxc+N7rzEOtZe
HxrFo35rFY0eD+KXk738HvANAMvIS7roU+H2JCy887APuqyoWqwmtfWdkmFumANv
SmO2/7jfbgI8pNxM7m9ljHQ/l0BoeiMPSv1F/FZX3BwAXg6ummi+ZvQMTar+bgOJ
gprkETgfxBhp6t3EKmJ97Q09BbdQ6R0nnK35upHpv9TMUM/CK/zAnE2A91r/ph8j
yRVnSAXSgBAGqQSGsb/F+QOkVzc5dMHdsd0K7h3EHWstRZl3Kr0vpjitWzlJSvlq
3GPDGNUsxqSe1YUL2OUqeCbj98JzNW7wVBPxJ7CKmXF65oXtOAHPS0uMyaEgNgp/
poj6AEc4vctUbt3ddwd4NilxIucyqx3C7GXWHNdglUJ3khNXfhE2Z3mTra0/SQvB
a4IfWGhvZdLJQT3jeXhf8Pr2CSmQcVcHw6VX8mYLgyH4q69sjZDfYNxItOHKEgJ8
11oum7i+fHpjPpfFZ83zMtZPvowKcnOQGSVucS+0PtLCQkYPHtLIIRjPQ+++lwIK
PbSkWa5x4NWhVWBzbp6GfwYvF/Z5JOF3tv5UcmqBH/eACM7HMTpT/wtgbNa5U58j
6773GDTmJfH3JAHE4/GJIV3tNbXPu4y26mMessXmrWjA8vVXgN4UNyj7nla+lFgl
350zxepK0DPZyQfyCXytAWWSUq5UTCrAro5O9JNfvRwyOiJlNerofRGDfg/veS8c
1KCs5UbUd9BQPnBIIWc+M4l8q0xXvcwbAdDCKVfUaIjwcI1fNGbZM/CACXKLK8VK
xy/togtXzUAR+jdgTjyppbkpKQt0OE0kBYZJt6pg9r1TMZK5d2GZnLesv0Nf13gF
ji9jUHAfg8NysV9eWIqGmQic1Aiu4NorgSRXo5JbqwX4WRc5lTR1Nr0Vu1Ip77DS
dZZbDpG8naXLBENNHlwP+eYD9c7bdMEFSzmkWGGozsou84knwy3hRSRHvxrNyDti
s0mhvAnfqEcwQ8/xGdgVs2kg5Pk//DtctOmMZzrQjayVMSi/XiCDr+BEhxD4shNU
sQUCpHs89em5JNAK05prswojcaSr9KC1fnQ5FV5uP10ngC1eaN4TCz8aKLrJ3wcv
Aexl9D73C6BlbHsxFgXXcJQrJ4SIxbmBangKl7lssGAWfvqDi7K/zNEJX/r29Slp
lQZ9IvvOJOadfpr7wQ3aHkYFWK2itwl4IxDkm4K9zfuaH4CFKfy4cy8wL9O1KI/q
KrDnSGigfM2uVVWS1lrYp8STMkvK7VJtKBaxcWX5wI+00RzrV2Dgrr51MXLHBCY9
z/qVbe8xJOjE+7f084DATcRu+88oO5p5vYx/9yZN9mbBz1vGoBOmiZ2qgNqOhMkN
AbUJxGa0uNrRIgU44639U6zYVLZK7kY5KBOvq2J1vnCK9kUqp6/IVL7pZ4t7t66f
VTldflncQ3F5YaixeuZJwJfA6lHd+I+0x7xCFgJsJz3CCDsTPZ244HlNzDZYJUdh
hM6FJqTX+ArNg+l4GJ9l+wz5pf10VRpfpSnIPcba3tEVqC3iXpn2FN4taaM31jwG
Xpc3A4bDscFRg/5JCKtKmxuAnYmwTGCFr2Ahwt1HHjF7YRBEB6u+JKznLG6+Y5Ua
VnkPTunUj3zArRFyyeJG9N11feVanran/2Nd+HW6aRwpNy5pKAL5Zs2PeTFJesLN
ZavjNmuQdSn1xN6Xkt1JpD+bksSWjH65rEhChHesCrBZKVf+m/DGuTOWZjsk6jj5
iQZr979Od0uzOCGlYqKd9V70sTKjGYWXFDy1qd1/+o5ybt1KWZ2U0qN5L0Orh2EH
mU2tpV5T63lC++tyGLsraF6tWZsNZRMjG2vJnWxoiv+2G7hbRx9251eUratYBd2C
NQd9xeIImv6Eoa8TOqJbNZUXTxk1bh9sB94xE4w3dPOPjC/x35Tlkt2G4QgU2mXi
D9QkBU27lsGpN+Hj4tdmXUsxCnFiYGOPUyC/BhwRu3N1nwhmQXdOG7hMQrMtjxX2
5I5eP+VmynygjD/0E31IuXmag0JmQGhKHvlYjD+GKl8DMAjNZL4IoCXTRENEfQQR
+lHznFWceZqrkvjZ1EIRDbmL4uiwNX7cvZ1fng8rDqzOHCZPDriO8SfWmPFRO7R5
bEDCvB2JJrk9Q0I+EHOGtV0u9Uprl5rBiPqkTQ2dNGKKZ26GWVaA6vRN6sJt+svw
uVhlCpwXgdcfgmKDiXD3SKPwEJYSpxuAp4u8nVeUzN7cgxV05Bg5sguTNycJDiT+
dofF9jNCVRTfhwdw2lhSVLoX1Xf1R7eiKPCuaoYfDsP9S4f3VIeILqEGmgxzfWnp
sWeTPW2il9EAzSsg922SpCW1QBh3ymhDdzRh5Ev0/hFvpAmkkASz2Jwex01a/WTF
t+GKlT4DQbD6d0U7zQ6m4aBkRP6bLUpBSsy5yYxKO8WHRrKe6RZ32ILMZWKo5/D/
jy7wmSwotzU5syQNH58H9hiGnALOVNewI8Kcppei4tY7rAd9yeDVAVcO4MpJasRq
k053IyjhzA2NKryjhLcP48ozRr52w+uHXjWCyOK5ra/hX4uhOKjDT6Ahp328M/Es
kBAXA7ev6ljuTjYHq/QRkVZ6ZCJ4FPekQc0FpP5QwOJNd45e1+Zm/BgQ+P3uqYHm
DcOca1vwo0rXkqPnK/Ov/566jSFnZZeLZVgJ62mFyy5PoYHsdrHh0oR5K0jRJ6rj
tpeMmtPZmCl97xLitu8sED7C5k6gFNogNmi2mHb3SRlfxmnkcuvpzbjHf2iSE7Mr
Uix1m/5XJ16Mof6N1AXvrpiLiyFb8pnDBIL8UpgCNcmaxZEuV116Y6xiOtuOXJ7B
tn7TWnOUeaz0xrvvUVzH+lPrDr4Fz4aWLNkbImw7vZnnS13n1jyLLvidqYVT4efk
pfqA5Hy/sQIgGd1rxDe4P9DzFhjvyDDgF/jhyV7BTYTw00pPVvAl8qpjh82mi1VH
N5y5fGzfblxiqSs4n5dZN1Ykce/d4380fg5wl2/Vkf1XhCrIhQ1MqBRf+D/rCjx2
G149nuyH/E06QwhARsr93BBZgvCvE4fP2Moi2q/uhTNMLzVYZCm19h+1mG0gjosW
cc+mlqkTakscGu34q6FirRvaGsEe6MH0lMd310Wjzvbwrvwja/NBYyiwHT2UuusA
UeuZYo0DBHZtEPHCFzXd9KswKuHvSZx56o1kEqCp9lnU3/gDDx5SIdUR/fE7iH1m
r9EoK3UCQBLIbdppEeZ0uLFpc8o8MIug+UT3ianioLl4nAipoAW0wjw9lYjLiVkg
eCUptnV3jy/twM5OWQMIIXIKeEF552hXRM8sezUPgao2YPhjIXlSCOm5iy+E67HF
CJ+c2wbClVC4ESspanSlTfJDjBzsVXZssGMIeQYahnDh17POe51wFj4qi5egFNo1
Hjpwocx+iXubOYFv/EpvIRkjGD82SYj3S88HWiq/3cWkkYdopXZLn0bxWzqZh0qZ
E8Vva3jFNaZSMjZxCk2yPj4P6V5iImWodt0NJ+XEgYmsbvCrLLV0dC5Lt4PmtvWi
tp0cGhhXRg09ipRDV5V5Z4FOMPQpZcx80E75Q604aHABlDVL491vyO1OCT5JrxXI
9ul9+DAURa5rWuSRh4IaIjEJXpsmMn0TgzE7Y4lZu6r4GffJwNA/XEHCacN05lRd
InjjTDkgIUconELK+k9kyPqjBIRewTDUXBo7nDwiygJtvPHy5p6dZp9O4WAuLzsh
CGyNlsrp+L/lE7Yf2M8MIZSQNXitJ4m/njQs1rzQzPbZM+fIhXzJr6g0KyK8d/05
/KlQMZ+EbZNGbckHlwi7MDCNhT99pEnII5gc4/+YkQOiVZXwAanYvZ7Z+1MiIoas
QHJHfxHRSQ8bCYJYKqdASmzvyEPMYw4DL37ffdPr4MGH0yAW7NC0NbY56LO6GCCG
nqHC1ccooTj6fAAYJdm7F8arKP5d1CGFLSZmfHWdRs+9VdEgfMp1Tqd0MdGVB3F5
+fogfg9j57MGlvmcskOHyFPdCEt2eUoaWnavdie2GoWVThGyI1abugUgJb9DHOOh
SuehoLvonDwMxgapDsFWfaecskl3b2LTWzMXQmBhuRP7iHtFG6DKCCDjXt3qq2GC
+5k50ICgyVvjh8VENgDjScwYFxs63qDEqeYq/PFmzV1TDT1vGZ4BTqijDFY1ZpzN
3nWJrQINmLmzRVf9jaqPfQz1gAC+U/oJEeoA4b47jDV4kQLrNIBQX9Lg8QupZDbR
SgONMjA5uMUT5/8noQjbayyPhVuxpAXk/IIGQU+0SzORGNYu34SfHYxZ8U3Zw+5y
t3QId8+xv7x6IbGjgQhAeC0ZQp1PE4AxkJmvr6hH8jqR7LRVXzkznRBaYR6iyX1B
2d8wwQXMDTyrYuffqWrXyBNTo3lVHGRDAIo1yjqrlIuNPEaToSd0S7jHordONRbw
OZFnQ3JFCq5vV2Gkg2xfgBmOZa45LM9M09PCHastfZ4Z0J9+l6bqv05Ly9MUFJay
6RS1LNRrdfrZu9PXf29SqwbAPk8Auw7ZCryPJMX/yYBAPXhUHfAWFJZdMGNCe25u
ZA777CGAFQPzRUPNuxcTrmHI5TY8iFx42hcNvzGl0TTRU4Bso2P6o0yVvKrUtDQI
BMhFSwHJgfcgB6+EeLOIo7wtgvRBD6liiVjqCiCcwQqCt3PioqW9MVl/ulvC6y9J
YvAp+3Cn9FWQyIas9OHJ8JOIs7u5TGtrjEqS1zWDVm6JFP7+CWiBTDu3mKWCAAfm
BvfmHE9/j23BzjnGTss4QvHrxJWPI1Ug5LOb4s40aWjNNfkH0SeMsps1Jnv4xLpz
pXYTK+fnXlma5cxFt9CVA+ejD1i60IKa0ByZPppdMSPp5JSMJ0cw8z7mAt0fdyyq
YGq9qQ3j54S5WxBqKtpBdBFseywzIqRTsXaRYZQuX29yAlnjT/7uLADCjiKHe+O3
4eqZAt8Mdr7IG3T2aNWmI/yYDNjH58i7YJLs7buvr6w37dC2LgusjIw3kZpKsH7P
DVq0e0l4Vin8GcMuBTs54lGowC6bULu6j1IxgGu8UkC88MeTFkdkCOtMEJkITON+
F4XtrXwcVM4aJdJwd8k2GqGtLllBTZafgfIFhel8ZopXT1ZSZ4Q8o20gBrOp4EOg
QLiydDwo7kCWyI6T9KIlQaoxYTZ6AjJEekhbcQpuBJZIS4ruK45TxXffAB9Dq2HY
DnpideUUYzs0JXskhCUEAp6HD8xvLi0S/TTA2VsKOdePQh52xDp44FnjZaM9ORO6
yZ+rrGK2ZsxeQguWq3jPb5X/6vOqJobdQGzR8NzCNdw=
`protect END_PROTECTED
