`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQVWYjgE9BL4jwhwPlWMli8F182gUJOpSjlPvp7edHHrM3igAcHYwwzxA8usVllv
wcpufmNIkmXwkURrZ1bH/OSY8Owv0lQkV5UF+iV+YmKVXFKZzRExEYDwsyK3s4NI
VWicCav1n1JlrXtNB5ZX5nxlexFQv38ZFETb5OGZmLrr+J5HxCNf/ZMw/J62JKKo
f4zUq61REO3dak2Pz3DM/g3TJw5gWjSpncBYgVFjgK1OHTgg//7+3g0kd4mXueS+
TPDWCoM52TNBC5WK7AzilG0Y2q7js+bHvpjIOjUNUdWX3pzLJrtaaYxwAsX41cNg
04uqAonLwUIwJH8qGrbh+Se99ZXzhSOkqjqn3lbQ0J7iGU9RcH05B0gTUKWidwVs
4MLGGlLl0HkyUfqGH/Za5LFpX442PRzJSoDCRBHLvXFsrJFa5+V8Eh5ibi3IFX4J
4cks3d6Fq7BhQ9aoD6MXDBsX69++tFuvgnk4srscBtaqty5T+A0aya9sNQQ3xT6y
dnR8CuFLc81GrtyKhYwcBtqZN+riy2EIgscOtsk/bneNltEQGtYJx6LQWQ+OYRDO
G8rZRHfs7+e9vhd+uqGai8BUFt3OYoMItMcXOPGaQoW0HBmnmlnq7xh0+hABQPLe
VMQbHeO0A1kF1UwIf2YwuMPsOMtxXzMNu/aWX4rY5PWWpKGiEtZnDk7PaA1zjeAO
R9R8QiAVgLbOtz5GdXFrueqbbo+JNz70jhCzewiJBb4klBt+q1iQbXwp9Of9chTe
ZfI0Pg+3T6CX+Y3lufdtJ2kEyv4qcmvdioeLN31OTp3UFqQa79+yCyoN9PFvOCaf
3BdXCy09TdKu4uOk8nSTmWBgoZqQsK7jt6xXEmZClxgS7FYG0zGBmX5HLEKhuSTO
bBW/ACYNaAFNVYSh1Ep0ojbH3orlqP3TBofuX4YSx6afk61iNJH+hLpjIyKqCe7A
8wROcEfibMwyi3opu7gmpN7A3qCXiEWBfz1gXBNbgHx+FRTIB0m5vG+NRpx9WUKy
q2a8Ln9dYn1xGpPOrg17sXHV5RHzRR86eei9RZTyiq4K4XAZ2mbHzwuTwCb5GaIh
9TYH6lwc63QqZ5qL6KW/lP5fnTmweSPGYDqJzombwCRMSlLyqGivOzquESESvkOQ
XRKDFbLIdxKT8cL16I6oPOB8bJq9zGKuHl6D3jXzz0CDppBVyKYKZdNE3ZYTAdPi
MboS+OMxqqXwVHzYOSun7/G9r2P/5dgE32zQArcl6Yh16Juk/WOIsC2BviXhFohU
cmwi03BYIXTQ+oPxpXhZq5l2AeH9FhkDst5nIkW8jqzDpv0W0Qn3eMPCz0Ogie4e
2MQ8KEG1e/9D6xvfMX/F5oYndK396+Y2cnJen7vpmBw1QvGVv180Wf53RPSJPt2j
lEVyfr5Y6rPfI1x2SXwum+gwAIivlUv7sufjDCz1U2mnxmmQmBoB6UePQIx8etrz
yWnyDx8ZKtVeSAZ1lyS4HLNe8Bih+R9m+892+urOfVpM66KE5bGxWQXvUl71qY2R
8yvss6K9fhFBZ24c2SRqQhDwc1GRPRSdCDLheJdfKCJPemLPJcYtSqwe4b6lmu51
EV9TwxRZVue8PIM6mlIcRykOPw3eqTQRA5sd6OT0JQO5t4osUqx98fFmZ3BUXveC
4j3AA3OmUT6uaH/UydyA8+WS6NVyFlEWrr2I86yVju3N75f/YHnkpWxZFuMU/W3y
J86eYaXpotOy57GaIEH1LrwzcY7ogpz8+flm+2aIvpGvFGPEje3oA2R5naegDDMY
lfjs5BNB1JJjV3KV/5TA9VezjsH3UYEzkByXil00u0+Kk+k0FxFtxuDsUL3W8K17
VHL56Ys60HevXGphAX/PuvaUhxafjg7gGOFzVIqiwkmL4NbuTSsK8vmPoJRn+xqU
O1aCTtSJVaRFkilQh2Gs9gEGBYO1WpE6jRKEgAVSkYIWzlvIEYLS5e6TZa2gIbuI
VuywGlAnopCnrZ7tZbP551UzWVgKe5gD2oKdEbmtHT3atuFsYwm2cjYJS0TmURd1
NeeE/G5I59eW/DMbyPIkggQYdvOFK8BfGoWhqal1VT0gb1uKzw+d1rkLr6iDlboX
XyoZWbReQD1q917SGwgIoMlPsgxwDWjBcmr33P21AW9hA0O6wpam1z8684qpX/3K
`protect END_PROTECTED
