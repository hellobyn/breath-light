`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y96ECB0RQQDXh6nb2rxFw2Y/AEtCxJKcVThMpYvVLukf4IbVgwUPeUejjhQhVY6w
H9FcMQ25aSQWNl5im5ofl0ICw9PScCPuDnPYgoEqGB3HWn2Zl6qmcL5KKrxT8ZIQ
sl7X31XYpUVAzgnEPlOpwlK7U7RvoWWGHIKLOXdIgEWhKUqne45IgTTXJGz+axVw
+RNR6g86ruIr4AFhrS9fLhVnUe2OXvACxODN/1tGl6RiHbrxs3y7dPZHu912Xzc9
/S45EEXfuwGLMS6nrU4n1Fj3o6ZG+ac/ptXDpELakIJHfZI7QVg2amFh9JBeI3f7
GGdcgwU8CT6tMYd3VD3EcTUXWlefy7Tguexk7ENQTi3OZ95QbLd4OAeRYjue222S
UJnYcKKQri6u3Jx3TFJuWU9NUC7f6JFSQa0bmtBxl+5qOSjMPBQmT+4hNvHiG2cH
gCBc+/byVzl31oMXWCD14VKDQTPlQwoDzTrv2hoNGJVTVX0WH29+5rIpr5WLU7D9
httQ4bifb0cTGz0Oe5mZQMIMLLf31QNXXdv+omZ6bmJK6ShWfSdJ5AMXJlpuhfp7
a59uKWqLXqUR33O5YJCVsjidNOieDEK3B/1x3FlwMB5F1RCaDWYBcspYcQbMJA5A
1njQ2fx0aZTniuUSI5CQCzMrA4xTe2f4WGjHguO6xZnztj5celgf3rLym3sqy7Hq
Uoh85Z7eOhGUdPfy0e5DgL01+QSH3dqlrHWFb5+/XpmoK6ChBA+urSd0LkrvS3Xv
qJ2Sh7oGO4ov6j2vogOWMUaMq/fV8WFNfkHCgxWJQcnPlx85EupY0Ka9udmFCsco
qzJ5yiEus6DUdAlvVGrys1xDvbOsNwQHrE3Q8LK1bujkAUzpg52M1o6N1LKQqKB1
K2d797C0NZLICZvCzhQu5eJ/AZafgpopKBgMRSoH1k9JM912bqbolMy5vZTc1zrc
MkfBsYzgYA8PtdWblpjw79FL42+4nLt5TPBrmKbG7zKNx9RHN4g2QkXyeumr1jt0
YOV7foAjUrCaVJaUmLeyJmhaZv8grIiA5f/pOU+zMVjjkcssz4b0KnfFVsX74Vjd
Yv9E8/YI44QMFZ+cwh77zBv2KFfoT4KTmlT6tdRLeUV8sgE+pYEpAwbh9703hvFA
kDWx7+c9/3CUHdB57dV//xPs6/pnjakqczLugxkOf7jjl9wMLOBwoiM83aBptopP
MtX/iZaCPA52m990ZP+CAY0flxY5Mv135XuqOhikEplovaqKzI4UU2dUaac9vZ5L
cE8nZuZlTQsCG9+ILe/gmgB9nFvllR7AwtNDXObwIk+XPbwhGirPYD7Q9xeO/CVx
el6yYJZ9xIqDl6wHchXWQ/fe5c/IjGvv4zOtmb+aRd25qUBKuRnPAUHyj9Xwm6OE
6TYl8Z/EMiybnksqjxiCPjHMcaKvIeA82f74u2zcHWFajYmicnqlXuZ3xAOGEuvq
`protect END_PROTECTED
