`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvc9uqVcqEy1yN9sVaYrmLyTTtnx0KU6b7jWVObNUnAIswYDrZABdGjwb/PuZV6v
UoDsqKb3y46E3rSZbUBU7TqNnL/guCGHofYkZVILCfAS+mA7Eo3WV4kcjzeaALVj
EKsu6bOwhYsqnVFwvKYABlVmwpDs/2k5zgUCel1O95xwzPlDsj5CoLJ3olvzj/3w
+5lTs2BeHXe2qiR7qfCUEgZdRP+8hVOz3w2grGHcKPxKkeZIa7b1w3Pzt2PhT6+J
5udQ2ckGV1iJdl7JBcgG+vk3pIymZTWrm/jdExiymTcC9ere5ZpKMz42uBKhCXwu
u/dFCPWG+Ed36sBqZsrWCiNjFY324tS74Gcy4fdhOvK/B6EAK/UcEEq1MwkkSq47
Ks0aT9OdznlnxC/n7rhwSyFJe5rDoYBYGre8VMuifYURmNc5wpK7k/STNpZ/m/6J
mAfC0ca/O23rsZgJXWzvAq9alg2CB/5sUApHQ9brGsF91b5/osM99MAbkzM/VR++
9qeeO+v1MrWYM6VqR9hspelUNKwUYXF5bXmt7OiRAGytHT9L32io/DgeOY5lUPRh
9mLVhrt82CwbyZJOCe9bLgJ8Fg+MHCkDZ2Y9AmyEEPaRRIJ9dQFqmTjf3ee8Aick
ZPbiDaXMoh2cPps8ehB2oSAHUx8rQUckLS3ocAsDBKN3SWPrJGTstXv7sTUTIVZ/
sRGx+kN0bY8sXZLotVqYL7Q6DoDot6R8l78JtF+JkCc3Djtm6Og9ZYiRtX/X/kRp
gjngsGRduHHE2CfJSj5BuVbKJKOTw/Du+2CS0TP+GX4z7jeS2Sw0cKHTzXgRq3RL
m4Y+BzdG+tD3eMyQ2vXHNCVT/TESJpytfRY+stjeqQKx75BWRJEzmkQKh9S6WJj9
gQ4qBl8saHI3nIo/KnQHBpcJptpafz0d+4I+5H27nfj2nuz7WxlJr8zzg1NWuVke
vAMDAMN5wFgyo8h+t6Mx7dWUw0rqMKSwywbAh6edftDeC3jlQrNUOavQmIaoVQpc
7ImqThNYwt1Yd6NUxenMAfh36u6wObzrr4wIwkY3hs5Fss0AuHNaN6wodtzdNVOH
Uo1+vp+Al4G3wqsteFDDWvX1I3RjqIXD/EThpvioVE/AA9zRLLHcGPAQ2DA9Xljb
`protect END_PROTECTED
