`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
974bQRjmUCDyC8M6T2umFPmtME+sxG9WzhnTK+MxHJTBEQpZuiXNyCpbL9dTg8Tv
4X5gKuQage5zI66fpO0cxzNcj2qn+D/8cXnLtRvGADv6X9AGRT6pPB19Q/oVb9yk
E3lxCXc27on3FuS1spHaY6k5ZBRaVfZ3sKpzg2s/9x+0ySo2pG1l/DmvTVCTh5DT
Bk/tZepPEWEYajA9KoFGmLXJgmpqlxhLFcgWl6k0PchZY/eyqjmbZDQuStL8Jgki
+EJXlEmM77JgHU9LFvX74EslEX6kzr1Y+pswLATqSDtx2gIr3uscJZHIp1ysru2/
cR72ghpj+jAqSys8esGla/YiXe5EBRrCiM+rN+IwWhacRp2MFpJtDA+trIAMg3w5
tJlg8WI4Qa2hsbNclT8H7OqEAHWbhvanpb/pBV/FU3y3vy3jwZJptRhgvCc49ic2
rgwd03ZuIcxy6m0RnnHTYlfuqbrF/eQwL3xLUW29mK5KWsSa9knLjD6VZOP5r9zY
KMAr9djwaHmkV/5tZtkK6ydPMyV/xVj1CjWkWBHB6ycpmdqUQ3zQy2fJhcgRPfpy
Jysqr4MnvPi5leQX/XLxWczercezgRW6IExiaJzpy4ZtLl1f++4L1IB8he6e5TfS
cK7M+b6aMyZ0KNLPNhbkywxZv5bfXXEdrx60Kpt1bLC0y6+MksJvgnIYgZC9TQWM
JgGjY9VoluPwNfTqyMRs/l1Ju5wRJgNi9ldSNka6NZ8UXfDPGp1DxPQwUfvNXSVV
oNTacwp7n0VYLGm9CIKPmo1BcSpHX7cTXADwRTCxiPnKYoAwEFr46JxL+yKAO3sU
bLaDIWIV05PWey4evnGWFE38rRMJiOtprLaObIg//GQZNGydNqsLlw3eZPvC1p+/
`protect END_PROTECTED
