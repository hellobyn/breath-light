`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5siBG0+Z5hM9u2yrNTPO3rhKwffS6qDbiLZ/ogzF5Ip2X/0LOMS/E2lLz49sjU5o
gVPGDLE2ckqb0Vyv4EIkIUvw/XHiRmfjgZOk2kcw2vDVgS2pDbmpeSl9LZoRAnb0
+Pm8A+ykufCEOqH+x4/88NNl2nhoIXj30wi92BAyO/Zjy93Xcnp5/mgGgYRNgNub
PK+88H45+FbIB7Bfn9CXc+TEDt/3nXFF2hUhukNhDp4GNUBCJhXlo30+NfSpU/3N
fwQ8SfoGm2OgK1yNxqtqQc5t322QJP8T1U4zAdFTHTzdo3qPhLkk2UuObr9UxzNQ
02PbMOvfL1JtvD+OigP+xNwaMFSfRDBUZIInO0zxGl47XX/TBAhUts7qPD+nKubj
h990VM2NAeGkTh3qO7A7rbNP0+2xPrn4tx3FStEiXAc7PskusIja+/CYEnMwz5zZ
9YqSpdM9B1RHBTJ8xCOmc/SzGOxwCOvb+0l/VnTGQMJe1OpJS4guJIerxfFtB7Bj
qOmrQ7DDX6qCkSngYnS1ewuivj54MObALcYx7gEtBO8OI/J8/f0lojGsabj9gNSv
OZ7ugL8wYpIxtOcPxNE0enYCCSegkn5Jh/0EmLyfwCzHyEkf9mS4bnKs4dUCA1BE
BoBMf3NR+lgSxId3PzLPaaeB0Vw5asR889x2vMR61DTf7IEF5+buyZ+255csmGQ+
1kgPxxQRRsV+/7uku3lqHyX/FbjGaAukXrN1z7dCq60mcOnw0MfDdwlZXNxMSkc5
S72/cK5iwkTt6cjzmyfn8WRedpMXEguFgAs4f7QwlCp5f4ZVK9K+km3IfiYRkdQX
elCVaSl4bcAmJuDh9xt2RrWcUcX32SVOTwB2H3k8YRaOgxd7YhPOl3g3YEMkzw3n
SsN/Ipyk7Rbzi2KEmQ9sHWAM/xzHwy/3VQ2uorf8mxloLl/Lm88a21Ac6ZFFHmEE
23wS6+h8iAOzkkG71ZIg39o/8nClQY218Caq+IGkHR6fmq0GQR3N7KmhfV52yfnN
mdvMTfHvAjbp7nnxa1pfXYXygaYL5h5hx2V4eV/ra4/3FSPNslgCHX2QhIFl8qwn
4kT6PzOMte8ZZlU+gadTqnJWuLTAzDq39StjUPAb1dxGwCHcnYcOg/AeoZGQkVMO
BuD0/RhGjcPiVNkwMErSL+S7S61l20++fU1js698E4as2YDEdZ+0yD2r7jI+/YUe
PXlgFGd38pYDhiiVGFs58QIDYyNdizMY2XnQFTrt2OvxLWO7i0NHwiokvR7TkPVw
kls0ZcPGDlxVLKc+VY9BaruTAssI18+fWBDIK5Yh8jLTctm9hGTTtxrJxM2gRDvL
08ZW8QIEAi3KEMGnbILesSPMx3xD64NpgWTvpPrzAQ60fzaeQDkpV2qtayff+g8k
/oLDPIW7fJZpgYynBgTfvH4C0DDDpk8H22SFQzG1+KO5nKjpLlzPWv3OFWsxV9qn
WHgdhJecXH+RJSHjTLzmrUIshn4vdvoCy3FEXvn1lSZakl1SLldzm8GC5Olg0E8J
Y4Ev59LMTG7FfFq21LEq3P7Jh6vnzc3YoqGNybBE0knTkrKPe9kMU1EjqMUNDdr0
Ga8HFBarOQjQdF/LrjjlXD3UzJo469/B6ppsd6U1x/LpP+HnI1mcOvnmfp3qM9kU
Cmc+pJAUFKIhHBHUTOUZHWu77ao5DGn+LuIvMBd349AwqnD1+vz0yuhm0G4ojiwU
HK2bnQ4XpRhxzSH8F4vPu5FtJw4u5UE8zYvIClvkZdYeNU9pKET8zmWAe1dI1PGN
+1vGTTDlYjcq9i+e9LCXqvYsZmg9wAQ5wRQKsYPSixz/SXPKkVHo4QXr9V0KyNG9
fjIPf8C5I9uBFJ/tXNtD+gVFTI7oUoLzm76U2kAU9Qa9gC65Ad5Ir7M/jaYVEXlw
s31fHQtqM+SX8hwezwbqFUI3KQzsYDcoVOqQddBDTk3gSfYPKaEQwhVQcVWpPedw
rQiCiwPJpm0IIRPFHCKckiFKBY2cyI14acl5yuPJdUBlEfFtI/kVJee58U2EOoit
AWJ44P+DSUW6mNIMQLuTGg3RnJupCvoHU5YbR3PTHnvsq7yw3yHpJ1JrkyBya0rh
l/rBh45PyciFpp7AzEMfIVnRLHHiFE20xMRLCAYk598x2wSApUV3WcjS084K4Si1
oaSHI4qqTG5ojxIxVe53zsT+8nqjr6GrUZ5vR15pwWaag20bf1OaSAjjxgayih6N
4Mb1Gr6rOziYwrMnDYko6QITd9lJxRqKgMoTPwDtdf8Z4teTmIVCV5j1mnw1OtRs
9H07S3gk10Czt7nPiDaSSPROiqKERxulNaQoOaD5xLG6evz1Pmy419q5OT/2Rthh
HdcM+7MHK8DYDjssAgVjTu3Y41QcyIHJyAUUqw9gaCFIsfDaoKsx6pjbvWMEJqZR
HB23o33kx1J78pqZGIk259sSz1Q/iet2kmC4xLWG6vzKbvZbaD6hE7Xsl20Bf7Fw
vCSnGz3IPtCiKAPxzcT+ghAVVenOq1IeKeUr9DEj48sVZur5FgJcWQyx9Epl7neQ
wt+rP2OXMBD5bKYLAp5gRDlipGv7iPVQJZ9o68UYxYpnT+n23tFQYPPZnGtp5sg2
qmvjI8IAWIOao6jCbVWPjTj6d89O2bYy6HB8POTkasbT334V8wiBvu0JOkvpHSbG
Q81Qw08WX45aeu0+m8/E2+ExWobcHXC7i6FQKcm4JlWfJOcmYzLea2Jv8ppTVQjh
xDqYjEMT+gfuR2vEq9CS/CjqPxApF1hcksFfau0dgvgB5MEH+R0t0OqJayV7Jzad
urJ0eUXDsiMpmYO2dhw41+pPO8B9P+JIHmRD5aDNV4yH1Z3F0fZPNO2+V1IpaM3f
FeXAQ8mnkI4VDgw7QpjW7wqaA+Yl9qRATXAE31xuXoaTSZxNm9mvdIMOSBrvpj5p
2MzMh6fxAwZkWENNAenTXy/dckhDEkUU+TfUrjkfRlqm8+eL6McznCiQczJOphWO
ZMZTKDs18cnFxAoKraA/GF1faCnVJYtcjFlIbyB4OpvWXekc5lZKFEuFDzjDAgXh
UM5W4oQPqmyg3uhp1f0Jg9UPcStWs2IOGVKXiTmPwj5+fSL6uGq1nJK8bwhkOuYW
pktpAACaTWARzu0aHsYZjQNOHkzjVrzx/qcdgRK2N5kksIdJtzIZg1y2Cz64dxU8
sOWL4t8XbOwlx/VkP4upr4wsr5H1xi9JhUt4c1IQSeVCapyc6jt//CYxrVtu6vC4
l4Imuc1D1eAT7YAljE3T0OEa/cS+TVhpuzaI6Zp9X8oIEnubuBDBg14sdw1B6yz/
iJDTYWnR6deO8rXOtkDN0mySiiJ2t8BrmDl6EYryv8grT4Zi4+wosn5aU7cxHZf6
J9U2b3k2XtEFPdxp3YdfxcQBBTG22uunE4W/MoM9WPu9gfgQrxTTFqIVoZvsIhd8
vlBuCti8dW0hoV1cdKLpVI/z6L7OROqlP8VFDowYjTJyAuUaHIlt5Zw7ZAWBywF0
lQfrgchgY5Gy/5aSqSpaawNHjhlX1cWcoSVwsPRn7im+FM5tX0Nc0kThVjqk0Syy
Npz0xSTxmaprFUqa0eyE+SZKEMH7bqDmLczMN44Vdinm+HbZEfTZX8euNNqGr6Fe
xQa3xh2vUyNXTKFZJm0YAe0sEjut/jne8V/cjdEZkhQ40WkWWoJB+BktDXszFkhR
f6C7eonh1Rt3z2MNYtaDE3MH8G4ZPsfEJpY2IPYCFQExQWkJPEjnzDZtIY0zY7gB
STs9O6p8xdVI2UJ65J4Jx9GNkoeB+xhzIdhjeLFPXDWF3+jFfm0f5mTKLgc08hf8
ay9VbAWFwTuwvfZzgj+BQfnNZWasmu2/Zh/rJwRuG/hrEeof1SFhAbv9Ug7IxsMq
vhHypJCn1Qh7io/PjoLquDPzldgbZWOoWHR2PnSSx18vqyrXnCSmWuA6EZSMYI/E
VZi+GGszR5hcm8eUZfxgfg5+Vt+wAxAlCT/4dAwNAps=
`protect END_PROTECTED
