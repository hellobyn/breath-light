`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uVLl02FS26MScRnicQU8guAIHA7bcyoy2ymYLDDUIl4ON52fvcwqmL4D6q1E2XE1
wi9mVK4zUvJu5KqxNz/JeG0euf0w8kjeetAg3EvVjHErU0x6YanJJ2Kx5hch2e/8
0etVO1Mnspu/NA4vQOxMaXaZkg7iUn39z21ByIObrgrDObyASLHieJqXmBCuUvwq
N6nh9wzlT6QvzH5TTzkmQJWwag0/afLiT6btUTr3qajO3dt0hQkGPo9AGmfm+UXT
rFlrkPwd1NDEZe19LbjapESl5kckZJAWoQfL33HNuMUnXK69poOa2fEGGqASUekS
urCUGQdOxyIwRDY9PwhdtrLUfSArKZIUPMrZ1NlyCVH852We4jxxzwaSYjhao+LG
QaAT39F2yh/bcl7rL0+U14g1O83dD+EUiKRW84Vk/5BasHmJBP9EUnENbGPIq9wC
VKLfmyc0hmeeCiXZH9YVWn68CrcVSLaNpuUOettFx2ZWWqo0wdSNbIgycNgADEAp
0JqFfMrNJR78+KgdNEPmQ7Tqv+bwGN+MEkVFZK56fszJX4mRIsHNTdEzx2VweKc8
iWO9uFOUaBs7KgdcNGkNdpanf5URuT7xTMbJPHAEBs3aExuRYb9M/2Bp31TarvE9
02O09tTnmO+NNpDRRppIR+iQKo+YCTkEaI0rPqcLHiw/WbH2XkGIujVI7NjZkpTd
rEq5M4rj+l4CUhw+7GJ5ozxWfHxHsPe6s0Cn6Yt+nB6cWl1FCq8V9+Ms7Xde6N3W
WcF8pUzr9tfESqULdX2y9qcs998uBCY7058T80pGQHrCDiyz+D9yHfvfi+VTsYyf
GCeYdRZ8BKUskh/bVW8QjEaxamhXYa12y6vrASr0bny43yCc7xC2ukB5+1PpQegW
cq5FMnIBNaeMQoyJeK/oorkYA+LSxgL7HXzydaqAM/2wnylF2n25zfwSBQllZqnV
JKhs4P6bgkmfAL3XedinSkfX13+p1682z4oneEakV7LFUAYkSjyowm5cEukynJIl
uEMoVaImYX3OzLe4U7HwvfPRL6TLXevkbPQLBd2vS3ZUc8EyeO4h9IlvrtTDL2qG
m7iTKT4fdYO7H0fMUa53ATCOn6P3rlDFCc8WbHsZ4u3pVfLbluTeaBLDYlyHzO4t
Ojnnv9pxRVC26f0fZeKlDQlSyLaKTEZFpPE01qrsI/zNX5g9BxNMPRAmslFTlibp
U5PZsvcUGiDUN7FBCPPD+8WF4RJm0/CTkR2pviSFRLvfZJJvtrjax9mTGoEZRZWH
5cgdY1VkSiD4Kzgpixyd4AVBrJytuDKxz4yCpgw0th/nvtEgo0t0XBz7LpQD/4cJ
cPaiybRPaERc/HwBZ145ZzzGcJC/cmNHCt/8UsaDcej2OKund1ytVpDAW4Wj6nIO
4LnP6vqHLdkP1sOBBJDnBScxzz5OY4E26oF+2fLsB1nfrRCBDihueR95PUUdAFe9
kDuqzrf1xGWqrig2WNB8aQ/yGeYC1kPYW21yI9MozjQqB+gQDrfwwbcqEXnTLIJl
yN0SQKedG4eCzgTiLwIYxUCbbQ5qGObOeQBjkBT1wKtCUicwvaqL9sSdT++arlLy
4lf58yXXkZEDTyzF7UBFHUv0raSbimAUksmgNgNj6ji2ODJX4LX24zx5470ps3Kj
jOhPeN3ivKrRIEyjzX9rQ3yJIzK4QSxhK/vF6/N5MWnsobik97/+eQm8kRevTO+a
vCF6b5XjWq67mDUl8TWTlu2O64fccXnanFtdpJQGpcaDMft+KfoA6ffvmlrC0fOw
BRzEwwQ8roVxZjDspxfXi6vahztBtNw3+45/bwnsKdN1k+KHGK0VdqYBkF6M5d8d
mt0Et4Yi/oqR2jbuIjvTLS7YKgITj8+7apSLy1/P16myBBJl1/2CIQcq2S04oNRQ
gcbmag9BvLV8tbcqMpqDTLLKUBJlL5zyNtvX7CoxUqPuC6imCLuH6Pves81ktGH7
NxvIeOJzS6Gy+0U6SSw5RFrVf5f68omD97T7LaEdTsafy6tc18Pkt8vvynJQBW6v
Mz8cJUuBx1/+miGvkrbO0FN1F9tbFQr+7ua5RrrqQE5Yjx7CD/oElEthcpTaDUBy
7jWW0hQFfZF/GyGOPNsYm0tOp56WWaaVsIALexeFJRKhWOnbXpV21qaRMWtFLCsf
3UbeEB04oTtWb96Pa4NtcbHBFmyC4AxN5OzraZyad1BznWnOaM62TAJUTVI04NlP
YiJVX6779pQsVqQdQtFu3aaLqcx3OjrWyDN7+oyREGcc0RqIo7eSH4gZQuehsAsA
8b2SNaQukvoLHp1Ra7oBpZBVwgCnfSG2ZvCjr9XbbfOJX66/N/EO68f37VvwDiil
H8BoND4aGvDki+z4ASFD0k9Vv+FTcSnva0TwXV2VytSJzNFhTtO+Is27MLqtKjGY
aOLIx3/oxX9KhFizIKZllT6NouF7LJtEb8UwrvU6i0IXes8Qb92PZzHnqoE4fe2o
FTUKJHYkFI9FeTEEAlmNMT+NOB2pQraofrMEi7mwADqc4Am7uOkmkgIIVSWI6zpX
bpnAbRRL15D97QbzqDfg5UhGAr0d+WNQBmCd4sZoN4RCYcsTtzJI5oEZ6nshJVXi
drZqMaJrGJzByuIdU4s2QkEnKVegWJeOeMemrh2YkutzCbWwbaz/DewOaICY0xsU
UW7nrs4VVTmLjYPcu5xk18ni0pkyB8xu+SZsDOPC7nL5Ke0fYf1F//a1LkvK3Zqg
+GxeLMrLk6N7Q65YUiPfBBNQ9BUnNetf5Sd7aMBS0zzZ3eLvUhd6JHkYi+9Nk9nd
AAt4cl7FcHuuQ7FAtyuk92E31d+b0SODY2ntRGzzYjUjLiU53ZZS3rjXnYf5gpyT
zftnYtKFpbCaX/fc55TSuL9yd3MZU9iYBkgVd6gDEUSdJO6oHS2i+H4GLkrlgCYe
GprLctE2f0yhpp6DERmZJbb0BmGJ/QDV3lcJ/Ly3QtNOaFusTWfEJ6da+PwT3DvN
hcPJNrMAKxrdSjAxbC+/PnRtbQbfLfrnP3Nj02pTWn0bdUT+SjJH0vj3NuAwgPwg
545SN1J2+BdZyHUumbZUTNgmbUEErCtaQLCSik8B0o/VCI5UAPuDbnfVYwsODz96
iJqjmFteZ4BqY5yb4n35uAhD9hG+1cOyt4m46axw+7qQtbGuTdtdjpZLsWWPZ0o0
1x2AKsA7uMx50U5DZw/+FYF0hR2+jQRf+1gcLQJG4PaO7Ybc5jB61gJ8gBGEaSEv
rf8e2lrdLmSiMoY0/lPUCUdpFOrWv9IfDJFxWyasi9VfjWQb7S44vxgImploZ3Eq
idxul5+UL8i2tq/FgYae3OiWOqlW3ACQt8NXtIBiQx8nRd/L3y/h02Bc2JYz+moc
`protect END_PROTECTED
