`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0BstZ3+VKR6L0OYAuRgBfWKzcrwxW6Sd2KCIl/R9XHknW1q228ohCGVxqOh3Zey
uXWQ+Ha6uu/tYqPYyVMfGxv0Xhw4bHVBifLRxhS23Qp7hIh8X1bAG308amWFcMwc
7EhEqqNzdo/oi3Z5N3g9owmt2R+L7YLr7iG7xVA1RAwgSAbo9tPQS6qKxDEkrTCZ
/j7yu/Sg4Jeg5fAkyDjKpEcP7oGWK4bH6RQu20IC4pRchRcICLswuonYiCjoD3fH
egiES/PXR54BYLTC0wb0NptuAz7pLWiRMkiJryCGfbwMNHphs4MHEUukmEBhI/At
8apph5UNvmr7ZolvNqmL/0v7P6sC003qSlhfuF/z69v3wZeP+BO36Yfy7jZSNezR
1aORRa7CMdVDxPparQJps88X43zP4C6pCwAVYTD1PSvitz21thyzsKk1rYY235zz
/Ay8Z4iLY3CguGLX2LONQX0ks+InKHuSAmApJ/M/cfCw6QVlv5BOpvHDQB0lHKB9
trC5QS6Loex0PoiZaZTI7pUqRSz6m3TsfAGRek+E1kpCv8EFeCeds4YbCS9CCOCi
rq7aHZ0+ILBK+n9MM3JM6xQD7+BeaVHvUjzINgahNG7ZWcGjMkfuG1KT31II+xBu
OCDOdlnsEysgQhNJwImjw3dMI0GcPLgNbyxuFr9I+NZ1Q6qA2RNAqcDyXhxZkUMu
PpAhICiUTfmM7ac+ge4843iI3b7DuEPReZDRCkMQPXxDl4cHDqeqFygp2CTzvdeY
lHwaicfsotkHp98cBTZR6m7ifh2QYp4laJYLTS7YWSpsx7oUCkGIKP6C4Uq668zQ
ads59ilBljI2x/CIT+dhGbkB+ER0Y/C3wRnFvAB0oVvxSwAaj9kQt6a2DYwEIOnV
jcr0AlEk8VleUkfzYqaDkuyPgiMZ1Ez7zTzuLIeM3S2lBmuaz+F9r9VvwdFNDepf
vQ5ZbXY27MlRS7xlxZXE1ENB8Ypnrp0jNWB7JD9tHfuLv4vIy6MYFyasxTvsJOgH
rg+a3PIxcBFbs8wNPKlLEnDjXNUURJ9DKz9ypZitZvaOhZagQpOR1P3mL+h3qgUW
+pOaclUK8KwnhOmeq7CGphvihcUkYQ10u7D5pzNVHkNywd2lqY0C2iO8g4gsklHC
`protect END_PROTECTED
