`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jEF9taGEj06i5xDgrMcJLe1bxhS3OeI9/hh8BvCeM0QUjP7m5hngHRBRqQHoWNb
H40bF36M0ygtPNeTtxDq9jXbvAKIK7wRzblTHHw5qgeJt72j/LvYpJBDAEeXr6NC
5gDYlZLy5V9hKH/+WdJqipn3Ra9HKwuQpCnG4hus9rydks0ipuoX63C3dovLH6it
LZAlZP/eZ/4/V4Kt1y8ZxyFAoNR0gjpF6HETlIPQw0DADoQH52amHws90gccOZ/o
heRhnhM4daT+sTwz7VTDpimQZ0pn6tdPi7xJebonGJ7epZP3/jGyFol1VzH6Rpne
AeQEm3xE3k9ta/u4H+xO/Ls/JKlONJ1xPWueFDJExH5U3hGFR1GWNZN0d7Y7sujj
ZI0eHzE8T6nj44n1XADRsgqEyluCUrDJmZwqH8C1L7t2kg5U3WLDQ01EJBFP/OXZ
DCVlqnemxNq6m/q2pyQMMNZ7H4ACUpTYFw+3vkFAH/eHmngke8Vq+a+ZkqS3lmzY
JICXt4ECAaBnlC1CHp6I06+vlWlgINBNuaeatkkE0K+TZfsYFimlQPgwhQISUzz5
yjvZOUj6Tv6W+lqR1ymQ7x0S7yu6voylYV/Fr+xJRjjdBPioncVDdZp5MVXHxokM
key6bQY9nf3XXWuHYw6qcbKGfoIy5HGFuyoovhPLGJghzYqZiBC/O92BznxdLPL5
IsUqf0TzED2bs3lvMQWwA3854J9GqP1Uws+6m8JYLGg/tKYvvPpjW64I7kMMuaVU
XHXV/WgrUrSLN/iIrkLrDzRQm5lctfjkTbIpY81rn112fpN4PqOAhFWlo+f72S+q
JET/HdJ4XqcBsMAEUJTuaHSzYhiRHH1MiggD8C9a+lM1C/iU+uITVGRwuATfKAft
Vbm/hGUPLHbyJ8hWHflO1Q2QEB3NFtibuMydS0EdCvxODfdqvxiP69/VQWf7tnWy
1xYHZDqSRqUKIwvoZcdlaaupEUrrsRnoES6eSZXaQjfPmFqPy6GctxDEfkwEM2Fk
FGZ3JxzbU83E9KbB36mNnWvvbpWIJegztIbjikER4B4bda7f5lk0OrhG0nJCMHuV
59uKFsCPI7cGHhj7AL97MrWkHMmKuTrHxSUqD1inPitPggTt/uKNXM8L7ukBSVJM
xlWr2QBnTN9byvRFQdWBX9qyN9zQBQtt7pLFqna2rpSm0EVP2/oOkRs4E2PX9Qgi
6N9ye9lHnpTb8n8ys05f9dDS37/TwQTeXqn5dE7R1JUaBIAZ2VWLcgv8AkNM3jCE
6oAaVJeO7d+cWwwIeas4yeTwQFS+nGvlJTIw1pnbtN3n6un1jRwE4AIbCBVexUtO
Xw+BJal8MNLBdLv1ZPN1O9f1U+rSEYl881n/qLaN/Q+YxfIJRZNK9b9qLcnfDna0
t6fMxezGstZkBFaPGSLK+ahDY4UmHTmvwhBLF1U80kv5ELMBtnlhf2dONTNXUQRn
Kxz43A/yyVSRLKU8P+ZBNLVjFy0T7Ak4xxS4zMTyQkzEkwsbVwd0V2argRtOfoG8
V6Y+4b2gN6H7KEcMzGTJQ7d9FgKaazK4+XZtKY68vwF1SHN3lGFWa+/sBNX1Vr5f
bgkQNuWlaLt8o0z0Y8tGPuhou2oXQ5LrV2wLaIU3LFkPljIpcuSnGYVJE77aUnGm
jGUN3C3YN3oAZGUUo9DpX24H+MNVxwrHm8uSHfBBHBcUFI8vH1+aH+nK8f8JW2IU
6rPkCUyYT2kUT5xZFqVwX4LXKF82TOfy3sLfyze034/egwNnGtvN8CCWg3it+3w1
Kp9F8ZC2hVykxhZ8d2r6TDzLd0M2IUCctyCOplQ9PeT3UMzR0Hn0iz2cT/tna1VB
OE3V2JRh+QEEDEZa1QA+hsXx9CO3TqxANibj6wAtXys=
`protect END_PROTECTED
