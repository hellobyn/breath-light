`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3iKRYpxHExDO//N7YII7U2Z3o2Lacy/Ha8x3bXGaTzgG9cQHt3Touh68NFlYI9m
P0ukprK3N1JNojFDIxaqi7r48F424FzOsHx6v7zOUa/i/hdX/kHRfdYCydfNKyfH
RuXp5YBFu81YSh2tQDu8XVxFx3EbC6apFYFSWPe2kTF7tjOM2pU9QuZuurvWXr55
mqZZC1jZdRhN6l11vPqK/gVFL/Y40A+27ZboBMU7TiNM7V9ULbFIT6xlmtUNCgiN
DJ3A/3wW6+0uORfl1DlT41DyA9zhmEO4ZCh5dNz45sHuwPHW5Hg0D8oZE6HkOWpw
IYwaIe/1w6Ti6PMok4DrPZLluRJqcufMR+KCVMg7i216bMwDM3e+9TsU/Vt8jNZj
jRZPafaefaf4tDGbbwC99OEAU6u1ooypdOZtojLWcis=
`protect END_PROTECTED
