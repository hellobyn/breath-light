`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcNxI0SzBekJvQIxMRTlHauEaHcfQraseKVzG1U0ntQkYgsOiBCcOt/WEp3JmYfx
LuQPkIOua9TG/jVwTi+UlEw2ZDwRDhCEcgdtBvzDl4Q+vvAMeKo1oVcw6Vm3roX0
ZBtXzRJoTtkNeLpV9IpBJMG6jELnhdbRRzc55tnhHhsaeamjyzUZbvENP9kktLUS
HXZgqqYNjpNZ7AFp1QcytQLy0NO8fwCKObMAcRRUfAs1C3ZXpX5dXxESK2Ahkyg1
45A4BiI4sZxW/qFZ7Dy+L7Yqzg2svtRhEKchhJBGxOVl0wjeCRuA4DqNb5fYdr14
1cmY4XiDZBtxyoLN++qhwYMEKOT76NzA9M6RJYTWB1Vq1kK8g6f1i2szvaxo+exw
fppdzALQBKr0pfZTFHN/wNN9mmRCmYAZFqli3BwXjH6OijGI7imjNMIwiXhChEF2
Z1TYHITTcjvmyCB7WCWR73SzODxh/2PCgCvH2QFVs62b6cgmOKF50F5pWyEOhDJv
q8KWGaZAz0kynQ6Pj+5xblYa7Dw4oOHZsXM0F1fZUoHCQPaQg3+S6s3dOEOoQNnB
wN5vg79BXrdAtioqJykbb8uVqUwZiriZnEBELWaGz9fNcYxm08W/YSJB44SICN0e
BcE4sViGZri+3dT4W2rDVyB/9gswckDOd7/Jbgayp3eVGzeX39uujj6J4k/KAQpm
lwBBxJwNq64bF9ZKDOahco1e4R30yAuqVqGxl7A3AOVylWuGYwYylB3hrOFRmu5s
IFrJzRS0vCVhqejBdajJo4KgW7lMXUEi771+cG96iQM/hQwW8LfoxRd22W/g0yrs
h1+0fnhg8yikxvVC+SOSO1GNLXipVAbJtZyuICk8uc1sGyHaJHffsaR/uTMk+zng
Flrx5Ao02AU9DIdCJOCbCE/K1PFLbPW9VjQHITWhsjLPywcwoAgTrRasthkcLUo7
HHZYcg5OZevhGg2Jrfl7jTN/US54++Og0ambrmtvRBzz7Y9dSb9PMN0F1YQvUzER
e/TNvrjZv50CZ91Xsk9gpcTR694nT+0k121xdxExWCsFHjN4gjtWFSlwZZyjI/HK
iIxtn9I0eE6R9qfrHXyFv+1uzmhe1WbOJDk4zootCyFzhYVjJBYaOYCmDrR2nWS/
gaO3p41DAJlWxpx/so3X+gkbdKtuXLrWnDHRxycLD7YhXI7UwQHGg3mSdFTBN21/
/X9Y1bg624AAbP67QfBC2gx2UlX8+I9GkJyew4zA6BubRQqufyBgjusYOwmcdEoG
xNKgh4t7kZkpby+RVX1QU/jHJxtPf6VlNvF5JpLCZ4cdbpcX1hIthZUK7Atgj42P
UIO0yRveL3lmrVhAGBMrNr4cAXssBNHoP2ocW4y7ag2BbFMVGfGOX6ST4kAP6zVM
gLKtNXekuoDrz+BG7rUGY0IVlVc157VTMHTt0Zr9doL/o36X6GukEumWm9QUOF74
Hoif9qNFnWWSAJFNJRfRQslrO2J/QC49JWuupKkEApabSLXEcLphsiCvEA5+p0YJ
4iGkzIutrDSUzRbqviSADcIwqla/Fvtg6SiXYExPy7A9RSHYKju8r4iLGZPII7fO
u4mxwWnkUskRtWu4/zS7aKglvYFaF3cce7An1DRC5AD0Mdw81DE2WwOfOTYK0DXY
RX0In0/vdSHnVOR2Rs2mKgEaAIH03O7IlbDmoboH2UL8A/yrpStG2wf14YHlCxBy
bMB5mp0pZCHEfmZ7Obw+CDH5t4aVsA7SueTKObCXiCbrXFvCl6Qcob0rQnAj7jDv
eO05V8vjapy6oZawVJuf0/pbwAgfFeANCVmRdBMk+kYoUZe1CkbdRkG/AqNnOYst
PYmQpLuBUqZk5Cxn/aQt65mmOIOXVD0iVKwFFrNKXwT5+EE/wxHk0ESqV+x++TRj
azLz39+Brg/7mOtbt8IUOUixv8OjTS13te/zlX4CqeYJwAZDb3h8/M5uMqBUbP24
SVkyAvPmxdGVwraZmj3KMpJuNlZePDhjPRZbjxZdapCZl0QZT0jt5rY/wppQfpst
NT2aMIimJtoVwhZzZVJFwcwSWcYeI/4cxqQvB5TxkJiQnDSzEJUEE06EcW7dLZWl
Zs+4cvgGfMHr2N8UWGV0SYBR4/zQ5pKfWwjirBvUMutVjU9imMK3WsHRviDINZKQ
DPTh8hrAYlu2h3o0akA9QcXKqh19YB5z3cMpi11vBFQZqMfR1Pa+ublT+TngRtiV
sfEFBb85iTFwfhLJZdLrxmjfnc3ZzpUe0awTzGZWche6z9LKxOKUffygLRDJdSDU
yCXzROzGoSn9ER1ZPPx7pCeb0gFO65abth4y2tQye1nrDtsXhy5/GdoGfhzEzOGe
xfppxD5QpTkmCzZfIWyWCKi/MibRFvioOjWBDSGbKVHovRkv25uNKUWIgj+60UJ3
vfi23j00SUDM+a7XpsqFkxFXO/zYOVp8wo4VPyeHowDOC9E8AIUrhVpXbKgtqsec
obJpzzz8k4g3O1hsygtQ+CwjllwB/YwL2jmWwfvWU44RAYplOSiNwaUE1CMibn5O
rv9aWHFn7J9n8b0gsHa3AIIR8wA+WBdDPFIKmt7Y2E99MLt8OXdZaI1X2kBxyJ7n
ODFTbCgn60NVWkNhQMKwHgUzgi7UwznMU2+dwmNAmCR/2zX/xTDQxSbiRvrztvQ3
iZ6jAQOFBNnBcGet0WDi1MjKFyp4vkc8jaaeTrGdw5/nB63cwcYynTpM3sPgctoA
W6QXS+Ib7fAzENhMVaqM2HD9mTKPzbWmqby+iOS8z5+0RtgNSBYTmKySqgCRWQsV
M+i6LCqRieXHon/7vbxgVlfRy64Hu6CefBc881JBC1jQN29rK7w+KIYXPe/GnC7K
dMbIBxTpZbhV6642XtlPsxJmiUSzc11uZ+XiOmaL54S9VFTXriSIbAZi1i4pOHvy
Ii8JakNgiCIeq47wPV3xJRKNDvj127pWrJIab3Q6wZeADQgI+YFcabdy1bzp/xzN
jqMmwJUIXbkVIK1MSlGNOkHhtVXYlw8cBtbdMD15FNkenp+llofuooExF+L5BKJn
YED73pxFbBGLG9BJ5NQZR61Gaoa0x0kjaBwX9rwqNrgST8PDrfTRhJR+qjug/tmK
JnwOLCb/Yj+OfbZGnV1hPaPJxJm3YeQq4kjlLIsIIVc1d3zjqbs6VHq0OFntwls+
gGgsiER4UKmiWmPr0hIjOMo5/ijKFQgc7/EZyW8iZNTsTyfqrUNsrqEjFmm09DyC
wu3OiwlYUYirOpH4Tau8kmKHNexdlzWWUiWwyxzGHqOGz1+VvM6maYHIBDebtLq2
SKy+1LZi4tnLbm5g+sxORjFi/hRa5C1vNgBUvklB33smyy/P2INphfVYqSn320N5
KC47EO5mKwUKGiW9lSt636u5XRN+tE3EedsNfo4B/So6qyZ/PtGtbYeeiONmGb8v
5KKZTb1P3ogkWLslkoulib4HpM+T+keJMk+QJeK5ASd0Js1QXH0nYsNcSk4Ix6D4
xemeHFOkgkdhbbl/Xt+KeGR5Fi8EWDSYi1vUROb6V5DDpzCLerqDWk9WJR7TcyF/
yZskuIegXyWTnJ8dHUErZcZc1iPeazpk6XRihyzoQUrBV0HJAvkRrivFeaSnnrCC
Ga4eaznAm6sayZhOjCJIliNndqPs9ZUgsnrWftAeQgdW9GZJTNRO+guiTH0RWEpF
ECwkoJ4KCXy0W5Zbmm825yy03F3XW55V/PyIB+NBZQlt/Xhb0OKPJSs5pb7d1pKa
bWPsJi6m7l5U2zXs/yjm/C9x8k3ItiUfe9dFvKR4rhIjRzhxqWhC/XjtoUXK7l0Q
8qkxJJjmljqiBZfkgUlBYqk/azSNkgds6yCDidZA6HY62kYCqA+MJn+t4wFEBA4L
I2SKx5UKg+yZrIS44ChXLMr+WlQSWhYiEhqvqUangrjzZBUnG9Jb0txqKONCXI2S
3D+xXsDo5jbu9QKHKLhykAThvUSETvOUbaSFhCZSS6A596tohL1l6WIcZyd5uNd1
tj9Ay123rPkcXKqEhcaXgtHpxGmvH7KibJKXs7MfgYs4C+2ijdlnJ7rLt4lVFL4B
0S8BNfLqWNWi0qhguWvtJjYlzzpxtQCdifk5iTY8/w37boH4qM0eE3FmlIe/X91J
g1pvJCEDbTTxuC49o93zYUpRB/eoFhONUcfRUeaESMcmM2j3vXbideCVFO7gBPBd
Zi0rkRI0jxEskephWeJstkCdOWzCsej4z1HBlTliY8a6m5loc6dLQyiZt4Yguzz+
/OitWH44liFpVd6zMpb6vTd6ayQi2WhDnOHEd0V8dn5anJqhzumSmgJDnTT7CItq
wF4g1EETsoFght8vqEcEbl7oVnJ390Dgqz+RPKcJJLDeRxgu8SRWP82DxS0fhIcA
MTVyrW0f538iomaDAu147NhDx7oo09cVe1+YZnS1zBrFpLK1WBvTrMOsWzxB+4Dh
GGSL55e5L/0yGwRxMmq+65gynbeMBtp3uyrqaZNoCjtjDiaz0l7bPYER1p+sfmyn
HZDrdcgUGlWQ/8+xmojGbUCUIPE7RAJPIO66LakKzRGPQRfvm5lodpbS1za9DXyT
u55QkxHezHJhoGOe5vP8A0dWhR5pWI204D2vUaFsK1t0tofUPZLY1d/FnPeng9+3
VWs3GsTKGoDoelDlytooZCvI7BoOCfGY01waPb4VitHEf4sEQ1xqE/MclfdiouwY
m5sZ4jovCLBNw8JdbfVUfCGQoZhPV18t7mwsrAueL1/RrZ/VAD3BZKGG+ymi7Lhe
d/qdfx1GtxcAOMoZv9hxCzBsGjE3TbylHeTs4klJ/kwglb+24jvRQBG/qIFAAyrN
w5uvf1I2pXGEkUcR08bnt9t2liZQE+2XpaVhVnYk2dbPV1PhCmqiN+ceWfuORlUr
6D41yYAW0nbmLivTnOKrwUXnHn4ohrQNMqsMN1wX/+7kyO7//wEDawMZ+vfGwdaB
6r6Wzq/YzOdhXxLn8AOciWB4XGDMltQvFv1IaLr4FCb4EiCn6/0TBg3s7oN23HDz
ax1LneikKwZ6/PXw5Lcq/c+u2iQ4mII+3lmL1Lx8LjGrb63ICvUZjqg58GAm4qM2
mM/n7pufdtKcSaw2vc4wyhY4yeGUHanf7ZLidfRxDDpR+j0gvoGVjvDrEL/OX0T8
ROBQXdp7cNVT/vNQHUFPRApAVwFqAQX//U9jVY0Wwp9O/Cl9ibnlSy41bNrBeYEp
MVU3mufh52uzRff15D5S4yFRiMatTNC1Fj1pa/WtyLiTiwYzKZBYPYvPyUWuChnE
v9edDKIrP6sE4/WKeUHSwstzbhLmDK2nZQ606kY2dczUpvCHALpogNleds8MzeMG
F7TatIl2bbBor89ctsnxU12tDPz42tkWRE7b3IBB2i0kcQ+eMSotSOfs0KjAzsyR
nwWsJRrztRwhMgfazTNkC0j9FuZRTEyRWKVi9TSnKEUQZugllPPHtCW4+axQxHBR
3pXq+mR9gJSNvYGUee3cmF1DmjMuV6WG6LJIWqbikij1FF2cGbWAcPxa5Rgv6PYe
jqrPjyAJ2jqLapQoJU3n2L6BrvlKWWbWNz7SJkORcM18AZQa3WVesCxPp2vOEoaO
RCV79bsBrRKUiIy3C7auCFbcQvyRldmTIfd9XVvEDmljfB1SIOoPX7iQpaYl0VbD
1bfghFsL1562KeOG2CoUfF5jrqcPgQzXXcwNVo4+2qmBIC7BDxcukTpz85EmYz9z
7lsNH/bOnRKgLepIRtGpMYf+tvgNJUKRirQXNd4lqG5D15kQPSBYFUZ1G8BQf4MN
bCJ5bsqofIs4hPEa13li0LHvNdoymASd+MhYjn/dUfkIqrfUYAqETNeZk2/UsjcH
9TcifQkVNWItIJLxY+2H2UY1iTYAuRfE56s9h6wMnq2seZJiV7XgLFJz6nZT+nxf
8p+/gTC8Ms43rXfNZ0Xp4keIpkd3vRKmjAE64+Zg0JxkZklOGWgyZYkYThnt9nTw
pLUwy/hCSdw4Sz5WIqRC6Hw48jkLPzkW09GML87LgnOOz8VKRIHkouLsB1epvZdD
krwtD2zdTiDYmGUJuslWZO5rVWXR9CSEMNY84sYZtPG8IQTQbPLQUODIiBHCbNrj
AG8qQwSyv8N2530ixqtSLtIjSZJodf4LQAAVjjXnZyqJQNzFsvUUppgIxFHsj3q4
yOZUPlDFsKVeoeR2lNij9hwSJw8Ju/Pu0+/RTEiwftS0AfCND8S4/Se3kR7jesCn
5R37CCwPwxZQ4ZaUSUoqMRm2KKmXRHVfMhNbz+y2c0+DHrbuSxwXccdK+6Jbef1T
RSK3PLZE0hmEbKU5EpCjbpLDUYjvyg32DEaFUKc71i+Cj6D+O52YfVpbWRkUn6Br
AfZD28nix9QLNgBwKKzk8g==
`protect END_PROTECTED
