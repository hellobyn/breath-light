`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpGXOm5SqS9pGc3H4SFFBThKXyCH6Z3RtwiAezugbZERQiCOSEs1L6IEzdBRh90c
E7IQFrIMYoVv9t5zTftHHtGGwm3ZKGguMsLpDBnuWifRcAf9qxro9X+rpHo1uXSi
2R3uSn7+sYpvrM0fU9Eu5zy0Kf86IVAhDKZVLAgQ31niBDz86hB6yX6oF5BUYCeD
ocBN1x9PFTnSXx4RXiscJQ+1LsJ1esxmvv+NisqqtpC3hK+mw/Dg5lNHozZvCKqu
CGi6rzwuPhWHpq/0am+tDiwaU9ffxzBT1e0fvaBCgcPGLccRKtEVyTCvQBgNRiOc
C1cAt6Rt5mg0T3gzMC6w9PDCWOfoFGf5SVYj4YYnS2/7BFApnqIm7SuXG915bDV/
6HI+Kawx6YaO/c8Z8vL2SqrOGJa1HfmZIv+mHycI/8M90Chjuw0IQ4jTQdcJAQnt
ZJLLxljv63D6Ku0XkYKDKAgSNfkk9YhKL5M2ti8vWbZ9U+uJr2O3QodiE7c+wARR
6bItymu+YZPmk5/n8QzuOqDTJRXUwo7IWeZbS9x3PaxgEwapRyd5ZP/zt3eUkUfJ
MZHR+In+rNwT/EiGGsI3gbGjSp1NOu/k0wZi9xaJ/BmPpVXgX2x+PvMGDkxQdiL9
FadTzSbZpFy6ZG61QHLhgtN5Dydg1S0LgcZlE0TgdUPK7+riXlgJnHCFKYGjMObS
5X6VkHQw833s9vZAox8zr3zbbG47SNsBBdySG5eTcQ/GOI/1mu1DcQGGecKmlztz
whE55adgdBDnZ/6F3agvwngY+1qQq8JIyJEkoF6pu66x+pYB/DaadSbXfBcLdPqy
eB2jmWTi41vbEK4xusXvyTSLoF/Jgo3z6bcE+5jzRxERDiXXp0WtijBIVTdqhm43
q7vERloCXQsOweqs0zg062kbgIEl6N67AgyiIqQ2YY0uFlA5yUcUGGxzdcKil+nK
aUfovlAOS05GbjR7b8C7ksMyOOB5IA+ks5UO/Bsc8+tjUpMP28rh8juyBXHn3Po6
RwHmzDG/+kAsVfl5+5z9wpHVYUkC2qL6AFbZwWFbchFbSehiRBCtSXJ36w5zRDK7
WGgGJyG+0KcUBZoEzTSm/VZeytKPO4415MTXhJ/jGcuiSlr37vyoKrfHDGNUXP6B
9YEn7/6qQbPJpR+fejHX2y5OnHLcnfalxlevFlgvYyS5vkhNZra2qMr0TDMeekwg
uaZSQc7gOtTXhFAJRNCVVP6OS3DJqVwmYtI2A2t4DzuMVNsndxHi9AbSYBleqjHJ
mD1D1ZZ9rZCff5tjAsAjDNy37nfxbFuYJLQSoJyQ+IM9vrnx+outyM4eXXymC2h3
pkfCIEdNIzL+jHrQfe1dzRih+stMDG6pOkO6mvS34s42+mT4vDuniNs6z1beH7XA
jB0Zqra6wgQtyNhdF2E9WfjKzVTBrsqkEiOywoA6uBLE+g3wgNk8fY1iYMF6mHZF
ObTSx7yIhLCKOZiIuPSs2aherOGsImbTUvpBOVY8f4MG2MJk04ycAkSRTe18xY8M
X4C9glbuOd7PHFhn18PhLdfxm4rCVvUUKKKhKdbdmCsgcoX6FZyMx2On45haG097
dZNSWZ0v2weGuGRIG87Ky5ductel254miP96MhbGsCS4F9tsOvS0i4gZl1P/xAID
NKe7AJnqqI4aPSmUb6Xa9ONcZPhDxJ1U+p7dX/ey3gMzuOIF5Vk7wJyugqsiIAS1
uoSy9ElKhcZDh+sDOpfk5fmO39W50Cko/eze0+CAC/+6E503rbw0Cq4ntjxejVHu
kAu3FmLYjMCmy1gnwKi4jcOWqyHn2kLCnFsMWgGSKlMtRSv1Gk59gCmYvo/ACJVu
wLUoMm4AMwg2b2DnGYxv6mlSbcJzYyv560unPbfaV267z0RorzBqCfLYeBoKbR+n
jH/yLlOdzNY+DvaXV8m34V+3/b4dYOAzhGj15uhOUdpN3f61GCcQyiEhQNWPNxVP
PiLfA/Tionixo5EuXzcVhc3lj6tdrhP5kT7KB0x46nDGITRzK9G8CAks8OrTTIB/
t0ubBrF+esSCxiASFVxe8nZiJnOWUsk5WF8LAdP63Tx+MPQY+N/QCEOFinxAKn4u
9tzl3e1z5EPeiaduSR6Xo+Ey/QvNRCccneF5Ay+4LqxOZqHnOV4CpBXU8hJa24WC
m5dqlMc3kakk2abIcU9b/DCbNAwF27dmKuV5miWjv1WQvHv4JnkOWUnBw+8doSJ4
8ygDNkR7tRL3/6ebIwOphDoEC0VnwW4WltAsAKtyT0O3u+c8IbnExirB0G5Is+OY
NAliE6UXNIbcn50pazYINUg2MIr30zDYiRSRFMdZmsEEbw7f3kQqsfS285kd/qUS
VL8w2HgsWnuCy1DbAkdXzizmJEd2GrSkMKNGUVvaRCB90f+fTQv0FjZdm9fpukRm
3Kxf0ZLRgHtLxN4TnYUGXkJsUmDfB09K0bjACtjHnidXHLFrZZ5LoW0TDvdC+57j
LzondQjeU49NQvDVIQMxuApK8ciE7hSf6bR0XZO3PYhW8CveVQOF3jDTT8dDqPyu
oTYAzCgir2LhaZPIo/kHvkNwkNPYgm5Po+BVBGLOIJYLF0EXX/fBJnzXrT0ST4rr
GIMlEJ6D2ZTuHnyVBs5BIN1gRUEaYD8PImz42lqAxJX9VpCP3WoBDwYB5jZ/psdC
eUDBa2L8PyktE5SHIKjiEld7aMV5G+5G+tGjsc8TtXVr0/P/Mpmp34QidLQvWPlq
ilZt1tZmR2MFO/QyXfxfgPnu2Wtp+RqLQDtLBcYAyJJnP2c8Og/BXFRhoikK6Vmv
CmyxQZ7hr5p+zXbRareDcBeynwUwrUfcZm3MX8VYC0Dios2nIj67LqZtimj9xy2E
2fkGKbvTFkvstL/Q+um0pePDtzWnqD/ZeVNS1WZ31yWUbYP6ACnsHcdMD8PEH5MZ
IZe62Dqg5o+4kv7/u6Z2O5jRjm4sfQmFshr92pU0YPt1OJhszelTE02eKJtTcmnc
UVrBJymXjshpC5MGVpsOxmPKf2MQWDFVFL5sdvewGKz6E9WPZrvBWyRbDIoiGCib
flnsh7oY4nD2hPgiZpbWBIfzbJ611xqcbzH+395ku0MW1ND7as37tqAVXSOl+BcJ
A91JzujiU1bkb6vCp4P+IPtThTOt2Vh5zaGLDf74Rm0lNIJLrQWLY/bWb8nSj4M2
WQ/JjlfTxI+dDYJyq1hyqqeXfZSq0/4s2Xxjht7SjsSREeCtfzh9ZFiIsMjzgWFr
gWbX7iCDv/eW/j+HQUXbmqSA0hnRwnnB6ubm/T+dJEVxPBaZy+SXkxQCeqJDxr+g
WRGH3Mhq+vZZxrlc3708xBv52bD4CqRfAmZcjhT4vCG8NqpQoGCio8umHk8CcMD6
lvu/J3tXWgWUYnoLbVzFnpa2Q43WtxxpF5Ixz3g0kBRGKoZ5jLeB1hQRHPoxowj6
EZaDYMQjOuiOzkGCiEL6JayJP7nQfrzfyDMsMt5dbfuCesTyf3osdlZnA+tujirf
B+ULcKMC0jHQAxDkjZZ5kUjLDiZz2fyJYEmHgqtfgqL02TlcbVBaWh1Xu2BBqpWt
4qd03bmCLEyFHEc+cNlHD8oi4H7FyVhEjSAirPr1o8JtqMD8LSUoKf+US7SDXUsd
Xn6EijoxtUeBfEVgrWgI7O28NTS4Fsw5MGaxGgvUdY3TIbyYdPOux5DfGn5bR7Yj
wMUhXsTuM53/SvuUt/XLGBSfaTMxiPC2cNvEpMehAco/JWWACf0NDwWKrjjcf1z0
qW+F7fALKwSM8R67cNVr4KTTO5DFGUQ6mo5K5c3VjFpQnMMX6w8UvDNI1+NMGLsF
i6kc6xP8ofGAha2q8BrqmHJ3U0AZ2y0kAg2/vQG/DXjzClfmljKPFJCDl/Ft+Upc
uv6W6rGzLzfOWafAyh/iR2pmBMUF7HYppv9rr0dgfxWVw0udZ8Jc7SXxVkIEeTfA
p8Ues5JmofrBB0XSr26LeIAg3HHlN7TxFjpikPCMOwNLtQDfFoRU46PHdJ87vQ5M
RYUSSPRqhxO+nLTf5nxQdthhIGUQAQOdH6awrXMIDcx4aVO96JjJyzXhXO0VqPld
gI69X6pEHY7tBkoPELerUWN41WUESPxF/nLFA1MZgsaOB7DrCSuYuC5OH9l+aFke
QLPYwIJDQO3rs+kDFmr/gl5hhsfo2yXeY87HWIVRvBPqe5T9BsiZS+HayDQGYUf4
jVJRS2Fg6iVdArkHhkc1YUCV4RqiJmXKApRLUlWRc9xmhZlUGvKvwMAARcTeoIpy
2Nx+fFqvIA5dcjDuXGP76EcltaHVOiECCGLUNLEtgma5DQL9ru2E7aAx8BYZ+FJh
D4AslXg/9cBMKLpPiXLs5ROPUlFqvHB+NtqUJSHm4KZY2hEhw7A+3ZgdQsPjUuCx
ovSFN7hFgLnfgVVfr4VR2bUKWIuFUaXdopDkvqmcWSM=
`protect END_PROTECTED
