`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqML0+6H7Xh366O5qsFGKEw3/1/w/lPVOV0G4k0jFbkl4/0qDdEGKIY+r237Ssdw
m1yWd3Be6zyx1imKnXNTiLC24a/vhauN2yxn7YKDT2QDsPuCY43nL03uEdF/c38+
McfeuiFQ2wcEQoU61yQz67RkocvbuLAiGlOQrnpc9SXaPCAasBCqQh2R6TDPQz8u
+MZxUOq53tWjm/45WcgHLFIFI4qi6ro4c0HdIYNPqDgTyzPafnjfs1rc/r+dqEa9
woM7j3ih45q2mC39ogD3qVbTPjXEbvHoNHWzhC3ntJflh3xBre5rJex1WvyW/Egh
+/Dlo3EuolK+v5bNJdLnpMjRbtWTdJH3/lMfGYmpPbKbgUygUjFDmRvH6XoCSjcT
LdxeW9L5WEcOaCU8wVFn4Qy5+FYVlytP+IApRQD5DR/0ztSY9QRcb/mRbctj6Z80
GphjSAOxlUrRt1WmeTnP83awsbqBqTnOBK7LLJacrzkM+Wd+dJvZ/ZJrWkBvrREh
4SE0u6mRze8H38Va3SPwJqtnQBNhbHrugnSBMlm/FsmiBJrEqBCl2KzdehTVkzOt
u7oPveGdTJy7gHd1mdER7Mhtkyh6vDtJ9rbLJXLSMQ6YQmkMmUYxtIfVh9GOeFLU
tIdMzFUMw8soyljNEuK9uD3IQgUeGxSl0bXby0YOtqf+SL/TVC+lIzFDTl9u8PU5
yA6iwIngAgZZ5hAiP0vO2h+teLzQqQ/lLaAK3EKgxDMZZGXYGAJ0snd+u9o5aQu6
NtNN6NuE1M4jKoTOv8taV9XIPz4n+92WNcnYShuaXAzt86xxegtqXyKCn9igUHha
WkUgMkK9UIEfaU5QNN4U4E/QyobVHJONXxDxryQhXZFYGw5giJcKGLRS0zOIsS9l
2dPmSMGf0opso3ex4ZmeHaGVYgC2xkwkFLMi7Cyw1vvAaCLTqE9vKRDYOfNTr7tZ
XsaFmQI/twTP9LDUVQqRrNAKlPbv8D2Wbi2zKzdKp+C55a0XukCvIIusOpE92K9H
JXHsEWnbZ/QZoKljVkysG6fxIBQdUiL/f8i8fNRAalEXbAKlj9AiFoPMMrzT94eJ
mj3DaN4DGThiN7cI0NnaEdXr5kUE98TAk4XkWald1uXlrwB2W9BpeWiMjKoXEhEC
kC/UUItRcZLXEKtwxTWFHA5Zh5RGeqbZztGEzDosZARB9wAgH4qE0ud7EJ6wcHYd
Zea9CXdFJXGOI8bEgXze+dP+SDy4v8akrtPhphlUzQVrodpLplVVFELQlBBNoBHq
ruyo6q/7UZ0TZ0Br/xXl1qXw2hn2lQlOxugHaZDiflxmL7eXmwPC6ZXUYpRkMAOY
A+7Zku9wDcvGB+TZ0JoH/hFvKyYuHGImkFQDYd7hxyEP+biE2WwkXbh3/QnwCbJf
QyG0ZsbHD17bdiR2TXYJYKM+oA67xBY8dK9WjuZ9pDARln5WCEQf4EIwoqkP4x0+
`protect END_PROTECTED
