`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqVV6jzT4WrcyeFkRhmT9/9NIuD87DDKukwEcPGxZS/UgnUJA6empBpKHHHNPbxj
ILeDg5+eRdxFODnZNHIcAZ3C/Okbx/9RIzVm9KwcdHSP2yxsZjXxE37iK0dHH+nS
pfpxchPA6PLcTdrFaiWZaQJgJJp1Apt0nfoCHUGk3v54aNDtf1waXx85vC0bGYHH
ml0vFxHPlubDTTIsciFAaQvSJFTddi+SACzDhLHqd836kMTjU7NEQFSJlVGzZiEh
LGesZx7CLTgmVfWt1NZhZ7eC5lh0FYVd/j0eWRyOlOS7o6oZ1Pxin4TvZ+BcMVV/
8TQ2iD+hT6Ywj2bQekDKggmY/d4FqpGV576ecBjBUbKyRRbwUqjXLK7lJ0j6UEpn
RqAI7ZX+vP7wnXVyOG0ev8cq2uiKPothR+r5sLSjaSgF6V/pDFq+DPm87xFlkT1y
jidROJCO/KaBDtsKxYGt1LD/rWffpNy6b2q6UOhld8EWEfmqiNCCutZWUyJhIL+X
ND5cbeun3Y/2KxhKo/RH5qESgSDlXXWAgEwePZdUlbR7iTtjj7IlOSSkhldO0D9k
WRrPANoAeU77FfHylkmTXxeyFW8lPNbkAUij8EXQfqFxwqcRR/17zqT2C+lnSuph
jU0BYYiy4FQ3B9juL9DJjdQauDqHF/XIfDYmQaMIycdYEWMRh6HwUrz1iQ4dVVAy
vghvBeurU8Nluv9739EGCyr04r8QUqsRFlLWYTRL3C64IqJC+Xo12itlGopwaraz
Xwcbtokl4CVZ1l9mSYaq5lO7qbFvSJMDB9193rFGiDFcMmB50kZVK4kr39TQxBLJ
GmPVwh6b9dg+Jfs7grRbBp/6D6ejsP1t3Ex4PaC4fNlElCwRBd+I94hUiGYUBsv0
wBtspgr46/gcjps6SWwa6ojo/O/F5uiPjMJwOueHHHdKzuBNfzWl7XNIJ4KnsWoD
JAiyVh+t3SZWhzf+3V4QRT8XugMOjs2jxxI9BBUPB4IkvtSA3ZR77CLGuf3k6CXh
e+96DUcPBlcu7YzNNacY0qXeXMOF8P/CKcRPvU72faCZoAIcy99bNiQTYbEHnvUT
KeN8Dt9YGHDx9/CJXQzhG8tp5RKys7rRdB/mG0sET4Bj0kUuF3LTmpgq7Bvu195u
hFVtjpPdIAWVsxuP9r/3b+EetTxPP2lICsIjpHpKNqPSSsT3XGbDJCY8aypV0Q23
J2coVgZbFEzavQXNO8Q/NsEXByrWqB9Bu+y6vbb8rzboITe84jdiy4IF2StN0SJ7
RYubsz1Tk1dlVyklQlkknvqkdPZlBh39LZ8MXGfXbJiyNWuC8g9AANSASz+xWLC+
5Wy4lhmjiq2cYIt3VCFAuJBzN7t+sZuG5FlY2plHzGXE8aQ8dySKos9rnhQA04ud
du+HmWVLg5sVPKTG0AxQgJIQ10iyO4p9nKdFg7z1nCuFUtN7Z+30qsF2EFnHtRAG
IfrQMj6jz+xPkEG+5EQ8phzp+OoXtOhM9H+AMQz4rhqfvrStzURZLzIgNIG7mR8L
rlmGXgEQbDZFMIDsJD+pXzqGylsp1Fa/4qfZk6+8tRlQ7HxKR4U9G+jAXChmhPmT
kYcd/Ty8I+BPIWK7aTSqN5wbKM6rPMORgsikbsjjqKxuj8WQblyOMaVYrUBzzIXs
qWV0P8TBzwTZJY5oezdefOrgEYNPlsZxiTgTYRQizz20sduVja6toEnxTcuU9rRS
XCwLBIy+xBYniPKog6xhga/o3MY+j6dAQGBBJTCUu54nfFbDIrghL8FZsZhYVU9w
9duO/AgrS8ExKha1vAR66Xumfd4UG6JM5pqpCtqFBnBPVTxzIo2Xy1EhmDMSrTrl
Xkc3rvYq9+QsRBb35IseWM1bkgHh9pfzQxGFcO1O8AMiXhESy/q7VYHZ/7uDv3g+
YTRJ8U/AJmmEAWEHIjdP/f1y2+Qmopi4Afw4jV4YBcfKgjvkXF4KpUt7g0N/fGjf
dWe8oRFi8U6VURBM0k9/Y1iE5z6RI4zrK4OjKdVLHCJIJMDS2OrZvq4i/8X1aU0a
MGlfz+YXt2NSxmyNkvNpffb3+KGm0yq7/geaH6OYErP1lP1WKzR6jsPGymc9QbXt
hHAaIDWsNMHG0+5LH9DFry1kwc1qNfe9zH5wbkVNCwxZNiGy4BJl260Stf2xzyuV
NPtm8Bi7/bPpDzOg8Y6IRZLLEAbVnJwYeI/gtLjEsCSu5JLH3OYEdVGZ9ooZsunV
ZecJNSJZVBTN+RiSHFtpQWMK3l9oknc7XAYIUuI0dX3bgbWivizAbe47lOMUISWY
Slwyj0KcKw3FnMs8C+XsNLj/g2xSidY1g+JpdRrnP9OVQeiGg7wNlanHgejykN0B
eMlRAWVioNTD2m0ajgvyYVL5NtZ2HKDbxF7yTONKi7yx4P02eaA+GZS2S2IkRCKa
ofigMGgAWaYV+bKlAJJvo/QXOOoP2TwOv3plhFGvCVHnP/+tpjoboFpk2P8QJ+kd
UDB4Lu2eHuHu681Ugt2jYG3LoGWDoV3ernPWrKFHUV6P6MgLtsZBh+KrdWkDM2nP
GMM8klpc04N4JrQGxjmickXYJIZQMtw2A3z31pprMWP4t3R6Z5UI4xLziS8qA9ck
hNrJCKf+PIn1L2SPsrkXBKP1fgSHbsg8n04Q6RaE5arWpAurnylfTQPX+h5STqL/
aySq1atGvBKlqd04/LjjLuZLMIV2eZRMCXSeo5zwpQBVeTIw0VFqCO4lXxLxsQ23
FCOizdB3vFID3sbChTZxVOKLr3C76peWJgrIno2DU6owdnPow4EEb0AdLdwu9k6X
IgU7WMfB2oGa9glsSvGu6bnD9fUBZGblzaWd+gP7fuUg5c5jSMU7laVcrcc9RF/W
+sezB9TMusHaRUuCPttgE0dUtcv8NeozbEttNy5OYdp+y6Iv7rNJh14qK+djIbKB
DKEVGlOHNZvazmXwtCzdgOu3e4poDVi66Pa3veh9l712Lfibrf/gZYJvhKQJHycn
i+MgAsK63Ne/LmtsVkZ21VXmKU9ZY41htRKjFt2xW3lBEucztqRhs/ulDT/GCrk6
lY8tHO7vKqtwTSpK1PgxEI4WDp/L8JM80YAD8VohPaoTg9FGXDK1hGU3x0QMNm83
Nf31DtHlL0UPumj5/yMHmD1p2BO3sj9bmKy0NuRhYu9jSvw261hfolZ7Ik4eye3I
mfU5xF8XNsOixLXwbEtw2bayE99HRZyBavuovjZYgixz6eYd0vtxNnaDsuI0yglq
ZEjjbgWGR7kw/IZuXTL1OhiGAVDMXuTsLzVI/tSdSmpQGgcS9k/FwYV2olNkcG/p
DlRu8coTYsX82ls1kF3QGAsTBVjeMFOFuJ/ZtUngwtC6+JUUUz7HwuVz8w1uQLHz
njdPwBh3uEX5+z82x1PWte+0tgqU92ZGccmMUXNuedSXbTOM52s8O8+GOrnBP2EF
1/f5wr2io6/+FPgSScCAYeyXelyht0kmHme7m60We6PfFSODpdp8thLJtjaoiioR
1ol+Vhb0OybSruLI/wzOkI3x+Lns7N5FlB6D+0IkgYZq3Igx4KTEk80Rl9zo1oS8
SEwVaG7NNhgHn/P9MyCP6SFTN/dazWpXj2pZXCxqmCK/Yrh+WUX/bxfWvKnq7qRu
KmjoZnHxQsl8lNp6gRHIm+WvPxIpaqUw6Porq8UAoY+dYwtcDPWY2o/UuwjFo6Lg
RcoolTMkBPphjjmryBlQvEQGqgYORbarnd7KzexNIqadSzlH3xI+AUoc112Iv8mu
B02XlvJDBnVkzI6fxmttX/Mb/wftaC1kvlPrh+N0XjIHqHrcWVF3ShR2YbAeJ3oM
bBAnyd5PBISSikJW9DPv03CedwTzrMkPpktxd4WE8Jw2vAAF+Wgec6MFSWAViC2l
mu5bhTsk8JIMriLoGOUULeLhqw2c9HsgHPU0FJDEPuhilDHumFBC5Zg/QNsTOzzC
kN+YEQZhkQ91QTPBKrfjxklbs0SdjK5pY9ibIZpHSEVkAsyEFi1zPMSYKFmpMDJv
0y9fBUpAAxooZHXe3GAxWNeiLURiJ1vovMk/1xDafgqu6pbeiPr9xtW7/cRnZsCy
KLefv0Y8fajb+NgsnyUp10lSxl/e4K4Gocq4rxVapu2awpC2MWNbiTNLtHXcN1AO
Ws/p9sSCRw5JRki1dconbsauI8TEFVN/TTg3ZvJ7zyKn0Z7N1jkvBCdIznGRswBv
zNANJ5lQCJ9ZeNEHuZKuPUX3g4718b35M0oEK/PmbSP9HQsE6wsKQr1/Pw0fklTY
OpSxPysxcDYKfhYp+JG4qCe4fPCoQRI8bfGDGhCYvcEdHnUZT9a1CVENa5rDvFHj
Vya5w2030AyKSq4NI5NlE09INH4hS9hcPdkp/kpZaA4bmH7jKWatHdgv0vV/ck8B
8SGAY6/of8OiJtLF9ywG818mS6qJimh/YqL83I+C4G06wM5u7F2C+H8OyzmPFUjP
AFaEuwwu6U3nSJUnnAh5RTj71lnl32eKG+I0uiM80vT7eKDb0wUAlmiwndafeWno
ZJkGX0bPnjmqasxOjtiDFgA2q7vcYEAhyYO/EHh+eSwlzEa/jpZ8c0YAlLq5uveg
zOIcZ34xA8578j4LzTd+99vdwv772k8S6Jd3YN2eCvMy0a3f9WsbO19LsmA/LCT6
8ITRPUEKLAJ5j9Xss5qUT42OSJ6leoJupPFicDXwMvtMfzj/c1/0bM8jXCMdmoaX
PYdgqf/BZah3gi50bUQdho+OcWBhJQexG2YIGgGQ3FPU886+aouRbzBkiGUiGEEP
rzs6s30R78D09haQ19mkqI86T+Ck5WoIaKi0p6aXQCkuSuF0/rFhLBNlFpNSCeAD
BQ4MkfYXJrFZDSPdeYHnabaTdwzd4w96qVXp+bquJSbjDG3QvVs7biL6rVxHJZ13
CAg08wlDAkH4k17cYtrjM+UVUYqp2AKihI2qMbsepYNRuf8yPWYke11QWBo424+A
94PDs64TrIsZJcJhGB9MI6yyScTTYGf67uBZ88Rr2JmYwU4d3ngFX4n9WmO/VOgV
aFRmzF7hyxNP5yc43do1phLYDkVvwesFCHtWBRCei1j5cAU8GRM24tnWvjatXvrz
ItplIrtw1OxVD1wWsQVxyWX9yqOZG8crKs3WEF7wZYsnQqiXxlEdU43A9DOGeO8e
716YvIfHOGwdLTIZxW0nlqJ10HKd7/9SxJ5SgzUNYoLVRHOcpI+J9/2OWTraC3Gb
DQlZzCMZdGvQR2wC2Mou03/HCC4eMMf8SnbaVguIr4JjrYUFZnjnRXdDqDDXT+8S
LTT+lwQ/B+Kalp7qQ9cp/d5GpAvhQ3VLHlQZSTMuf3KF8UMaFMJOkUUtaTc/R/TC
JrG0HwGBiVFnG51rVN3aFreKswwNT0pwUYyFslwpUxCUkPEwNb93Z9xu+srMe5GH
DwGaNQaWkWjWY0zR1YFB1HjnXT5UhBYNqxmYwrysjdtPzIk5FTAlDWveWEfEnwae
5Ds8udnnTGaJgYoHRUxiL5bLMYPyx7oxguHY2BftJrPY0IfLwv7l+cGgj5oTbrpn
sqrDtaGmv0kJ5xWAympuC2Y/zPCF7H1aud26Y6mxQHfrtiK8NM4mFCzpdXedHQAy
o9C6A63G0ETNTWILKljnzhoVL/FZgWe5t03etrmPQwV85liTaNWoivJpvb0D0t1V
aOhn8T/yzs+ayIKkLmHur/JXZfou/Fhz5U3FTfGNLLxm81QnoCrKJymWWls/HXg9
1o9WwkXc6vHDnzAPsyRDCzDrSnueP8hLK9pr451i4oJKXxHeNzd0Z3xWOGIo5Fg1
K9WoGS7FuwFsouy+n+SCTOq7O3Cgci49Tko6wiXvnKVaOk0aJJQ/rJnZKzHnJm2i
P7RW4S55i10km3jiVKwejjJ9cXpCHykMMkieEDy/eUCUpmTk1REU/meTaYa2Q0aS
mZE8L9T4EsckQ3HgYAl1Ct0Afw19Uf1lxs8pA4ZbNkCFu+vCFw0bJVtP540zoWW9
d2xiIPq4phFjR8HaZS/G6gnyfpgP1LSKdLOQXwrjFECydT9qktqyLNTml+STFFhL
iOOQlZwJN1ZJVElCsjkY0RbBlFs81Iz7EEYhD7kxsUEuVaZTzf/V9MExq+OLqWpY
AoFq4xN7v00vVqwwDFoJMdtwYveCabO2GnDyandALr5HEAbOF8IPGM4fJxOck4gV
dKdYcLzChNytEm/q9ZM3+DDBzf1UkPeyOFlqEsWvXF3OGvZPm92in70jX7HzdLLy
yHB+B3aUhJDaATIMsdUSrpUIIoHXGwplqAEX0AfKRKdJaqH70v/ZiBkK36Jc1Fx4
oY5KCrgT8AJ941Bbrctg6QCmHgRaSHyBrIS8yIP0AqNmcxo/ifNGbmOteeM82pT1
ydjc21jOW5D+z2FC5MiG2kennemyk88pIlBixpdztvE0TkpRvq/3U71fZkNByjAA
9kNlrPpyWuAbjnnCEcnfTx5PMoELgGvqc+OCYYv5IYLusxPERy7X0gcQYYL7n7KR
oDKq/i/GPM0ilFoHufjvyODN6BXNiwtB0v36rMtmRO1b2Oxy4BA+ZiNkrDLk8gtE
hPAYVLr2+5q+4Wz699C/yMBDa08aCtGrf9fxLmjfrYNzNSTwJonHOqyCBrFVMl1X
CKGej9lvQMo0pD/O1vWIv23NwrjS6eO3l3Iy1PXHBlWBnbJcfSD7ZshptjRyVquR
DCd1CsXvHeXhfkzNHCsj5YjYfun4NF14fTB2r1AaPEAtyLUCYqTatx+ediBJ6SbC
lvXSFUa0FcXl6jPH9fRIok0vzJ1UFQmhY890anyCKEfMo1dnKmpbdqyfvy1moX4c
KT6fwTDRPCR8aJo9PiIfGyO2jrk9fBIf9osWE0ih9ILXASUB8n2r8yIThaEAUajJ
CrRQa/L5oTNWEIy5qMj0MEHWzTL01CWO0PUUXpbibNEpq+/hEZ2RhgTGQutj9hR9
yLTNs+oO74j+pt3FyB39mkTT6O+DrD7pOTK/EH+jZLHVe9pgyMt+qtL4gMoinpP+
7uLqZP1pVFFyLRPs1QpeyI16eqncqNU0Nd41CiTa7iu8O215emJyRvPAm0hJZLd2
1WCrWBUkGQwlS2Wqd0XbmCkpfYEVftE36RCL39QBiWYbWfUU4quo0eda2JFTMB2F
rgHn0YUY0s93tMNz6uZEaFoEr8r0Bpyr4EgYPV5uA9rTJ/Ko4Oj5GuZ6vGPALsqo
wKZpvR+ZQINpDRpqGM2kuUAqZMCeJfB5gr5aCe2kzCORzAplQVQgbRW21y8O2244
1LcCnCBmxso980NqFEoy48nxvtNTsIghqkHtqAB+fOgjWiesk/kXCkQebO+jbLNA
gGrNF9OXe1FVn49alrIp4OiSYH3UACADUO1cTXSp9hz7LjRpjCMS38/ctaXBPrGG
MKTtt4lmZSkzYI1L9T+NCpA51bRlvlajZwOJpKU0vfkeRLpYgmiTQykVDKzu8sxZ
PVfpUsrtAWxSBCybk77vcxttMaeFty33ANMgZISC6cpm6z9b3HyEr/+INLCxgzMz
kPGmCteeYNEQ7CP7xwXcmu9BH9mQ1vJu88Zz9Jli/Fvc9egsk/ApsQarQwbGrJEi
8QH0fHRBSLHXfGxFTEi/JCOLBrIYSvIXQRF9zA1+7NHQMf6Io9hzSdA/th0oY2ow
biqnom7VcMYXEbzMv67qr6ppbR4F5Jvi66kDJec5TEtE9wXMu/+LY4Ba6twMR5NB
nnXjKry4uItv9O36QNVvHRazy6jszMR4Gh2NQr9LeRruEx/6ja43WEJyt/9f7tK2
nke97t77xMeKv52eV3r3yB+5BcVlG3EvGuIUN7JR7ubP4bO8FrE6CoS8Yp8ueI3s
G8fpS7YOQSTIyDWUC4j3ZhT1k00csaorPavs5Mhw9KY/+4hl0MiMZRUmwBB0bMWP
r5/m+zeJk7TJihZI8tdpKfMrb24SoorjVKkATa3NcYqCjIIIRofmUejzYRxo2SM5
sG39w0E6MQhd/pJIPP5h3L9aaS5DqgAh0oqk4a4H2l0VPHoiCsl242wvlcBt8Q/k
7IJWBEWvW5EZyxmQqawZa/eJRj105subIYL7XkNxUS7MfNdoLEP554AV0JbCBiIp
A8JwG1gSOTrVY7K6xsii+wW3nxInRg52I23e57O/2Sr8mFXYkljjFo0fQ0fv6enY
F907nj67W43D1L1vS44a6XUmrMLFPHpMAia5vjWrIsYRLvrKMDC73HyWvI3ziArc
x/61xckf8NeEN2/Qp0uj5+/CkZEl3i4d2gqfAzlB7k+2rEBsrGPoSA/wa353IqF4
5yLkUi3Al5KHDYNfY1kHmkH7O46KrmlQhn9c3k5rRlLiT1yFLyjSkY4Ju+x19OqI
h8W+5lppqeEBunyG8wF2TlZspDJp7/7x071++YDWC+1PsLAf0HE/cNfsdS+x17Bm
TJwwtnDpzyht41TdBmEFetFBHE59XddKMtl7XUn4V9Kr/TZlbt/tKfT5G9mpXViH
gbv/Q3bg6aE6xVbNr+BEDRcFn0rB8WBCAHOjzHw5JC0ti7nQtfphtAtERUk3s7AS
NN7KL7ftINri4+0GaNZ7pzdj4PuGvp8t2n/aCi3eCQEM2Nx04OpG7CT+2lfw7y/P
YO255yuZtynWLI6ohlKysUmA9arO2HerMsVyA5EYC1prZgp2Ze1GULHUI/mpibs3
g3csj4jZv4WJUaGpizTh4cUV9kYcTVNNHGDErzfvOHN9LzsIQ6Y7Xfjmsd1dvOL7
qGql/DdHqSIymI6q/yPzob6NQoTTTCaiNwjakABBe+NlkVXvvJKjczC/2+DWlP9h
19dh04fA+3+VYXJu5VrLYa0F3Jr9Y5cfgS2j65oFubwQy/rwvrObeHyCxZOtm3al
0igAdSNralu74FjavS+yeRflUrn+/4lQNsBIJKcMBxFUPEK+9JTerwLzIUtzVY4r
1zcCJunROtnwQzK6wWLOqkbCCZNxPLTDJ5InJ+Fn6JKl83fqUMTU7n3jXPEHFtJC
Eipsl08tsvX8y2ihNAMnyNzY+I4M2WLjIwDk0pbbngWYHgtPeN0rXKIKqK9eIi6A
CfhEsJuXD5v1N4YOKBnn8rB4L0wRMsqqaWVStf+mU/3Fz4bb4mt5MheAnr4htn/3
E6qnjOTh0ycMp9w/QF+8vGx3bOz816yxnFZPSNP9pv4IOOxGJILqFV1u4vCGYke7
qxeaJ2YSr01e7wF/o+Yq8kv1dadPSDemVrVqyJXI5gFKjYz1Hw5Wm02aMEZVuNib
d5CJvMFeEBaT5wssfKpS8rQXcc0vfYfmOXIkIDm13czZ56IOBAQiJQlxn3538bwV
c5cebt5e4bsWuiYVY7oyG5mwc6H8H+doF7qw02RIlCuOq+opEQqvCaaLhhkx+Ttu
YOiM2dVapg1ZkYdfjSwDaHi7KrwfCVMQqAnDR6GV2gvCTnQ6PFDuBfdU+ps793Z4
oXtmfrIhFUkgTk0YP0UxZCvKiQhc3o44uIdHd5Sn7ExUB49hY1MSsrp+woeP+VAY
IARrH5/J6CvkWm+/0oPbmR6aBNAeUCMwsbn5Rhhs+jAXOg63ZewjW4nxCdmVsYZg
iblhvmW27fAowZxsmD4KYHDCCmbLpTsuG8xVdX7mhwRIXGv3fh8QhWlEznm2edR0
xJQ2CbxZLBkpqVMQ58MNzMyaEBoZmE8XcPJjYg0FlEHA0b3AA2M+4WmAMlN6slEp
fUna3ZFlB+/jWQqS12ExafzBfrSqMcs/03FIjJPzGgcDFIT5mfaS/Csh/XYvbi6d
vgT94U+JokJ7roZUlLZG0l7ICpFQ1R7pZnrTNy9dmxcVdtcYhbTlgIq58c76dcwK
9NbETz9v0UPVidOrBdigWtcn/XLK4JQOhItEbv9t31vwl+AdZ/I182MO5kHWpECh
fpAL7fheiEIKXz7+B5zi7To8xgwCFMW98j+FNiW8E+J5atbnfqH7QyK7gvEpQBO7
8xeGBHh2Lluc7/Hto9up/JGCN72dh4dFjJAinVZZ93tQwpUiABKCj6xYqW80xLJ1
snB9F++t2MxFqo0Jp7IALcjP0iWxM+vvaLPAGxs7CLjPKuM25mlMbLCyjaHSAP5h
eauzSVMZnUF2XrH2wRA0pfGKvcK7WW0jJ1tmpk7v2hYbdG4csSqKbLXa0G6TGErl
eXa9N7wgFF+xTtS32PEgIpW1r5307jlcmB11kI75ONbs3+eAMoJeJqr9MkxTWMcL
wKpGJZHvgfIs0lW2pV6xspACGVLfYM9McmLyOfzDMIAlldfLPmSeGqANep/6bmc7
syHvKqYaJTRmBqoQju76rJfNymbwnIBU+Zt7AO6WUHSgy3cpDO8BJNL9juKnb5W8
wmLqSkO44U/SmTsL30Ca1TX9E8S2qvQYk6S+B13QSwcUfg3bIg99UdMQg5woHkaz
kohcciNcesDk7MaaecF50UqGeWrOh0NYPRk4jvgtGVhpgMosd6KQlUxRuAJ0y0Rk
98Ky8AAnE7W4Rp/zAnIQ/v2esyxKpE4zaBZyinKVMx3pyabUCPA0AykjciuPDbHu
eV+gFlp/Vayhzc4eRnVZia03Jx1gl0hoz26aU1MPJK+duvv/xxSWT4w4pM3JBRch
sKP14e+6fHkkD9+vn/1L5jSecC8iGoBjN9tR7vtZjiDdikTDWu7yz4BZeN4A4JSS
ONo4epI3VWTWCKybTFMghsWcMmI8FFv4W5rdwnGpwQJLKazy9XFQ/BLUXKg1eDw0
rZXWB8yxdEbkudDxkVh6BP1ys7rCak/nTvx196KKe0yroJwAg0Ctax8asDuQzuCp
4F7Trkggd8/gVBUeoS6ngcZSYllScHPwlDU2Eki/F28zchh4oAysp/pnY72uhhW6
DljtJe/mCardgpur+AvO/Tx5UEAQknf38SA/SVr6sUMYRC569PKwvY5jHADu3S6j
9+M+vTlOWz9bUtoRx2BF4ye+PMpgk1UY3qR9656KxexsYHiiAbtnK2kUSxsTlqMf
EhlLY6BL2O/ZP0Izg1hZ7uxcB/w3QAs8Jv5CdCq6vQokw4MgQa6J4Y9eoFIq9+JR
Mn/kAEgF9wYO+5eDCtKhGbeG7Yx2G1jhWWmTDEyJ8wlBx1PvAmXyRUS9pvM+Ba/h
w7OLcDAN1IJySsnH3CoVfaVjP/kroWX3i9XvgQoXTMLgo1jhbX8yjK+gZ9X2zjQO
gpbsKJPsL+8v3AHxyzcglxb3Hr20yVAUbmw5QsU+mPIX40a46rUqu8owhLul/0qy
OeTFy2THxBYvu31hE0iunjBozpHmw3RYrzERIWJUjFIuMGXREQXdbBA4VRrXdpxg
bID/ZCOwVCZXUKh2LOgZ2QjXJg18UO6uTry9xahrAj10Gi726ckXdZCjhV60SrLR
GWoe9041+7yc+dkUcsMHj1qcZtSeh68hUMl90UEEVrYQkZCWDc6OKBZFPNOjgicj
ag6FBEH0DQ1zMcNk4i8To3B5PR2+93NiJKhOmloEGkQsrua6G5wH2ZauTm2TOheJ
IzHVBmV7GTq7irfaV85A10LTMGo0df1M61L9pA/ZtmUjvFr6+F1IYVnCa/QlNWJz
2OYX7baOu32jtDRGjRu5jaqgq2mh9JsVT/hPVfzlm2zTTBmQk00U2I5uRsDV2HL0
+BwbCrlyVNJvovfoDlKHx7rw767jv7CMGqqiwtGHYZEYu8b90F+X31ILqVWo1sHD
daRWMgzWmUFnHnN6EDEG2JfAdHJVV4N9r9uGdjMKFRqnBYVWPWMOYSavHKANi1sE
iOgiKwnDAKtKwFfSPRZLgzwsFoT3I15UpDrQoxernaFPcJbGV1Li7gT7o8IsPS3L
klX3OqaCF56CPpRqsfRYvjPD+ZEt4SYS39WiqWnUKzHb40KyhoaASacR6kn8xSPc
DEyW8Sw6Yse0qukcS3wKuqNaiHW5qYKYUQ6YbV0a8aSWsDinHC+Olpelb10Ju49/
zKgp4t8CqHNdADOBPnsf/MkMzmFafmB+lVCswJTtiiPK/QJCg2ZXqrAN45YEe6xo
ITurxZ1hazvohxSBYA0TMzBndrZb5yYKaVrtWvv0yHsxi2ZjvZEAKHT1OegwHtaF
xIzMwioERR9jsVmtUDEVyPL9Qf7VN02uKtR9M/vEwOsT4jtmCmyGU62Blfo5VyHT
RSrxrhJ1ajDjcHalWp1H7rodZ7MBpKlT6N7Y9o9aNz7UFeCezeIR8C0qB+sWRQOQ
iZhGmIh4n++m4BmC18zw2aFLfajdhRZPGcx1dEVfudo8c9OSJfpqStrsHPLuX790
js56IRkhBbPxsZhzcxTv/ZgK3PlqP9LE+Viu35ftVT6ix1KaPzyYk3knhRIv9Cp9
zYaST8aUY67+wr2EfptBDj04TDZjhnQZoEp/5C1QEz3sodNRVpFtBWI3xAwZbzUF
+qZCZuChqeBCXROx2wpjMi33aGlkrMdnvT5IadT39ybfnFdohQ8LQFfa82HPN6st
tpjul8QI9ZCjYcZ4H5+YZOazmAhnx8RePVO6mqDQC4S8C7XNQKfNhcO5ZxaEFSae
yQ2sngsUqLEkquNCCz5CFJ0QRI+od2+S7IK4HHGE/4r0UYJAqo44cjBpPKqQjjT8
nZmyCd5w+fC3ZLd7DG+YL+NvTWa2SV/h5zusWEG1Ian/7pUG5MeVofqGNNVod/oI
18sE42MjDPzQQRIfr33oNJMXlzpmrnexnqSIeAVdZwm8IFBv6XYXU8Yh6jn0xkdx
6B31HwhcaqjBCn9i7l0j/kleFEIFCKAIpcX2HLgvYjty/NTCcRAB/ZFnoKVM5bOz
XLVauVgKOdz2JXnOhy/A13SnGKC4WfN1jaB24kbiPHBAWZ6CQl5CtvwvovpqJaME
TRfjToouM/T3qzPGuDzxHlw3j2HVq6QffVhUJGgxcTbEFGZ4XwkI3Z6s0PFMzWho
05MEi61kmuJz1jSPejWRyVHsKtJ6LcewKT8uOtnfIGwgPPYkUFf0vZH+5R6fgDJs
1vOqDKyxTizUZxAlIJMKrhJFyJmX8PCNsrkbx/7KPDucno4c4PEhD6WYJhD4pL/r
eUynyXy6Y+n7LZ5dRxIeBP0uYEMRikZCiu1AfbxDzMiQqIxtbrZ2xbTpMGL6Upyc
6KMz+1wfj2cYvC8WPts79MMWmSPvwJWyZEvt3lVyOqTo12Tnap+mKmACjvoKNb/a
ZMJzKq+dVf3eF1lfAypmRZuOyCt1JXudTccHxmM1lLICgI61pNZPhJwYoSLAeuPk
Rg9UhSBukXZuUZSUCUgotBO9ldCuAORUmjS82NU6iAAxm4Z16iR7WE23RIXry7Zv
CnukJ/2Qou11g3NyNANYYusooab0GOxb+hyo+vrvDHaN3+XcmJN5RVJY9hU/pvR7
rS+85DPkhm6f9y2JEGFSphgVw07sZ9qZ5B+Mn4rkf+NByE0OIG9TFGviAITVka7B
kFqyVIulbgWdPquyVaBdSJjkN3jQFhZIjqn4m7dM05dx63mPN3e47VQU6NoeVFxR
5HyeH1utoRE6b1aAmwt9+wAK+rMvL4N8OeiRoaUj0zwwiE64YTDBmwmeP36ubNDq
dpJsi0E/iULGG/7N0xX8RnHpmK4pRgxzY981l40QB9L7w/d4OgEzJ19N+5HnJWTa
67NmtI4Ivg8osJJGzjE6TOe6BEzuM0oq8/io8TRMkJxdi9Or6dQUR3WcH2qQ4lIM
joOk9wp0/QnvWySJ7udajDniu/Mw3Hv3XQh7Qa0+2HfxaQMlyNxLYi/B5mcrNRPe
0F8QFzDjLzn3JxSqQu6ajO+/2ZfR/ZRJtrA4DAg+L8ImAQA8u+iohXg7VH8t/Ljc
AOpedakh6ySOLhqgjZfs/FBgNm3P4j1GvuNlkS0GwPMPZDqqfleIbBRe6NDVTDYj
/d4NqnUY/fpR4Gc4ctcPSlrhJrI9maGd+1ErdQ5fl2zoRlLxSlOnVhi4CZKQ/NDx
AnmeegnHBW5XgI2NiT2/0PHyt68LXSdOPxlTuDmn0fwPhWo5nV+rjVeDj4cf3KYz
BLlCqPSFkPEwVeOkCRvgFjNkx4QduXwOV+wiKKqLbADhl7T9yJLUP4jmU235kpVE
yeO99oL0q0mJwze+zKBaEHFDmzzueXy/YvmelJyWsQhmwQb3Y8YH0jVaP1KQZDvE
tLFD54j1INX+ejoy7r1tMvne12nkHpJAiRsmxwZuth57yTLNdH7img19eCabeJJY
Z43PloF0OK98/wYvLP1VxKeipQrvijGxC/CJW80RRVxOtj3svAvGLcL99r/sRgJy
Da5iqyYkmfAsGaylbpmRUJF0/eXX8Re+3jw1UDYMM15EokHXric234qmsGxgkZKe
gp6EA9VsiXDAIuWSnvRP4HJqNgdZhzIfu/pa9imzWOauVivMB6rdPS5BnZOhowsx
ATjNv4JYVXCjc00ZU7Jj2lkCUor+qxf/7HKVQEFNfXm84dEEdIN1PLZjBHiyT+3u
BOYUUeziHHnLAMmFrRDpxgTIS6abK+QC66pmW9d4Sb0CJFUPBjAJ1iQixQu5DeoU
uc9qFGLBtVeZ2o8ZE66RgOKR/H9LmGT77E3YwcBqDe1IpPxsCSTsO3qNvgBl130u
8JB8fcvsxyBBrGiQfAer6+cOV9EjLp8ljKpAMZQ1SN+RFpsSr/sfLYgQ3YBpDWiJ
WYf/6cxNFng3+Iyfb/TqyqEzmPzxKMATSW3B6+xepLjYW4kFE6C/EfpkHJhtmvSL
BiGyZaNzM5idQLVyAxw9ZCo33quyQIZBbebgQ2RWw79uktCGXbXgPicQtH5xVUPL
b7gYus4U14UO40DlfEnA28gT0LO9FkoB3SzH1X1HfNFCLnaHr6AZVKCWcyJyR6Ee
EcS71au50nl38kWP8IutY+s6lIVPzk8YzlTUJYLoBWlZNjMAXQRvx1qEg3O/MNBl
PzVNJVrQS/xk9OxdV6bY6ofk/x9JvxBgghycX0tfPS06YWWwVnHtmdnVt1dban6K
jsFcO1tBv2ymNlNeH8mO5HJpO/k8BXj6Ese/MaLJOZO0ZcytKczxoWuvlYcd74uK
f9xlJQ/4xTa/BuCDoZ3VrpIgvQSsZGjtyD4CkYrzSUTLlzzrkNM5tKJSAgx7JcHx
VYL2usSMhBS/MenQIm2RMGYBx/dMPCREYWz//TOA0LG35Os0a3gPCf3OM2fsQy5v
YQKLN8puHPDwmiuCMsJZK7H7r6rbtCHXeqZtOHZRHpg87g09ZHtnwv4W/JcxcMu3
QcwPbIm/JgU851U6g8mrm+1FjouhZdpahAoirLbvmvvs4HMQqeebGyt9e1aBAMUt
HY9lUZfOfS25jWq1Hic4/vlLCybL0DAzPfJID0N6kmr7jeFKYBFQk8ZF8u6Xz6z5
nSOz1Hg22cbrijzV+WfX9o3MZkXL/b3TGFxPOyYw+oQdderOu66K8eP07n6GCIh2
QIZlHMoWvmJn6YJokephbI5r0VSf0INyINRkH+H25DZuAJUXTmK4w+gDIwsSTIwy
ABoHyFFZ2d860yn4+lsGV8HNUN48hCHTL80AJw5VWPgvECpLTaRNXcUe4rnWKSIq
KXxg4RMn77hiKj4ZwuPvFFJOPEGl7zoR4gPNNRPMustUUlXLgcMYs8yQ633/jvLH
AhnvQUZQ36Lk89xcwW293Q3s3qCJnorqnhullhhTqaLnpEbKHaeK304UDr+b9REJ
tw3jUveuLvoxeQIZNBo84iOeI33pL2v8pBUjW/Ga/nRwPFgWdL/cp4VhJ4d70zCU
wZxKv9UxAOeRAbugMWQY9qjNQ0WFh0+ikwImk339P88raT7OMEp9ostdqIdY3b2Y
vGH6EiZS7+LJgboTFC85bh9PwO0Pf6L/tmPKll5ksz+paM9t6AO53kXO47lB2woK
hPK3PwYfQN8PJOHfBMFk6ogZVR+admaGd0vZmBHEE1Dw8BWbVYK2pEBMGcOJhK1M
EJvzs4WSDnEEOnFRlLTIPCWH6e/2z3bLTGucOtNgtrYJCYGbQaUPIIXdA5nAmcnL
ct9ljDOc/croCfWGtfB4QLNJJQ7Li2J2QTUJ0XEaBOFYGUKzq5UyXLV9/oiaHqjU
QWNTpiw+aBJFUy3eT98RC5uWdAPtRTJgjlOKHb6+DfFAiPNLNnwIfh44X/HRo8Qw
5P3Qq0dFjEg5AZy9GLmg3OATEKCYhG4MI3QViv24bAN+/F69IfmEjplBdsBPwa64
oG8i4ioeHTDTglTyz5WuiiytpsNMDFjyA5fxUBLILFI2wBpsVfsRw8BobFqr0Uq6
+yfXoBFKTjCi2JHn4ujNi0UCemQ2WLBFMzpWhHSQUctBl7Pbe2rd+QwoY7Wf/WVu
mSIKx34DxHF1ekwZ3NjThb0pXlphctyCRXgndae0ZJu+b6f8gSCUA6kcBfqOdETi
gx8Yj1ClRmvK1WK9E/LliIhLSQaUbnGq0ge/jWTui9ZFqECExSnishYTp2hCXqPo
uozr3DaCDCXUyC1p2IQMS8O7IQS1YV/Y83XRpW48TJsegJGVbNmp6w9bWGqz0qMW
ZjFa+J2ob+bbSpTduV5o6dWavas9EHOvC5d1smAZlUqGWq5M1BUCG6iPmj7XE4Xn
w12xsyMYDBikpXGM/tWecr6lyIRsKGTp+aO2ejeH1cXrcLAddmlGTGv7cN4KDAhs
HuN7ANYODEDAADM54F+vLrqYltq564bcBdo+LhoNeQhW6PKyahuc/SqJ0DKj1dfQ
5inv996fNwSN5oMpZHHmL7j7CFOBXwPMsViapKkZKkHH+xthm/uVE7CpIDfyMzS7
pZysQZzRWfg7uqfxcniFFVCkgca0pZY5Krffn3TUGbFBGUUpDWdJUW2iZeO/rqyk
ywimHL3jKN+hcipXaMnPdMYE96iRDipi8PtHPbctm8U3R5SCfmjd31OLn1kc3PBi
VsMYKGM1MHp0UTo9haH5aaXH7Q/SBbNQGJV39eV5sihQP8DWyqLZkrNsn+7iZc4b
SwrL0g5jV9y9SkdBixyDLj81B0FqjUszbZhTLsxM5QvaJKJNFvY2nPVTGXNb1pGe
fKCaMlDfX3pRF61oI+uP4/98uvu2qqQ/WreK6QnkX2DNBHUnhq0pMR4wYy8u6oUu
bBfPif03MGx2Sa1J1ZTKSXwVCf/rkT2ihnMBfvDyw3HAEX0sLc94f+G70Sz+s7Ce
Xqftp36V8+SSFEF2QvomZvEXw2ELghmtM+N0Nm2UtOMYdN/PKzUtM/zbThxv+XVL
R4q2YGNfw1zJBiLrOtRYMMqraLVbM+oV9lG4HWAO1a+a1Hs2WkN9U/YyhzGSy6gY
MmHiX2jYnqxO4Is7+g+qNQB3V10OVYdUEGvT+q43DTh9JNVeyjK8DGbcjjehwmwL
N1UN3cBSWrtfke/wxiTEVq+ZWceCvsNWrvcTERI8omwCpa4BWBfSnF5+gQn1+6NG
6x7CaJ7GpRjjff4wY5oiUX3ZNXLUUSGBIT3z2LKqzd4H73UQA3w1Hm/C7YC4Fm3M
hok5xCbz4X+H010rHQS2xNpXKvvUHbJzJwHeunMDSpL29BcNuqgX2/+x4nxZRj0B
wNQChsx2P3gI0mOweBgSH09MLxC28hytMWkXg7ptfAPrQMXJI/dp9TI4SJ6R7/K8
V6+hYaUc5GWjQeOuxviolDbcvQrq60rSolhc4C4BQBGNjlRn9O0lGNrQnPBhmggS
JRQ+krAGOmd9q1oflara/W98l/SiJFLD7lUrR3+tDCp3qFXscv93WTQZqxyKcadD
yAJVyz+R2QwRLuVsmnRKRhKP/74f7fFqKz89jCBD6kbcVoJThJfAD5ZA4fVoBC69
WtBxQ8kP1sDIryh1PfIDpi5/QbUshDcgFiEQk7mkGuQZEL51DHG/NxpVp1yTJdLN
7qLIeafB5Dyl2BqZsDIbrGNy0gVJuzfAlPm5Cd4tSUMx2Lb9LhM3BSZegzZJDtBD
F6/tF/t3+VuEcmVVZt/86lRThoy/1ClqHZISQGT0AtvVgrdJgUPtgMz8CyUFgbA0
tXqRQTZ2GKqtuJz+p8Vc6wSS6iMmNysVGRyB5Qek48M6MzL2h/HIveKgCOfW2Ez5
UQZ7PFVD2NbhUGWJx5ykpwikVDymmTAiuYFivupsv6sNQhVm51CdxpRChEvuCqXE
+y72WQ1M9l/U8uZiBRXeqURBDHk4bG7UDDvrGe9a4Dli3bPjq/oIydBr64eBPNRn
nTyiyHHmGmsRKuqLs1eKUpuRxvYnpyl/h98Wdk8ascll2OwyFEJw0OtZjCjzBU1a
a81FlAiSVuOipkOkReHWU9rTOvJTjfosNo6aLv9gVIq/wFfs/mSYA6ZnyQmxM9WF
CCic6XbyUco/qAekhojG/qHo4kXcAWjF9gOKALWrcF4SQ60uU91PKGn0R0N/3j0W
wL482rcs/1/EfwPOe3vXgviGzcR5nrQGOBxnn90ZHTMwETCrz84QM1UP+cpor43E
mfP1DUuBFXp6eP3wBKzSWdXsC5o11m/U/6GSnINHktHI9lS2QDYPk/27+caZU1Qq
+/6WAvx5yn7NWwK1vY+wHKfeV37yn1m1ZKOFOUktXFCAJuVxJ+S1b27gOu240beO
MMoWBkjcrR94soeqFJI6S6PnDoL/J1DL1sstcJAVg3MrRKJ28Xqa+zUu2/gT7Sea
FbaeJ2+qOsfxxDNzHV6psa87s8eeEZS7YfZqGealar6UbkkbT1m+blMIuIRpQI4O
M+vSajeK6KI7OiknBwkdLr6JM0fYafgmGbMM76iJ3S/vjzTeuw8FcBnjWZUSg+sm
rp+b9AXNX1IfDLbFJZLlE/Jh8nR+QhXyvKPETULxXXQWVfX9sbI7H7lwu7dW0g1H
qAkeWsYc+zHs1WAfMCQAYWzBuID2VYq42OHocxHKiIhcK8hPefiGzVx43xcU7n+M
8zUvGruLEVeXI+lnnu95/nnbc80qFhIakCEYOecEithWvwzHK13lblOVOWiOG91n
5hnyBeKaGJSni6qo1R/ZziLiAYg6e6/D1zjfOqiSf2JPHt+lN2+SEiJpVnG4gyAO
u7CflgN6uncU4zhepD2WgpjTTnx/9CgxA9hKnezjE2o83zFBBbfCgCgsX6J+pBvl
iFM7ejDx3uYQFKjQqfOQWKRdQ6Xx4XKSrGvpCICAR30k3Ds1c5MVyGD5Qxo5B/Tx
lsjFZvslD30vSL3DNU6rOFFldEFa6IHdCJ5EAFOzFl89fT3FxYJx3jfFJC0VklNw
1u1EpbGeOL0YlsNHCtmhQsAhoE+I2S2Cdkyufj+kSHJoTsfsT5lnyz62yct54c66
86t0aJ9WQbjNhG5OMNa1JlZwhZQOsXjyrfCsCaNepv024/VAJEGKYjuPkNPv7b56
tnC28p7vKRwGIY/KEKUWqLf4NfboKtt0HMFfTs/4+8plAIKFOZe1HbCI20m7LEX6
xKQwwiZ+NGQqrMRq/q8IIYyEn5rcfTDSPZ8gwGqliztrLpcXmrjM4CCmuyCDjxUr
FJqe4rzLRy+6wA2MfwATKAlo0CSl20kzkNN1GrtOnIWSmIaGb1qMXmEUjKT4iub4
1ZaHzSGSIUkM8lebWPcvwEZsh9HaEq71pYb5ggP8f5hCcZljEQv00JNMnrP7+tII
j6TyVOOTb8nZTWKuHpwbd9cG7RawZT3Va8rj9Sjmw1dJ4gOHpEXf2Xu49yrhw4qh
YRbBmcAmo9bqRvVmp+o3aAfEbu1rRLuPStO/XOHo7WIwT03F5eWfN5yUMqjrKSWq
LJtIyOasc4GGIJZptciolyD8mEjs0Dg/1dE2rsMgf3b8fPmoOnj3j+Xl0JSE8SC/
XSp+AXl5klUvZiCM8OiwVfbXAU44Xq4nOTJ8PuXOb2bbaZ0gL8LlDR1F+sOx+jra
pmk4Rw05J4jlOgspT7P8deAmiHKumEwXlWFxGMM22DazDxaPpaCwx4aupKJhJNSV
oM1sUBv/7KMrarbI+pjLr0tHP4Abn9TmgbrWuNxdRvzOnn0m1Cgm9GhNuwW+l6GQ
MVvzAaE2q7LLrqui2IGIVhyhl6UZsNbHgtv5vK26Nqj7wkoE1oMZTuGjOvuVaNVu
/Htk55KTxOU2/CJUnOMeF4TAUBZZ/+aZLT3augTcSWBWhQKpSBVvoLVwM/eOxxiL
LHtmzcsJUSRiq3AXnuQfv5+CK/tZKwsKI1712PEpNAVX7f/Z6EvzZ7hX3mi3ewJM
Sl8Lr4Wt+be+ujFsVJTmyQQM1B4NVrDzRqLLUiah/syZusy4nIVlMVzKa6Ufrwnb
Hfu8EeTLfHi4VfsH8HQogQw2L5/8m+2HLZl5mKP9TQv5NacQZyXw8UNTVCHMOVXa
VjyMy7NcDu2iH5tm7BbQ/KtcnsHcfK5ZeLod0gTnDah18QdO/2GAy4dzw5zK1kDe
TCRxMgklOv9WkwjBzpB+l5I1gTvgaNMnebgG6728b/xZG1K6adI6ds93LFpEzV5R
9N0qt8Nfs31AmZ35B02K8bn6JdAm9hZut1pV4Q35zsAx8b7NZ58YQ9Bki6oKwNQ2
f3AoQH/O84lzspgOtMjlJFraDT1obDEruA8Sp71yNIv0eR5ODKpg7d+ONq9yCQVf
xb62xEr/2dmCK9ZeZx27ynwE0somov34a5adIaM/9Nl3/+cTJh9zC3uWgzbEyjEE
7CXL9NE/0NUeQxj3rNT6cGsB2cettdoLWqnZa9ODxI/CLPO4KY4sd7aOMmz8bT1x
UmP9hIZbLHBb0QRARh22o0eBZwwDsAPvsr5uolB+Hti6hmKe49jNQObiqrkMlm6c
dC6tDavL9UeVazQJEcRb969A8MJP68z1Olr80zSgXJFZKwECV2ST17j02QWeFTCn
shbJh7Chx7JMTXv18MhQf4MNwbQ5EXWXcFH8GBkr+upZ680WP5UMEWCpIfpw8xT7
XSz0aqTVj3SJ2fg7IgWLtEDG2dkTcFNnqEyi0tsxB5BzJmu5a7+mr8LOzQers0to
19hycHOQTVe8x37Jf3mpohcaG8wfTrxfb1IMdEJtWHy7KMMakzIGfv5PkR8c+s7a
r904LKksVC9vZRbTyNs4yHNYGg3o2BWuCB6C+BZWJGgrn0C7XQRbChL20uskM0oU
sHbI3pNgnYERcuTgXw9cVUoQ01+/Ya4t+z9vtMJYOf78AranTW099tuvfwamdzjR
HWEkLbwFte/RMwaHqRf+fEBfZp/LaVXGN8hj/KYoW1L4eiaAWvkYV5uEKonc7Zml
ADw1pw5G7olMWCYs/r94/4ZLGgh5sdIsns9FlD/RjBvuJuUmNFjfFTcO2CewNrkJ
Q6tCzEeL762lInLoLRmM4bStUw5xCLmY14tRTe48pPrweOQ/NiOveHOl7nQdxtLP
+9XdRMAJafbsdNQk2RxtkD5iqC+K6NoQem4VCoFQyb7PBJh+H+aE2j571yqeUXcO
AEvKixkwtb6pWF2zKQGwWhkIOfe8y9KpuKeFRkNlQvu6tST2+07Mz2k1IRl+9KHY
XjaOGBCLvbzGVqvKTdfm6BaPbUTVy2tvTkR2wucwSKB75VtwNmGthgoP9hDJm5Q2
Hy9oniSRyjoKIawyp0F6H67thZRHPUUvW/ocugJgIwZfFlojAVb29vjb0gaZ8HAr
nDaZ5H1Oxed4hYj6Yvg1dBWiQt4FAsbevPKN4K0spGqHMsCqG4dZy4SeJmk9TF37
lAf59GSEinYa+jKYlTNJt9Gw/oPWHijOjH/lVqJHzOOQY5rxqia533MxuTJqxtbR
oJYPjoWZ4zxK2lvLjnf/6ZEM8hZio6XNPeSjz4VrvD6PcGA01GlMGzuWc699Fc13
Hm5wfi08VBSkJqU5wmOO7XrHxl1AGr6Wl/xrAkhsvnlaIYH/5Xil/JU3bA1gV+hf
I+cCzg+4icunzsKZzL4NTBIREx7VFu7M8AV3J0EXHcctxez5cZZt4Y1aArb42WxV
x8EtC+nmNImAyS2O3hXJIFt9tI1vdEhTrIsxhCqO3skY0u8p3tTzQWLYF+g5BSQN
Eya4DQ2gWbyn2z1BfqU6j2neUT1whbHBi89LRkBiosFEP7Rafw3Go6i0QHiItoHC
u1SmzYtWDoLnzh3/41cxgH1LBi1SfuL2qwldF/EQUIFe7afOI4ZXO2MWzGu0US11
ncUuRYgAZLvv3fkUF8O1a/LTC3+alJYa7cgUxftQnZTwyQ2z4kNV0Kd+POGr1JQz
0VVefgpYWVcHB2dPiAiaOMhzYazv88QoeK39/So9GYpWaY7840Qj43RvC6mGuq2d
nU4YcOycCQmQXfhX/VT7ANSOj7kh/LZnLpW4kUHgPaflLuyDFIC6kMr+rucx8JFk
YiaaIywQ03BckyT6WI5xuUMWKGkd4+hquB2wCcIpQUsxhhPnPfOQLkr6wuZg/wx1
eg/YVOtovS69Tx+gYuUgwnEAEHXVNGetoTsUM86hAu0df8GkknxmPEQMdVjXfU0n
eNGolwH5qY1EOYvA2/u4GLC71ECVb1bhsnz5OdZ88qZnknQuf7PeHFSuN+pk113R
uJJha/6LLItQ7VhXRZbDT21Hf3El1aSxW2ZYIAioL8oMOxmNRGVzxZi/Qs3Q+lMN
p1Yd1QiYPPynRVqZeNopMUf2C2o2e/2TLTbshN6NvzjtfE2pbolGrNb7Iji1p1ms
aD3X6lifNXTv9n024g33aUVvOpaCnGtbzaaoJGu5SZynPwCVuSeQeUMgUNt/Bq8u
0HkdxfjUS9Rz/JZ1IfNk2/oRbxhlL3PTFbO0gIPMQytOdBgdAfM8WB/EiJG27KGo
gSJy4NZYJuMUSGCHWeyQ4hvaDkmhpf0rzWVHq+PLk1rgJVQywp1q2ZipqG5Qe293
sxF2I6f5spNbknTGHIpTXtpOYsOdsOK5IaEtbwPYS2H6gIkdJb7rCodghtDvjHeZ
r6E/XeCNYSi+yVpmDDGX0pHmXBvcfIioMm5WMzXEP0diOQnKjxkHrOzADmwCwr5P
Xo7kXsuDC7eI4p6IJFaoi3jbk/sAOcCxIpdlyFo2BPTzuuyU/d2GQzdtaxbq99cd
TA9NN913nVmc9Y+4SmhMH2wHlAecSz4CiuqmMNX2t1DS1Ns3eBTTG2/5ICb1Ers2
A7oIe7e1gonoNTZFDCseKj7mzjRkoleF2MSTt8QmtXNpMuOkK4GWnnkHWrk0Y5H7
AmhjPNNIOzJUXsjkymTuRGvYvWNkHtHoa9pkGC+s2FXbKNVFNURHRutwdkaxz4u4
gLJrGyUbmqW27QwWOBbUfTSIKMQHS/IZSdzUua5wnvNbKdCih+AC/EktSPn1Ge4e
QVExLUAJoeo1fRSlQ1vahYSKLTucCRZO4tSWLfDSRgns3GPgkyPVvofivQlwrfSx
N21nVBOpC9WZbtWIXPwbTC9cc4TqxTxvKiC0/ktf/ZkgkhbKdWFbsET9oqCbfFcX
QtNE8tQKl/aQKscx1EEXQ55pt8fQUyWtDDX6tNQ5J5DXKyESY6SGtd7B94b36fZW
2fr1AMcaoRAIGPbwC/Mrg0s3vVWZnI4tfk2q43T4MYd/7VVZg/pKGGhzrLmsuPFb
ZXS8hVPN+V2KPlYI1N+fYhFeId02ES9JCheEhnZhFzSHeF378bviDX5YK6yyL1Kg
NExdaGRi30U2MLoT8RTdUsLkQADb+PvuYD+6n7DP6n7AyPULuswF/GFBiSLBsfku
z50AKUGOVrb/6OzQPaXXHI5qRqO97Uq3+qOtcZv5ZS1xV9/8Hrl0dtflwgctsp3A
cz2XCb8+VNAbGIHupRQMt0yzO3AeSQxW3vUxpWH0z7f4gvkTxbOfhnpyzov/xt8D
LmVDu2/qn9sqnq/A2lCzJBXnidyykZsTtl6g9GqCofNWbl1ME/v0+tf0h725j6pU
7O0/sleakiJ+VDwvR/KtHcKm4kCPhJdiCnfNUkKVPr4OAbJCkTIWrMHjQxRmM2Pv
UjxBqCz/9LFt3vp9GFrz+DwSm2ETm8tvKu4Ep8iRdYw46WPZTKZMOZsIGKXxtq3T
KAA4wCAat4K9DLcc7Xbb51Fx+eTKWca6bzxH9GEnmxDptYugXR7FnqUZyFQ/GBur
eY8W6l2iAiY/gN+dTTFaHC0VMAA4ZpWVBQntaIcjhLRfW70buMozvm76e3Huc4t6
HlpfJODySNdiGnaTlo+Ik8HVMU3DRCfOGMA3/6RikcamDUd8kbT173K3CGZA86S4
XSWg/KYn/10y9kn86OoIC9Mm5MXJc0LkyTd3qxePOUxuWyfpvg3Wqoz8IyXiVMyt
MC5XdGjA+helxHaN2eHHTArDxslzfIqyk3hPrsi1wOmCEJyVHRM8YjZW+TqosfAZ
lJsnqUPOk8NTegkODJ5qZkmnyAZTI4zv1rYy1izBLkGSguLFIB1pyV1rpZSwmMIb
DkH+hZlNQUzb2gJCbbNmFnioznFTH0u9DJeSPZzNNj32BAjHSyv4ZwnnzuDaeqYC
6ZMYdUzyoDSVcYShVFg9sV45spUlNm+nqVphZSSIPwrrYAbOzPu85UCjY332JN7d
OToP/HntmGRQq0rypTyhg6fxNJxBMKPSvSI9M8vUxSsTf8bCxBIbiI5nGiU9OsPy
Sdt6rcwCv6TMyOs6x/9l+wKbhV3EgneAGymfCNn5A9yiUGShaP9qNbKSU/5+VZyo
qVOKw5FxrloPxpk1bc6jOtyn+Ac5DErJ6FPf6We5nj1zQw8dUE7Kh3SJoSZ4XXD8
XOW1haOLnUwOQXFV5A6n6PYsply8r9YDjQ44PK1zHFD7GHOSoYISevz5pKeRWig8
Au2pd9JQz+hz4bYbCC1OEefk7WWLErsEhmmTdr3cq2I2jLdidP/2EfBFA8YjR5tC
Mc108YnCPWBrancizG3KgsuqGwYXSkBWX23VW3/fqGwEaFso3t1Akz7HZ7zHJZkB
cbb/PFOUPW16fiUYqDtf87IBM1REdj+caLowz+J16Fi4z3tsQQzVeRWTMQNh5l/d
qIQ2KclePO1TsLOaxNp3bXdYYhIqZTYrrB2bpNHE3UB1/qwUPRICQGE1gRXAQ92n
EGWmZieUQF8OgghiBqUNAuprFWXDGLkA44oc2+ImnHMntGTpYIc2I+bR/quzI/xe
5aLLXMDr5oEjgG1kjurAZmVHUFQUcQ3ivQKq30LWhI5+FwSLfolAc234Pjxytzlh
KAI0Jsbcl7McxhpxqyIO/HjiVI/lN89HmDwV5jOkE5/+9V3DcSb0/sWAQ0W3JDHj
rSFWhVXJdpq9E7o1uv56JXzPiUIjxGZCmm8b1z9xbVmTecv7t6u6c14XnfjM6tgl
TU4pDa7kqbcOXvI+6xBEZSI5MKZj9SLa6hdPi2WOyHAHSoHXskVJEFoB2aNFlC7q
rtYbOd8H2WEWkS79b/X52QnosoEcVYOs5k6oxDdB6JSgGraZHtz8eSwSWy2TKwvc
Yx26aNuUrk6qe+IeGQkhMBo+agIEqEaIIH2qqPS7bjp0oJysZTXeOL6oDtVmqJKn
R5EgWwpa8VADZ65qxmDCircEUyhD1azMKszhFHtMZSR3vM1zBeQBDDbIyC2FxT21
N4gds2DceNN9kK3vtK0J4foqDQ95AmnUbR8lNbJdh6GhN7dCBGm/QT6jDG0ZgrPp
V8ivDpLmxfxv0XaXVx0Lbqr/GMpleAQ2C4oq5DoU+GLUSQpQlOly+3gjoULjrmf6
lNsSdzuwKXO7NLPnd3nzdTYtuJWuW1Qs2yB3B+W3BOBIMzR37nDuOCHeknQMNpW5
885IWe2uVkhTC+j18TQ9YqTAvDdWq1Obap4z98Pm1uKswyrx7yK6G5IHF5v13VGK
4zbjLQTlt+NMiXrHp26iFrMxzfU7IcgR5EmBOmd1jzI96ZPh0goHmGQPpAjs7tYV
qAFF4TvqOVvlVdjO3HAMdRjSliVTvqOTBhDAGuShV0Z6/QMHXB1J7m1X9IJOG3uU
hTPykqAWAB3q6YQ6h1skwvnVHTSopCktiD8kATqn/2PyzFpskuaChjzErz8Fk5hl
F3fbsQ8E1lHnegsnBuDRukHawVbpXUf/j6HYC8Tbfwka1IbaKv21gTGHn3VxL33d
AAOE5dNKAPKYLHCitEHfLsdaTAUugCRYhqY6e6dRmYsIXrS2yUxI/YxIDow4TNSt
d0QQcKiSOiq6BuaiVz1hkrrCgcvsvgsl3qonKKaSsKrX4ohqA7queIhgXextRKvd
6Rg3fpSNkrS031kuwjO4NbT71gcM21+b+eOXAg/WASqTwwnn1ha7+lWrQD55SmAg
MN+sVvAYk6tdkkz22hI6fZE+tS+K/LSgitLgVb3WoVZGeyM1ZSF3M/z0eg84YF71
FgGI/5Mbkp3cVYiKWsYgcLizo0R46OCU1sf0x+LiTAfmJlVXaRSeRmk/5VElLuni
Fz9Mg/UWXUxDTHXPmryqkAgiRrMtKSMK32teSIpuScc6e2vecFSgigQRhrOhO7NG
/N5CCE8giZ9/38vnZPOr2fF5fRB9LkvIbTtVlgW3USvwcO0xRW/YePCDgTB1vEMX
EXNihZKzofL92optVqyKXB0nfT/+JCNrpFIZC2JGQuWNWK4u1thVnJa9gSxnwiS6
3qy+/0ejEb97h0QXnTW/YfqTZqbqWOS9ZiQ4nWGQYzJQ8cEY7HVYKm2A78vxE+qR
e3bXFUvPlE1D8lsg7KEhExTLL3XKcIgVlUjC1jGxyE1/njfIdKrr9QUZmAeadt1O
NbfnAFnSqUadNhJiY7ptbZiuFYpdu3s/yPJJBbTx4QkWC/sumA44Km4NpMu/fcwg
ktTzs8Z/nESafEsCAwqiE9HR95qQw8pns7pZGrdXzqodBJR8IzbmgPrRMs+VPUPP
lUmL5SGMNt52R23z3VprkXjAFXmP8l9hU69fi2WEu2W7H02Lkei6RXnbj/BrZKMo
J3Yxh3GJSx7RW28ONpwf9UOOzHNtD0QfjmXRy3eqcLKK5ZD8tL7FoDecXMrJbGg8
Fb3pSXwTdK4wwmVLnAy7I9308WAJDIwTf1EsM/6F4zWPcNcAoK5vmG5sb7y20SMF
H4eSV48Jd13Rnn1/oUmW2NzWGy4CPjmckxXSXzI4rTqwVEiBBF0S/KecMF0D7lCA
7uHQTxDiAHBd3o/93cfwwsD2ORkZtfjcRLrX0OgAX6N098CMTo+rx2t8sm+oB+C+
VGu1wpCs86wugdUm0WHwvFdgwDjWCF4UeiRwlffXaZvALW9J1eUtJLzIUyNIIt4p
SDzd6y8Fx+DORkj8cqR0N14W7ZlOj/88mMkPyjL9emrLihw//k21RDPaTsVNssoU
8kgEP8IeKFYdflRgpyQbD3Dz7lbx8h3+FQmbPK/MZLb2zS01aKv98NQwPSYjImm+
FHHol7LsweZysFLzPNbV0bUVisjw/Y50a0bcM6jNdVTDLjxTWg/UlYCcBWazsao+
yk8+28UJ/OnPetyoGFtRKQVOLoswvmcrCJtq+ymqhxO+XY2q7Xw51Tl0DvY5ScYU
8inY/GSri99ptjl/d7hEf2bk9zsg5WfdxEqJnVSqWi1zolrSdH5lhfYk+PTd2eG2
mZytBUFtTXI9AWI1m5T1szF3HLpxLerlgBzsh0VVMAr3G4Tb6DK92OZKlKnUAKAg
hsatkaI2kvXaSYV4t3q9CKlHTsqz6xs7nmAr/NrtQbR/UYK44AsEo2XI4JuN96x7
qIGkRZBbPjLePibRWi5LI5Q8A3ff20pWc6qPi0u5DIsyT2xD/QzmyZi2fDj8kHRJ
T1W2t0HhstGVtAc1wCApuyj236irJf23io5UwVcaazPISMZ/Y7B8qfSiSpNXbMhU
jtiUmmV6GGgLJakYkF1gBC5CNIBCWvTGWyTN/fxlm6ei4USQAj5VLhs5/74Sgnp9
ySnuqrZPlJb9J447rgFE6/QQ7y5UdqLcZQLOdR0lXc0crDlvvnulHj+tOqtuBAPx
GEmTXin6vyeWVSzVQJMYlZq4cmwWidVJ5a0sT/nyAg99ueUE4SbCYNe3NPeX3Bzd
Kryh0KN7PhXu7oUP0kRq9NgEYH983lJDsS646vkwztJxqvqKJS47Cms8E9Z7/QK1
7V/tE3C1ReC/7LbzTQ0Ut6Ssrtz0HWcwCBfzGoVPcv18OUamYBS8mznG//kXcRFE
VYhxL4L3GFPyz2sl1QobVeGpFEe8dvD1VRZTkUcL7g+r9X3UzP3eh23AQeSj3uog
3NGGCGfxncSJgKsSBNg43u/FkwW4tQBALZUnXhBBkN8JeXBixHe12njGI9Hxr1M7
4BG8O/sEjc5snRyKDo5n889AM8xvGNag3/ultDuVpKeEbA+RMjiGmzbRggAjnUmU
b3tVPvmdGch1xyJ6L/I9yYsht02742/xKgvglaLV6iuW7UiotDjdTkz63GC4Wo8Y
H/BLqMXiOfuz2So0Ng/IcChBDYfsS4yxqEPGLcB5WhZTnLD7P8IASNH1iB6PeFJp
C4ow2B9vDED/oZcao+KyqCP9P6XLhuwYAIcXPCNESsr6LofZfn4wC4ogpLzU5I7i
vx/6iVmklmqf8m9abAjPUOhvfkmInJwCZ4vN2F3zhHV4LnfqPLwY184bLcasQUGk
u7syyJySsOPhEwft/+nKt2HNK2SfShrCU8+0R1Dh93lc0rfZYYPFCm2Fd0FdGDVM
ztnNtE0SpC2C0VxgEw07i7avmhauOjZCTZ/kH7Gu1Y0BkEylaj33l6LhayvVzjLU
fj4+T9AiLDbXqeaH/8r0aDPYLkqwWp896AojxlcZwlHes7rx8S6jvQc2sHKeUOxy
ZKXBfz2h0whkDpfpD00cWqSLrFqNedG1UFKZCIPeM63XdONFRSuzvMlT8cGEk8Vg
apMqoEkcwzVS73q6F3+SZYryaSD234amDBXjmlkIT3+PbE6iCGPLIJdmumtAwrhd
mUwskEuYT07UhS+CfoU/BYeJ+NeH6AjH8zIr1ijRS/uCAGMqcqDK5jfLMs33mHF/
zrtQ/WoLdQiHisEZNe3Dv9mFAaIskWsbqauj5nGCBH82DOoQeH6tHY20wFE6ltFD
BCuN2fvfDYAgCAz0VBNUo4fGNtPDt5h4kq5o9LSDDUrjNs+p3rFjO37XgbNnePKs
6sv34VKgcfZReXdY4LRAtjVjs2jOP517ihdanhiDnbeyaQ4ftX1OnqEbeqOBYpey
idm5yV6updLgw6VY+3teZsHay/qGr/hy5HvqUgJh2OL+WOcRK/KnkWHzqU9BwNrH
S27UHXP2qPQ4G/yqs4udWczF/jrfvkIIjvPfWpVIjQMm+dIvhG5DfDK90PeaoL8J
l8qEjNW4gEAn1J/PNOV9yddI7GlYyf5iv5iZeXuPqTeP8EsKq+mGKb74h7Xc+1Al
BoWr2LiYeO/ZsjB/t9L3MFI081y30RKrrbMeXIC5AJ1dI7zAG0GA2mdUoiOhZxtT
iNiNnIR1QPj7Edy8XfcR7lZ93wOK+5KwxXBXW4HqVtvjw/6NKpOFsTHEsffTW71z
sC08umHkZPbpUvGhkFiYDl09R2Ss86NsrHP1Mm1DC8Nnt6wNakcpurOhCiybKG0o
bSfNXOJHXxiC11w5c2F4B4aDALQWgcqzVYLJRMEHUhpIKeyflmGZVzYX9KmNIZzS
SeH5gdQ6edk9MvXKD/fzyM/ugtk+qWUHO5a2Q6bNQNRigUd4ekQYI+TaU+04Q3M0
21pT/6/RqojhcS5hLI5odH1q31syCAIC6YpmXg4volxNaPegvf0zchAJFnX/DFOp
5R2Jw3PlN1Pr6e6/AjhIoHc/Idk01BnhxVrwVuxFJ+B6cFejXZqi3Q/LGXt6vRqi
AUGrPuTDT/fK30MrZnx7RK/Fb2ne8GPfy0Gw7x5NGY60sUgbWeZHNbDWLqEVA6ar
kmdGSuZuqozx5chpsvaIvLWHm1IGzJfPLdVtB7MmiQDuEOX4puQU7id6CLeYac8R
HpbifjP/PhXTMZeDB/FIhuuPwKFsaMbBfnje70MCYvXI41fRvLFBzCBjW4ps9C4Y
XKV6FzfGeeZN7ZkC8wIGgOvpN1ti2pm0sZQDWPdYW5lD7xTjSEKCdXXfGVEijino
Z1kxlevFY9ijxsaLD0PkLnGIOYyKEBpYL0P9tfMBdLCiyp91jS/2qBDGFqRvoMI8
tGumivhEqBYc7SspttY8MUWwVGrP/gKjCSmoXk/4xIwCODlDCfbutdLfIjRET47e
0eTHuCQ2FbW0BNQjHoOkbSrF8LmEXGLVFD6bltCHoksInh9LeLMTCLSGuouoyF/7
gKqUS+FpmiGtGHQ7Y3y7psQxzhVzzTS+jOZ3/NIPVkvwY3wptftSUbgaWnxAr/g+
5bhRfmamm+cKnNrfc72opF6MJyn1Lx3Miip30KpnHR2QGVDSz4VXGZGivXJ+tLH8
+/h6zezM8v1ff6OVwWoFzW517BRBzAJJpAdx2rwRdl7GPBc0O9jooTlnw0dqwRhP
Pqk0SdIrj+yBe1of2Da0Xfv/6Ah61F/qngPJxPBy5g/NTAgs/fQ2xN9qE7+v5XDb
A/bJsyH+y+HIO5djUNTdbHNWjnpTFcF+psCBh/AQBZbN3e5uBifOBnP6lWkgkCR6
C0V8RCIYf5jIREnP5e2wVj6nIMQLUYsii/3S0RCasKKi/+Rx8e7cECZKvR196ay3
fUhgKpX8qpjNNegn+bTbzNfu7u0o0uxtTR04YLNes2tSxTlLbIfE5hDOlxxldaOD
fszRejrHhBFsxushuOwZe3+C4cJthPYX5wz34g7tyaFpSOVo9Cs0nXncXWZK8LZ+
XGApYSbQjoOo58wY1WRzW8py/LZ3pX/8ktOZvFXJPzIxrMd91FdsN6iyrwUA4JLf
KHMuqHasnAJjTpCpbGak870nFt/sh9JRVAwdA8euPehkQ6cqiScWdsnsD4FEwtzR
3GpVZ1fuLRU117XWUwQ1o8GOIMurepldfyv2J0aNqebNSCDMr4HZ2op4KODeuhV9
v7MPswwyGApXFq9X9sziBUUefQNeCPhvuSDdjSn05K8leBQ2XRBw6mCVTaUVRiG5
43VYoBTA0YwIUFxslybdidC7C8GbYs34KLbdWD3GcuHaIy5RedQv/0WD06oOLdrQ
iOp1G6xSDWAb6DkLp7OR2rMLV9UVlyos88dhR9DjMXpbYgMI+Whw9qDc8i0k/b06
HSCg3OHb4ZQRfTDZ5ocyeinfOgF3juCvWgYXW5X9L+tho1PAxF8ni5WlQXYCJHrm
LxenVP5l1sfZYh0XX3XtbZlx//WszAhi7NQhjjLyfCHDqQLVmlgi2KG6CMVNFZfB
T2tTTpOKxyi4hRiPcvHL4e4wJF/YZMO7xpn2XpypVTqf9QfzuKvMTTzHJ3cwIry0
VGkyLr3ABJ2Nd5NqzB2fxN54pJBIc2ERWuJTcAzH9AvYzHqI7cgS8TPsDddU2Ug7
ZZuWXigpZdEtxWTkFSQBVkgGJSLCP5cqax95QcnoifWLkHeVB8fukODQFTevUt3R
w3l3bUkXeT4DyLyEXysvlJVi7MrZ0oJlny+3jDmYIc5w6gKdnhPJP/5kckQ+M2dw
BvKQRYtfMLDptFoEBAUir6jW4lFr7giz2Cp4ewBbqVfbrnrimefcQBPqq0CIa6OA
NZnclWDrJQedt0yNbtUe6fpejpPXk1JdIHKlPptSWOCEpALxtFHxTDsOc9y0YOR3
eb+s2PtdTt9lE7vb4t10tnRr3wd9lJqfITcMYTLfalCv+bJ/V/yJgALwaNRTVWRd
72EK3CpD9RQ7dLT87z2147fhso4BwEJRMjYsCYbFKkcLVCtOazLZNN6fqUJaKYbk
dfpIO+hjxUXkcTxWjuuZshybjbvnGFQTB2JZKiXfgDynLGQeqTbEWuwW9m/6fZQF
N5mbIJIA5ld3ofEUCQajjIxvHwMvwM9HbE+tih6Y6gltaCSNGnsqXCUHXB6uTPWc
rL4HyJy1LLtcCkMAEKsvSn4Nat80OG6NEDSTlS4Gzw1rO9QdAp6bw5UX0lD5plsw
pACS+6r98Xlz+aOWoG+/NQsfLAG5TLWcIPCIGJgFFRY=
`protect END_PROTECTED
