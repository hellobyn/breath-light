`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FbEAc0mhZTKeUVfh8zB+EitVfjMVFAudIS2g609lfXr3x6Rv/T5e7TuiWlMbrU5
8hov2wHtO+iOz7KS8L0CGppcK4zuseQYaLNypy1vFeLCY3A2TTxuyLISA7JHTX+f
sQPrE6e66bJRx3gyOdQ+Tb4duO3WachY8eqrBvmJoGbADGygBOkPLp1UDPE25LbB
BGvMrCPZL2Q4o4lpgmCl/uSUTZ/3JM7bz9Vh5SXiMpk76gnPKhLZ+zm7hVsauKtX
O+gDUflv4yEs6JM3+nV8nIiW9uPWVbefvHofELJKn34eYaVAlTvBzZNOUsWIwP2b
RqncjbF9cX/bqGS7w800iULcCpTUGeLRDNZQqkOJTNfrCDQZh9f4qyZGgOmIz6OY
tEjvUtD6wvF9SkGhdQBqsFSwQ3UlMJC3TFFbpFrLSb2n5YeoJ8UdF8NfYoXKW8ic
zdoo+q1JBMMGe3exRpLUqDT4AtnY3TQTXmCwBqjcKggDMzq2GnYsSql209DTh5WZ
jVYtwFS3mayrXYY/lXeho+/rU5CjYouLZc+DC0opUZyasuZNLxB8mmm2OLfBLsXu
bQGDxy1ZXAeMhnKMt4Q0Opmd1PREbk2/7rfrwF8aUohdXGo9JqCm/eSrbEmHfTLy
p5TYD1cCLcvZtQlgK81aN0AwwgUn50mSPMXQrzBorKvnTHiiSaVryYy9fyuyNcqP
YE72ksvkvA7wZsB9k3R5c2sMmnte8fJfTqPgzDvYzNG+Ia/4YOsLot3T2eis/t5F
ieSB9PaG1OAXnbyp7BPIYU09+dwEfDUXDyTYLcG/ppU1kAGxUdQ6Zmw+v7a3+qNq
/8TJ8GXV+1UasyXPPxPHgTdHtKPKW5ECiFHY4dAaJziuvfgLLmvzPjvQj/OQiuqJ
5XribOVKa9UmMJpWw1Rl82RyI/dYbBL0EOwcWwRmiR3BaOrDVEhLiWcB6nPElnY3
T2PHv/R2lGUmcOteEYQSbWYKKhv5Qxdy9UMjPZigS/24EUBMc/gUPV3oLOjXvzHp
A7r6R2dnXl2JAyQVYreSkOCDRsDPDTcU6wZerdOMFJ9wF93fdsxgn2fTM8u/kbhf
trMIS2Rzf/h7OL2WH6ish+657sWEKStvTWgBy8u0lsQ=
`protect END_PROTECTED
