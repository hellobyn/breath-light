`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VKtVnj7+EzhM/C5c5+bulND2JrJwHm1Cbx1iXt74RjeIze+0xubaWA7m/RrWs+Ov
WxEVNo2/axgAVdkDbLYxo/GDiJaLQIfoCAtvp87N9EEmnAzh44hdltL94sNte0U9
MWQR9lRWgAOjqHaU85wHKUYv0U74bgnJIP12P8JgObCaVJl5Ydq6lAZTzaqJvu98
dPY7hdvGGHEGyUiKFes+I2YYkGDb+bQ0KsoYP7r2+pkUqtQJ+x8MBrAZNdbLecz4
pEECEFYGxAPxo2z8LrWHXZgw4AII882We0gLvTkdx4epI2v3LAEJsubmjcEQmZ81
l4ZB+IWrsR96unswtVWlAccjiTo9M+UHfT321XDeiexvOS3WMcomk+XOsHz0OIoM
thegSRYO34WXK5oGm1dzKmLJcyxLWjQ+mivZIMCShrbvFePIhWTcyOONKDGq6F+Q
p8u1NlQZciHRx3uuStqGQtqxcZSLs6WsapWHW8OxwAp2GnuyDQLR7kByxn7D1Pfc
6ksooBI3QwS6tvK+TwmklkKF39mV/rBpk0gJaZW5rr82KeMJR18fO+WF55C0eEQq
Xa1Zy85slaPkOpht3SJH6lhwnUw/AgbWeSP5HuJafoK2bjd/bVTWFMPjGpC+vdyJ
RB39jAonABpBZN186edlfeKzsHi22e595LFjMvRtmhsFsgreumm55cT2ZP/ZVyrB
JKuZVmKa68u8rcsrLzUr+ZgOmbu7N2Smh7IKDGjFhrs6rilo5rmOXLm/8YpeswZI
MfnzclFg71j3KcXPqQ3GwZQR/f1b3ClLnEk9xO8CbRylJ6huJQMfQ15HGj0tVKcf
CoztWPGtJGzWuLq/vcGXF9psHOq/REckf/pvqI4bYeuv8FxvFs3T8Wj1ebvfKbWe
1WpiTVLJfV/+DymeXKLbUIOAgFear19xbF1HURd2GYp+7t10zzIsjLQfHJoCoCMF
wh0ubDu2HShPV93UdA3IvduFuvC3LftJ1nXoQ9w0+kpPMZiW9M2oiYkO6QyWBH73
CAPjrRpQCViqDk749+9u+uwlArq+hw05BqVnNV7MliIk46ki9epP6Vr9tFR8r5oA
vcg0ovnVESRL1FixJwumaDRPHWJHqeZ/WP2T3ByJciE+q2/b8lAvEtePxAU2ceo3
JTp9ovm114u1TfS+mRDJE/zCNDhrB9bSNnGSfR5vA7hxL4rOdiGb0xATZ2CRNbjU
OdyqVWigu8J+7AfjTu9R7hJi2Zh6FrD4roPUc+YaJGJUUZb4jflfIND2qf/iIX7C
E/yQBLx7lAEuYG1uJbMN2OfLy6gI0lx3BgdzUQdl6VmG/o7YR0xY15pSOES7Xgr3
OaomYl00hpRvxWFu3v2Bt7EVQE4dDTi6Jy1ydvltU7LfHWcL0jhtyGHFv3nCcsa/
ugTSXf1UQ5fw0rogHZ6DAF6Dq3usLDLTEVCiFfLyhDaV1EKYIKCIFQwbhsDXb7Pe
eUw2Sul/ncd2DeiI8sfs5Ev3LQHkHNiVXM9zfrHbFRKieqACjMaS60HL3s8I9/MZ
F6WT28AMEfxsRR6s43TayIweHNBNCiocOmbGyyHYLoX5z6gReL4vEaJUaKjxxBI3
E5hpH5FnKtTBWVO9tgiekhOzRa5yCo9eJxDMPOziPIJ/bzMC5iOY9Un192W/5Nv8
1OeHVXoqgGlWcLJTjTWaXq9axOhDpARKiT5dRsDXX7dQCWhfigb+lHa1lI130eUY
mXOVNgPYrE3DaH6yhvSOInU7VeX3ri7O40oqA9VsBBuv6RtRcT+oDlAsJwp0y9Gq
wF3CrCTEHju1aZJjd+CPuvXXhEleMRl9f9Tax5zaWH4nJyj9UFTQFHD73wpNQtca
yykrruE2UG2QmU/56JVas2GdDYpM1FpfrFJMzmDbWpxzPA4w5MGIwsU4tJYMwU+O
xfsOLfdJHcfcvKyTgCLMgMei8RPsnuRCBxj3a0L8G3/TlnKQ2EMTPAsq/BA/WNdB
inxmADUtIaW9SKzfDlt/mS7nSIzqauLr60cmiejv2x0OBOcoGw2BrRrWnqyAYjZf
AZVNQMCrfKQ+4TtQQBG9w8znRcvMSOBS5RuXiU+0OeSo5u05ZZbwcl390XgfI9fn
5xBm0v6RP00Wx6XiQg/X9SiFl2tTtL1Fptm82EjMYSgum4Y5eQF1OsYr1QwdZPns
cJHlNLe8gKaYhUcns906Vy5kk069Ws56Tu7qrTDWdlJhlBKW5euHp7WF1465TEak
4xFY3WdVLBWVh9uNK8Z7tbiBBxT3sId3UWseLGJHPtWs3OACNxHDMTVZnrQYArSv
rZ15VkAwVAfnxN21vGP2JkKysDsQ3DtWEh709CLb+HUtXuYh58ZlceKaePdnGegV
eZ5vdtGYbjMV4qQ8wRJSdI4IU7kn1JylA1vsRnBnyl+Lbr3fK9wrJNTXNJ1NARJl
qsEBkoF2EvIKdkCXyJHDg/ckJX61C2kLR/JTQYvKGQtxLehpkQzX5YMRiv9yDKTL
ndhVm7+ULhdr+hUNGpaf2d9zuYMD1bIkPAa34oyqyYb5lndJNsHSuTA9ZK2xV2AR
HBrimJhO4EDaiApyow+7pJIGhWgQej5wZhhudd6oGPzS/wsBDWMU3XIXBqE0YTOo
O2UeR9Kbs4XxWlKL5Mt9qqIKF/5F3WD2RIk0TBWcHwHR07BfcXgPXSdgP61YpHnK
zuG4knoJMgTm88h1uyJE3Ue5HDjO/yogrxGM7WarUbAyh8sPn0nihH9f9rJ8yKkX
wz6u0jrrkTXbIKR311kILwQCyuJF+tM2otV/Nh1ytUHhVc5TPp8yL1CKlJmvOK3H
TBm2tB99Dzqsq52Riqz5lyEu1hkKtPWZsxj512xcINsGKszroV2kvEA9GSb9oiHF
HyhGozH0ibKbrd9uNvpphsAzQj9XAkTZQBtYByuHXQzJX06DNpWRtTPKQGa9Eos9
dwnhJK5AT35lrLOLKuEEMHIJ4cxsnanP54Zz3kPWqLEYx6lWGCWp1ATzDUMP6109
P+hbJh3ie8AIV/z9svFNDkIG0wdfCx2+gmXmVwitmhTWhfqRZVSWEd2kzqwV66Pn
nqRXH4J/RCOHOOOkcq166g==
`protect END_PROTECTED
