`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dH44mz5RmzfZ7gFyY/jitNjbp57XPnaWfCfgdJL+XTKB7YNM8GaeS1TyK5b7mOWD
nUfLmTkRt6wgmAVXsf4sSvkJU629hLi6M9UP5b4NbdNpTapIf9tj0bPvQiTUN+G1
sn+Y2wXH/3Uo3mERC3iTOsc8i5cGpX00hwM0xNEJTqEJ32hSgVfIp6xpj3vq+t9F
91ReCU4qU7lyub4et5tO4VQexqNH6Z/E/zpa1+CrNcFIWnn8KvrGd7PAkD9dj9yI
TyMjSBs9z3fifv6fGwsNY6UHN858GPlx/Z30x/JxsoMJHTAWNjToBnJf4QMeoEyl
6OnMNo9M7zpovE+TC3592NADHYV9dxT9LrYvrBVmVANetRgZHxZQeFRVRkgylba8
6T9nuG2gimK0zsq7RnQuUK8bIZRgW+puIdp2oRIqR/He/XOSTY0tZH7hUl8fpv9L
H7/sVE9NqI7zCBMnxfzw2A7CFZtNUIOYCn/gqe/68TuV389WLrG5tr9U8KAMFWFV
adRNwkv5WuCEP8i8uJSW4NmGaBWIe+IP4ru1CoejkWAKlPUr8BZRTzKGsnVmWW2k
t/Gzgwqy7owX+IwNe92dRFeuvlwPNaVEvQL7BSIs41PsW+8ra3Qqh1LuEluXaA+V
2oVadi3Hn+YUqOZ9ax0pGX+b4Oxctj5Lc3TMkTT1kl0KTtjrA35a4OcMF73AShPf
h4433ehtHMT5p9qH+nhnSsFpmrwT9Kb5cd5ZlW86m+rJ+ACSfqQ6U/YdPtm7OpwH
XNju8uvJmUCWE+3/OUGUyU4uX2KmpkOgMb3XsE2IwgGXzzHrYiMp2ucnPhgWsZKW
xpIp+z06jE+HjDu3i81WqERIaOSe60VwDdh5zB9gVLeQOKIX9CXOOeN44Xh2gvw6
n0VUUHow8R0jhvviNtvdDjaVFiXf1FIYYQW6TzZnOpxkHYv6/R8md53Ftdh+mYGv
2Ed2KQwxt1CPpMMv02jsvyLv4KjGqJnWatOSuNkuIRTpjT+/pTHAiY1N+eaTowx8
FvfrZRFG5kUP3DYNVsc5Cq9lfMXCk5aLXA7BeJBwU6LazKKzKjTwCZ9KOE/5tAzQ
PUTz/Qwm2HuslTF4QzaGfxhLreLzSe6BsuMGRETlvRAvTgfK23tvklvxQRQkn1cH
ztmiMaSh1cs7pkZ+auFrWsrPjbDE+LAuK8cYFNY8JvzHBwo3w1agAhZt4S/zaV5C
VG1fT+M9qcPqh5JrsxJZ1a6wDyV1/qP3ZOACHahV1vmfXjHJzyasXcb+maIqMclY
si3Pa41xVyKOE1/D+HeNNX8AI39be9OeoMBujCDFLzWRCz4p5WsWVq90xLCJxedi
Fvu15mOurpsxRXTSGgIrAHvnbKHECcgwNEjAlRi9kD5kD+TKVexCcnkSvuo4y4Vc
op/iIGrOox1lpLrrNnXm57h0A6g4HbCbmswjByOozUNmp2aBbuUrtNdu6Cg1iAND
08gVdyFUwjdBIp9Lcg3984smTUVI82aIaVyO0wr5pBiYw96/+ikARh+MEQLjXGUt
XVmeu8PtHVRi6Ugk8AIij9lkO83ZMo9IoQ4ws91lXnnH/5YLWdgDnrTm3whBEHkt
ocGw073Xy/sNwvRF1JhQJ1V9Ia1hIcksbpGBwRWwSgBGtkwKc2pd3bYk7g360XSA
emfX2HYvm39UXurkipbtzw55r9O6UVUel5BQMwF2WGw8z35fIPdsJRibfig8H9V9
H5jySEHvcH5yN+mDDbNCkxmaVGtnQGeYG4aM8pZ/N09WdloTtv6BR/4wcw6GS35X
pPrMdDOdAqcKc2Zk7FOqO/jQepy0gy4cXqV9b9/6sYyfP8XWZRx1ciEFYIE7XJvm
y7OW05V5QOBw0oZcCmwv5FrzFjyjv/PleczKmXeyQQdq9rV3i1jUlE0Abn5MWPTt
Xe0FOxPVrgGZ980srLTIp3Ab5Wex/nwhCT66fIQqTv6eLoUZvBoeHryDGlY+fT0s
oqyo0oVMTDPGgjM3EL9ySmnhlBGdj/mh0PiCPzVTWrbP28pcuPie6IhDlv9OLmHF
QxbxueVOO20HfqwBmiRfN4SpoKPuEv76afM319cPoSt4cYq6566htZ7RHImjoq5D
2stt4Ey9zAKrxnzDRZ4PI3gUZFn1CIbO/pcRDYC9U36lOYMP9g0aUOWFOxaI4CZh
Y0Pb5ek5xwwNVLAntHOOFGHzFsGyTtPtaPOAYotx7B5crJPiZQSkIEaJ36C2vLGS
Ju2orCMjU2EAIYa1oC2zKNxgUmMhDr5oDmjfEnxBtz1fftzeOXzeAsXt+zIB5Csd
MypZLEoIciOWx0pdjJaQUVuSHe5d8kg02K607yMujk1rZaFJDXUKanCqlTfIU7Eg
Z03cJgSvEhZQQd75YfGRYRguqWwQfOipBzjdWGsiHJZ9HzYaIbWM4E2BdFEsGnf+
e6odG3G4MmQb0nhI3A+QSR59xug3UTk81GjDRFGwM5aJDMD7/Kbzzbo/PSpk4sg+
yuGxenhIIP5CMsvuFLrtCzzron3/shMVtyZ6OMhhmo4irUGPzq2KDn2tXCWn50Zn
ofQNVN4vpXbRK/0F+Fo2r8vj37RCHg/KZcJCxRCyA0DoxZnoqJPkaLyiap7FFKTG
9p+w8+c0bRXZe5UEtxq11Y03yWajc2PzOi6/ngfLy+ijTVjuRqVrQrUbyKgEgYHP
ic5ayZXEFnrYizW7A4mW6rgg274mkiw5VJSKffTqs7mQ4s6nBivqjV83FSKOqobf
9TWjDr77Fo4YHYLq7CHlZGky/JlRne9WUk+g6Zg6/kV7Z+/B/zf6BpT41QIRxONR
5/elubBT6/pLTehNQPm9aGjI20MgjVnd0pOkXGuwmYKe437hZJuzpUePtAI1/yy6
krVkBedEZjEkmy8TA9p6zti1qSBKNeqE6iQyVTid0jZ7WKMfklpEOY9cnXhY7Zjb
ihQAuLTM2j3ZTTc59yeVRKLBq3BH2QmDr5kwLDTrvvsc3gzg07uY4kYTPujBbFaa
2YWe7fxmr15736eDN4QQXHsJR7qof5h/cuQHymXCMXRYFLU6zpkV9IeA6rq1fqwo
yTQh59/TV8M5oe6w//iguZ/8whUpaAiy07anFs8CBavUCBWgsTeLVnegEnC+1qZk
CS5UK+KEDBr8Gq1U12+yDHP/q1QvBt9Ii4YHvqmURcq/QfqalW++mCwS/5op9C4J
PbXGljTYb2h4BdTOid/DuhBKF5BOiZbGfFvQ+v9r8Z8GK1eE+MP+X1WLdx+dK8oe
fRHomr5o6FiFnfdf/jfjcaN8DyyOFm88ECU+nCtUJy2CWZWm+4VMSAuHDqc3Pu3n
oNqzYFBP13peSYkmWKjgXXPHJ+tQIfjDKjPcBhFGiwKNjD/MFz0MumLQCbWzzO/Y
5hvi9Eh/eqXn1swiZaFPWQTm/jVNUAemCy+1gv5j+t3Y8vBz/k/5DRxEIblrKraJ
sirs8xt6Lj0KcN2q5md9JM9X6+YOiKYZwhrS9N28qWDfJmYU9rmYAQtCzcwNmxKq
BmdDtBC8FcEzzTCAuAk9FHTM1Q3UWX5Xlr+6HpP2zwe0SX/dJtubJPkelS0Wn5f6
gbe1W8yeEtTaY8iQlbOJ+2kD12vDS179qc8pxF243YFk7EzdhcfNZD88gOhw/0mM
z27BHEuH3JNrWOtlHGt1q9CFLB5C2DWL9N2fn39NPgrhUk3uW6hfgYk7hADwgsju
s/zmaJfZphKmUxQ15VrlY9EVafqi6Oa8fQNTm2kz9MvvlnWSvhUZxM9Ue13E6w/l
hE0c6BV/1oqWH+9PO+qF4FOtMCuOhUE2qAi9sc+G1VqBRLGNkkokV6Vftqjhvq4x
M+bO5ESF4myyhTPAKqiguqPbcBcty2+KgWLtU+mQ906pg9l7oNbJKvjkJ2kzRFSO
pMr756rhxa21C8H2FA07cak4aa/Jsd8rRJHeUk1vGwwA9ejXQwHVClU9hn782g7L
wu2Wxu5dfcfpVnCkf8WlCgaNbO9sEdLTW81G2Y/wchqgG1WNU9qaxxV3tazBrAdp
uGJ4r1nlYggXWRe7ec4moMixkb2Y+c9oyxx71+SyD2go8ONvIzBQReri2HR+xT51
rJoaNbkvrWFGxf3H4qNyEYFT8BosANNX9UliqukI9HYLAHoDd6EgKpl6T2qNpR4d
EfmzoRiwDUtXqcDWxik4S/h51fFsBuasuzbBd9T55gfAuupOSWQKP+ue/kLBrKb0
m3lSCv0v00mXE7OtOaDSsILqQGwcPtbRkggGfwVHMEngqzxdV4FbyEyCs7nJkS70
bDWu4QWwakvK/anwRstEVHwXbm/ZR+lGdnOZK76EQPVf775tjZCf5ghUtIpeDmbT
M3Xuke8n0TzA1Y2n4Z5tkVo+hJGFp4821RE67w4XpjITdUA1EYN6ggYptJUdcaI1
vgeZtmNlRfVbOoT4B5wjPBiU9mdK56A06BjoPRUlmgviPjFsei2bc0xD+UjpMd1Q
N7tuX+tNiycpmkwsyIVYj0/JRYGtuUb400l7oCUaAvRlsmvgkq40eRmkd0MMpdJP
BIQ9OnJoAr+2vgaQAbe15MjswWjBStvJjxRBgEAjQSvRryOkPJYulhBKOrTY0Rl2
q+/KFrWsJbECBnEyLKUFSMNOYubvJE5zrp9qWbjBxPEkd5v+xzUe+kt01RjETSnM
YC8q9VKIYNq1Sfpem0QukkX0dQPL5JzYV93xdvrejrZ3BS1gCQ7XC0qyQJ4R9SsK
pyIduvk0fCwiYxu0/Zh91QbvtSrhcJxddR/dpkkW7VAxc150QqKhfhS6R35GfcF4
uukm4jbPFKJBtaC++IVn/G9v8LS43RgChPmkrtknr3mx88eE0ii8tfhuqj/5a2yQ
/cdF8F9qQD/f/uoL3tG//y0jGHBXaTiV2/fqUZc6eKgkNVIwjekUS8jRT/uJL8Tq
Zd55xih8VHpD2Srou4tlCeQidJUojX3ndsTbF00h3rbPHedAy+AmvukRsf1jVqAW
YyyEPbJazS10YGqN+vMDxPTR1mj2x3eLnayv+nraMjh9wfzpHSeFEQ14PTfqVT4U
IJktksih0TdgYpcqs0iFJa/AVuHSVleSBD/JLCqx62K1rrGr45e53E6HiRRZfMDZ
l3mkOwbd9QiERA5qAAPtucF/KuIZVjDBos4huhaak9NcygyUU40gJZ8Rc3vGaAen
v7gQcFKW58QFy3GF9fehbZPObhKHx2eBJu75Hs45Q79urhXv1LDskNveuR36IRGA
Z27FbVAQEC11HKLBagjQXJQZ4A0SnoICd1z+HX6IO93apthXDmUGgeAcVdyAyfVK
Ud+U0699u6MJHSmNxFqlRDXdehbO0kCuZphgHMdr8kF5SC+YMT8TVFp3C+8K0OL6
MwFsAp6K7dk6V+9F/rA3aow/TGCEmWtdbnYUJbk1poAoDyfgSMBTiaOXRZnc42FB
EtbZEdO5th+zG53QdrUhUL7zohiDWHAFSzVWBw+w8NAToUfDVCcOPwsNQiAcsr1k
/zJtZE7yCt6MlscawjXvqLUUZN7yA+ar4KNSsXUC7pUXKVq5a57Cz7YTedy/mmnS
gfTjU3yXVaQtoHDctaAKkuyh5Wl+Z/BIDNtBo+II2bBVaf7IIHxOyx84IyJhIBuw
R32Ih1iKmARdqKTVprgfjJmrDokhg+juVvcr4vgqOy27s6ffuF3TWbwC7v/HcQnp
7BSDV9Pzkyr6OMgH9srJs1T/kMDne3MgKhSSYgROn5ZeJbmzx9bvGrWV9eTCnmvS
oEQDEyBJd/2LuKJMg0bSowxFyX3XVMY0W2eSyWNWgUR4Bm6cH4Jrdq7er02Efotp
iToG3fG79vrrfWCamYpuI7j8RknQGA4Wcg55P+WES+0btqOm1dWNmt+fYtVE3aKp
WDzjvDfVOq8liyCQNedkcIdMATKfuCv03QZAEyaSFQcvDWKyf6P8GCEwutcK/ShU
6DAqHxfEApLCci4sW8IcntVRzJVK8O/OkF42iS8JxvlDSHbg/yfuJpli7yCpD9GJ
FMKpz4lk+sjsss8Al0MrlC8GluhHhxVAwTW4mBoxake0EEqqa5+M0vX48MMmSYcZ
Z8pb/sN3GiFTIvDPNuQlXZK62Rt70WCCtomqXjgc47HYU6dEKt93pOPAk2K1l7tx
opiUjtTTLRj5qAk5u3h7M2Q1Ju2GF6SqBaMAK1maR9gdt560NUnq0LQySKDRV1Pe
Lt6S4ErE5Rn8Z7rBlkPzfCYhTjDzzjtgcDdIoVgwv8eg+ndxS3buBSX9Q/85XOPp
d3iSGcmyKoDdrR3bhTb4j5bRHfx1mZ1gB0WY2/aLNphSLGzn80BBcY6DaUNoBcDI
yBPoKl7zc0VZkndNWt1MWXb7z+p5NV62yGqIS9zGSDPA78VG1Jl7f35MI9WQcy7O
xiErzSj4bPYVvibwxxir4QUaYrjRb7jpJbQWr+HvVZQRO5mYwSZqgy7ypZVnLWl0
ZiV96cvPUxaSdCoE1HkHa+iYq5QeepKqt9yieJ1uXXeSXZRUtlgRgr+DbxCUPjFU
mripjIcpZxYZGaF2XXldinLJHhvrSzr1wf5NRBcGL0CB5vRVF59wFVwBsiikdZU5
+DoZKu/O5WdUMbN96wWjGcOew3WxPc1hqcUIhOvxO4nlNvD4OfOli3IJQww20L8J
590cBjccwxfCgNtdZpR5V30Gmf4ww2bH/1Euaxy8FI9bs9yGF0MOgqozE8d+rZm3
kN+C6owJSumsA/ZWFpwZFMepTEIjuAEJ3GbhO/O1epE/ZNa/oks5jvven1spJ3Qh
9HayvbC5hko/M6hVmTk7vsMBfdzn9Ml4MCAwxToimwp4Tue3vBcUxGOr7+dui/mf
zerEr+56KLfDFBH6Utr0TinOSyTbNTrOFxzglZX2yxbe5VI9Reqfn3ePHGdDyP0J
7XXbNoCcbzqtem5XXikZRXosl49ycHwuBs9HB/J/fWGaLECvlp4yhDH+GCiIcDk1
ItOJ0V8vEVjpMlXkIrvA4LsaVISGTlCmAKSlsA0LLEVxKjujoi8G8qAcPw2kAQCp
TRksCAIPxxpc5qXPPpmROwa2vNz+v2Q7s7ksY/la6BHdNjRyt8ay8R8mwV8wLX4z
AJNnzCB9tnBRZvEOLD19iJhcLen+1dziVzm33TkXdDyWufzs/CgtPR3fP2M8wVL/
sfNk2BT5ZmwnoHLbilIrZ64dLAS0OsnMOxnZAJ4RuE/jupmFIJ86jqH5DSV5q+5t
WEilyj2c7KSQIlIH7BqD370yOwMQgNYqmFCFffxvSmFLxI8nvHA6/SbCzGqmX+QC
iiITqvniT3rmN4b+BJsEOKcHKP+RC4SsTH6bk9myrmr2IyH0K2p21raBnY29S5B/
gJ2tfJ9oGVS2bvKgx5QRxU/f29LezWxRPwHPl66CRvzq7q8lwPIDrz6pGFz1fDCx
TI16gerqwqqs8Fgj1jiRl1szMKKZV1Vec83KrltLTgy67OipaMtWrsiA/gsX258Q
ci/HY7gz0GDztEyitZfSTdrdugo6BinJPrx/KqD3xFm20wCrBg8KDcebSnt9aCk0
rZscnH6Z7Y/u37Spm/CQVB1jEH32usQVe3IFLfLuQfPyTcTGWnYc8PpIfOUbTIcC
Gr4z9SqL4yomGvxPeCftTqUqjDdgX0GKzvdML6o1a5pva4BjYpcPYgQwBl1BAoL9
g9QKa9g+RhsQv/rU/MvBA4ZHCY/UjJQiquWoLmcQT03iIK1Wx13bMMNh80itIvoy
6Arv4z9Frt2dqb/LvP5vE+gsqqM/le0A0qTe+cTD9kL4ctuay1dvYnZj+CgtDx/V
ZiJ/nQf6HszGqvVX7dZ+xbr3+YqoUcGbDOqP/wUZAuqofjn7r8yN35Py7ygxTIFQ
VR+vfWyu0quvSu0FK9N/ZSQnJkXhE/qDgGbeMum5sCQoMdyRQn/TosRC2rJX3ZJE
qWc8TrKbfVGlP2T/fWkqJqcHrUtwfJlZT6l67A04fTg/vCsGxw6ZrXNqXUPk4QcM
VtwKlfoANJMFEHSlZNhlmfNsnhf5qTiltOEwGP01lrWBU08psouNj/piYp0ELkRi
MD9gHCU5Wzk3pccdvJQA5GnLgMafS7WiPcmDLZTPhtOnfy+1oP7hyDUPq/L4O+wR
EB1ErZIyCanSra+1jzTb0vqOuMErkB4xkIJJIGdrcEGGFrOjLT7bcvw+tUyYxDIg
q/ZmtuZBfKxKA5GJeHL/hf1Qoln4Y9JzsopfxdnUnSbW2tJSlF4DZrgIEJjMtlrE
xFmr2OuVZDB2EGiupmcrk17j/LFr5OmRBTLOY6ojwk0Go0rsKcrgdKm516sjH8/A
Y3ulzFhOCsMadCRFs3Z1kcS4N33uMjy2QWT1cBGkdKj8iW9IV6QMh8x/YpFKM4Sw
gweWqVETx16py/ez2X2JOCowHQZDi12w8IC0tKCZtqyQ7m3qPBrGehu/s3O6URnI
rvTznJcGqRET7DbZNVtesGzyqXs7l34cor4L/+8bYE4OHuhAStJvDFZIZb4m943e
/AxZHKUF8LajilnIfQhrLxTfyh7GDE0fuQCOzFfOBRPnk2Y82f3ddwVhCE/13YtU
c4nyTJ9G24HIfO9OCwuFLNReYFSVc+2chz9EebCSv50Z1NXR25s4AySwvmcHZqIL
3YyF9+7VHw1Wi3owGXSl37QoUYE67JBIRaCR1bfw9qbrYf3wbymZY7tgvUFsr/D2
ns/r8hW3wUjW0JvCUFZholv9Z0G8pM3yIKNdvK+24Rosb4m07Q0ae/7n4EXgIzgL
oj4M/vsE1ZCbzO7mRswH0rUEd2AcN9qXo6lOhpDdMleTcL2dSGXs9NDa5Sp/Wb2d
FEUuQ1QUnj95TC4Yi1+P9kYuKVQHI6Zzl0Dvlu2kZFgJKEJFgerKTyUzlhw4b1xf
HdHUBMyC88JiZZhGBbD1Tlx1u2ij7HB90BBzA/YHZ5ULdCVEU5mBlVOdOYt382lw
IEFDBtniZSKFQr6/831mqi7jaQvmeMSoPGd/64CyaXzskqPL2PGc1tf5Fo5J28P2
xZg4UcEJ+XwdLWvwxKrt4H9Npu8Lc8+fNPILFcJklkoYxuRf9pyyPijpNAGJHeZK
HahRukzyGuwjL/QBTDYo21eb8lyHVFq1X1Scgc6uf5caYMYu6JQMnwFTe2/8joT2
tJEPoylyUcax9yfxs6+bs+Y1hCRNaXssOjyLVqDLTmwWtgmBx0DmpBNeJ/2dyfRo
KK+TdJhATRbQAPy8N2MDCmQ5pSNqVGDTcUynz8lVGcwpIYAubDG30Zx0RBH7hv5d
m9oBB6+SaWiUEIsz0GLs8Rjz1C54tgxbOqea/nmWQ1MznOhaSlbrg0jdNS3ufbmz
t1qj5yTzEapyQCsTRCrZrYl3WltidugIdE+CejDqAunL6V/4lxiIBfzboij/aPku
qBf2eYyW7G4B9vTN7Fwj++v4wJCBpU5Dl39aPFGaoS9Qn8pXbStOvUDPvivDGn2Z
Mzo48LtyszLmWt/ig2AcTg==
`protect END_PROTECTED
