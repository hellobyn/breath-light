`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PB4HRyikFJOCtFtNIbpXV/D2tFPopGJkNVcP2l2LFIqs6A0xuISBYD20UUABflQD
jVXZHWWDAVJsD3uILrro5ZOHA/9cziZzC5FuTZtdSGVy/Azkusw2D3dWkXHJ2OKk
mibTvdc+MCfS63vXtsn23j3cu5C6nBo86YfkPtkQZkRwddiho7VzSrnjbwBC9PI+
nt4L6pI856BtaLInfbbTScGsar0wfF2ndtdBVRtR12DfKhe2Iy77YkUTNqXU56Y2
k61PidthPFBS3QdoI2GI5TwlIm6aP7gCRRqq0B79m/ZMkR7M0yYeFYbyfmeEzG2X
RPdZALBidM7QtsbUoK707rEor6YX3cGI70vfvvEtmlnEk0qpe3J5KznVfXWF6MIX
O3NtcTk3lFsGbYfL/QTVkEhj7H2K6x67Y5llV1ZoTp3WHgOkYRwZ51CBSpbxx02U
dqHfhK7H/XeUHZo+UghElcElQKYZWKZNZ1YDIc24VhTeARX7ADmVYLAZAPhSieUw
MedH3RLr6MB4tLmTVFz0bhBjpuucn23zbMU95ZLu7G5ScY9Y23EMyDYu4cZlbUc7
jzT35bd8wvcVErMBUrKDfNwBfuOUFPYRNCwcl/aO+rvHAnnzjqDPnSyKNwlIQdah
Yfhd93oPdWUlfOEK3PYrlr4lc37k2yfwdusH7zZtNlP4SLAPSGQ9JXCPYqtQ+qXW
GIr1mbrQmpWVdMTpff+knIeBhfqudySmY2eta25zuebOCBLuVESDgWrmUmsv7P0j
Q+zA+KZv0ybctf3ox6CzfAMuRZZGzksXywRIsKwEOH+XLlssmE7LlB+Qn5L61sD4
8wYVrumsgTS1cglWeMQe684u+DI3XVUROuAq3Rctgf+UYWsxQMsiYPiH7XlkEXAv
FvyFDgW/Z1O+vjdtqsIBx7zi6D3KZ4JLfa2567yD7oWhMd56SAQZtLwwggnNCnf6
ddTWXe1mL0OF51G+LKfwYY3xCF9MUU4KGZ3XPWYZvKJrmkD1ukzJ1kdetkduWKS+
wiqghavK9TVpyKZIAHem/x5XMtWgLKdmVZt3qwZtTYfO8czF0DV9cGx8mqsSfMIt
xmlcgaNn18EOzsxbu0gBz4EIVmMVMjiYrLce6Vu9XAnJJb1zQ4PQ+NW9Zx+9jYeR
quyuLjkI84S90SpcA0bGqaKVOxb2SkKcoPfAzTi04etJ+FVLhekWIFi38VLAe84l
LVb+AbbgSf+CiLgPQs3Y+h3zgorotAwtXyO2Gyox0Rxl1gPzrKtiP95EQN2g/rYH
0l7uU0G1YwCKuW4vZcxpYIoxs7QDLD+6uC6YT6w6Gp/Nqr6rShVR5opwP3kXR4w6
fBlUTUzhrtswHZygl5EzID+ynhz1uL7a4XJ5yoUtNskdyiMX52zCnyqPHbgdavZQ
nxg6Je01SjhSmC3IEkKpRCAkcJGh1A4fE7IyDTWvYZ34xc97NREBJVqdnGBQw0Jv
6kLYZucH7Wa4P4L7s45nwyLGdaM9sXE3jzpUHt2AdRIHc5ePitqBAJeo8N6L76Q2
TOacPzOZjnagb08RJpxE4RYewKHaMdnvzk2DimYURPS1wA+NBRqsIHsQA/l80Nzp
2eunqC28/erTqn9Kb9xZUhWwEOdM/oN0qNBBiS1M4IkfpMWJKZ0DbBvvgCBOXbG/
IZYP1XOfoPOy3d1KqsA85oSMH0WJ8tj2cuVPr6Fimc8Tq0gNekpJ+wKkm/FcSSKf
FNCePj7hwhm0Q6vMBIynmR8fZGzfj0Ckgk3waQwmR5FWE91IybFw+1y+THnQGo3w
fCQykm/k8WsHzrFsB/BoX6PMH5p/vv2hRT+XSjRb+QtMTb2bDtG4j2mueXtiUx5Z
gU5IZBTNkVAkjNoZlvODIvXVC3JLOsjOrW3WE4EsUhBBhEnhvu6ONIXu9I+pk1we
8wr8s8/y+OmlTNDq7arLnXa2a9qZlcEJFX56C5aHLucPK3wX5mtja3hn9o8+nV82
q61qVHUp/XbwnbSLsKGz8i6j895um6ewhl3+OZy9JPl+4GOqeE2lka63ddh2VnmF
g9KaK1u4Q73KCt3lbs1jNjUhIrPvuzv7tMzG16/VavH/gCqa6vV2CgcSm9ETLihG
4xiI+xWcOGrAk72DRmiHokLvBiGha8SK97W0GAysMCbZc6Zj7r7MEW1ZAB6J9g2F
PH1HnvD0VFsfWINxrB4xDOYzdcU0C8Wum+ZwzWDFPOcle7RwySp8Z8rr3Hkqf5oL
DLMm+Ru5U0yP6Fs8DYBPWc4i46lofQ59nh704qiX1lH1UMnUrHActQbfoRpzZ5Jr
DFP9deH8vHulJc/HdpkmNwsDaxV9jR0m6g5miP7RQNJ7XmQn4w0PpW4wGG8OJNMx
/YjjMeqwzOZVlV4JBHKTtre8zAlAdavr0qsTFbRWYziHOjyhDkHg2uO4PEQlbaTf
MXTHEpaPOlBJph9l19iCvEqTTnEawB123IlsnV+Q2x85iuYel17KOyVlaowwCMSL
VNpC5eZtfV/XG2W+ikRQ7ksVb+POVHePdolFTRq9W81xor0HW9D0n5st/7MErYDy
IadAMC0SdQpnUEGViDEljMp0cls7mu1E0vEER374PDUAyXNqr97lZ23iUQA+wFRp
Q1VswMNwlpfH5hnHrCedEUG4QzAgHKbLljcS7vHRjq1JPATtHgj6PdxqT2Vcnvkr
pEB6tj4MNTbQc3iYpRfg93labc6qPJubDSxBd822TYp5pfI229FsJHUN8MhbR0Ac
Nv9X4bkdtQQaJKZBSmRcFMIEZ4Y+DBa3NUySQVdm1J+TcgiLUNropqinkhH7VbCV
hX9qGtmyxny3pNeGPwplcKB92eID3DjHPcfi347nwZTkGLMFipdZncKJgUXis8Wc
LZArUDP88IVdE/t/69eBISi9i27E6UC0W8/RlG7GcCyfk8Mjs9zyBhCKCZfP+d37
ayRp7yvY3trNGxivTYbvngM6QOxnyH/JU7wR0YlY7c/rVjrLUjQRijdzoGAtTDWQ
dExWETRu4wOa6Ryv4kmXYGd7cJQRKduLFYeij3QEzVi09wsLe0gW5H9+qxMnWs5U
8JCuJVNHH6MenzrXmZ0fsKPK9np9NrQoHtMgnpsuk0dn63cMiznBMoBg/VTJ51YI
IZ+HBqVqG5srQ0Ei234Laulk4aXAtuL+UFzmXFb1Tl1Rz66c6urhZgdmDe9osi1W
9tXSHtwI0MxML9eBfdX8selY2StZZdsEVTFGzhuZl7Fx6Qp0dclpO/JlOS0TNrOj
m34CkMAc6qKkGq8P/LLj6A==
`protect END_PROTECTED
