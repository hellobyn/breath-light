`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raablJZwSd75z2wVzfBqVoWD1SRslufYVUs7fayXZCB4HE0X5QkwVxudDtNR9tnA
35ibbYoWssMYI/c06jLQiiYXQWs9YGI1x/BMdyBnDQi1IYvZRW/vUTQvi0jqo1VR
0AUoo0JvK1iAcwHhONEq0pJc+CEPtbJEb1jE0vCv1Jh0YJFALAO7NOGZesOsw2N7
aTBmlzWsOHm5cz0elOs6IShjomYNRraolegU3WPy0RDK4yAQmOm5trC6mGXGAqP0
5t4hWqZtXnCzr6+fhIZ2gp24Of6dOkKJ6TJxbjbwcKcryAukvWa4oukZbbOUQMXu
o8gPdopyChfUIkHO0vEfy6/ifrpXMKt2ycBY0IBNq9OE70RkeHbeO3dh3GoppP21
1OqaPNGfmsNLjqQzpm73Kh7j1YVl4r5BJ4oHGM7L4XCRT9oVXyFi3M5zpulPHXEw
pL35ZRtk6DN+B+BcIeaIs31bm+nfPuqlaXXJy1RpC1euCxsKaGHWkKGk+McMmSYW
7t/XNDfCXKq5lcm+Ew7qtOsIgeWszQDAjIT6VidknVd1p9F9lBNrZB5S+IXOZ++X
0MNoPb03CisZsax3wYZYLQWljWcIBYc6ycI1nYrNDLruhWu57VkB2zRyVSm4Ohec
AsDSKbDBXHXtnaVwB0gjwqY09bAaGwaLFkN1cVo1l24cmAb5WYx9Xf1YOu790FAY
cNhBwMkm9JHDWEtxnBuTyRCY7Q8Dgj9zKAnjRkREEiOQ/SAWW8acmOUUSNDcNY2w
+ei/5oYP0rKUYHlc4CcZF3BqPzBL+XV6SYhilAmf26u5jNwcOH0zibxLemx5StLC
mz+tMmEBCw/eUW2mBACLQt7kR+0dLkO3zKk7Rxpo8GfvHgACdN/IWNPsk+2BeLUA
SkipRpbRkrcbfYSLSs5TspUbwCL9zz/ssiWb4nqdUHYGHO6IMYl8b1+3uzQFi3mX
NaDT+kydDEnh2GKo5Y0wva3FDyJAjjf9yZSDoTTXlttvkbtRPdNVTZuHDMG6PF9S
En4xiYv2feqmF4WxXMN6pjCtMhkL+uXG/uOqJH7EyijKYPX7O7yadJIGgkhoDW10
11sj9cI0OSmWr9xc5iwRCW4fcs6icv5zxM/y42qhrSPNAWwJCaEnxJ2YKNpCYX4Q
x+N6IgUeM/coE2Wq1osDHY9T/XuCtdSS7mxbRQH6EKDUOcYlQ8z+0gjxE9OSvL1u
ihPRszpQLwzw3aSX8upRzu1Dj5ZHuyt2xDrbvtIpumTpJ4hbQZYZq7eazqr7GP3R
0oOhSZ/fgoMOLM8SBumm8i0V1H138fG0lRjIgv7cby6uiKipm39ubGQCfI/+1eCz
RgJ/z/Y6icegX1Tk0xYhz/Ahjy/SBJLiqs7ONU5xae+uve/wOMFcXE/Ahz7HRrJD
4FWTiLpFy0hvXByNJjKhlNI8yINiuBzgr+4slZgzpDpym6xkrieU31saGDSZ2pwF
X4Y+tHCC8zvhkDi9IdpXdA==
`protect END_PROTECTED
