`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkqlBZRNKdHkP8kqxdhpqSPcwGqIsVzjd5SMOtgBST2htly4jcMOdXSaBHwCpDtb
Gw0aiXzVHf0fWzM69eYvcWSk/IlNhFGXy/aVEPhkfeKo2E4C0NxWJ/0+JTD42k9R
XQpRiqKa/bLzwGJA/PSWmngrLszkqJvzorG59DD4JBRyi3PSrMcTlcdasCAcH/rN
iPY95vxpLLYke2TGFhDdfrUryh2WIYqYbVLw5mOJQ6LBuxEMXSGumOUVGeRiiMY2
PPSF1huQxUuR4p/1vjNCNuMSNefBmgTIAYOIg+JWHdA+5goHEETdM18IjyrDliOJ
T260G0wxtjp04UW8eQ9+xzVMp9cXQbtNTgNJ5egeIfvrVqb/j8Zz+f8Vd6hc/8WG
og1m3RQ6oF8Fts7XMOJBSWKk0aMkS8WU+DAMwxFgS0UGSv6rWboQwk6LC36I+rpN
nQyKG+k+DKMRu0bVpedeS/QXlXJDGtLKqKYa03agBLrOsM2JZmtvvt8I9g20ZR8d
tJvGmdBl5kKJnDgSmeol+nAwMQVSDlBchKZFUj4o2hn+141S/U4Mepgye0OInCFu
auyOYFutCpHjkZoXtLVRcz7f1hEQV2P2qEg8GgKp5lF+JjpyVA5wuSwrkLC1Az7Q
Tyl75O8z/o2vfFwA6PNfycaQcIFLLEJ0k8jJt7ZC/bkR49ri3V3T03gpLTt10UxZ
GLIWvbNm7aHjXfoiKd2IXV/eBlIlY6RKDR3olK9Pdf0zz/XB+Ct7PRTYX94jlMda
xrQcv5gR7jaDKlt5U1br25G9x5/l0kC0U9wMj1e/+vMf0FYa8REd4e4NqafbUrLz
VV53LTQO3qUlX/rjxN2puQSMC+jhk8xa7CCYjebaTahAhOzwzbj8TKL67Xg7O9vv
SGHo7+ChEnx3MeGG8fHwVfTg2TcFwqgRjpPdVjRj3S7bsT7et+E0/WZpykEZHLi0
XZ+THyWEJrx151vrFpafiL20S0pZ3rEcs5xcrTI5veuHiOjfjSgee0CEJe2w+7IF
cK1NEE9pOw9dY7yGhYZiKPSLGyTHC6jrvwrSWdFqKDdfRkdJ3wZLqzADiELWLW7m
teuYE+KiVFpeEW+cgiz9WcUYWS4cSahfsriCttBy1SWAPWgTRMTP1PoMEwJaXZ9O
U9GzAaZ9eod/lSg+aCVsnqolD1QReYC0vvOfPo0IPr32Akb6G8qmLJ/IMj8uZOLU
4abRPJ9qkWmZyS0LnbG/MoXKWEI5uzy0UAtCa/Gi1bUsAVWndibta3d75ttCGMTd
p7Ts6EriWX9wfp2P2o/YzZpftvR93kPC9vG8w+D8zXK/fqp9x4mDbZIupf8q3RJ6
QofqNobOENHaNgMGZEdOwFXkrxJFAhIJucsSReednHgncJ6HAS9QpYXK+NywdNVJ
DiMJfaFiFmaBhYrnN1bH6yR11Vbcjq3bct1A+Fy1U6+urZ9CxkZvRHqaiSpM8aRt
NpdXUYDBc1q11tGjcKu3e58KKp20gCLnqJ/oYYBdQkKIBfzp/Tcs3xrmo3JskON9
WRdDW1usciBEgslEzasWMOKKlr1JHBut3OCdtUvpSrqNJ3GxFe/C0GFcPh9hZQGE
GfxA54hcnJDKVeYgD+qyP47hJoHxdfg0dG7sItfD4lRBFRdLWfUxqsqscF/r6/GC
2IcvhXkxV3e+ojSbTUsSxLIjW8yMk6JAotQ21jhWKSTQCSMPp1WKN/p3ovYmtga6
xTz1aRGR0+znQrmKcxgMKAPQW8+Ef796R3+4WgbVqtt5EjkchRhvXabyTUNo8/dS
FzxuhKRFa3wPsHcj6qxcB47d8lBYCs7pYKLd5ahMo+IT2fzWgbOsTu4fj6T3yRaU
frFV7vrlY1v4OSnrDCLTjaJV0e0cQvFGuWq/oPw9JTouCOty0yyLZpFlN/7usyh8
K8F2RGS+wH8R2VEagcUiA9Qg8N7TiQ0X57/yY/2aDps=
`protect END_PROTECTED
