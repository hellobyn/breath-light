`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yf61PFGM+0tvDJIiTRnhxkVwOcZZZsljhGs+L1ZJ7XJp9KyJBIpBEcmAL7SjiSp9
Fag8Z725FmmDUo417uQu+S6GpvLSBQRNqCwJLyZH/6WHML0poQXbYcnuYC9/YYdx
8krCn9DYDDo9v3v9LWCA5HQtqHlpksV5Cx/Rb6qL4FIhiU5nABcR4pKV9l/996F7
yL8VSipbGtxzAv84lz2OrlGigLEc7M9/BdJoZl+gn0Njm3rh9/q5ztFasjwHpsdK
nc7/4E6kH+zJLlA3lLW9SI+g90O7UbtKRo/rhDxMVcjAiukWEMIupd+w3usHOK28
4zAXbWMDkd8U18Bd4ZMFfOr5tHaCyu92OiydQaAlsrhrTK5BbHnEXE49bxlhbr3r
HX5zIUWp9M0p0qJx/iLRJi4qqPI6JWX59AsUFKmWXeN9WgQZaSGakEzrJqDRhOd7
LSdBitcjEv9Q9u3Fb4f4h8v4C+Q0s0FEC9nkbKUWuEkmHy+jsn1zi4vJcM+iBWq0
o37jW4QZ/Hi03fh5A87mwtu6Z2EhuxjWomCDHXSoW15naQbdV6WkAir9Vk+db8nu
WS2LewjFXuDbwGSzU6Wgwc/gUV/xm5kCboh6hGsrISi4eddeGh2yqjSuLPHbo8bQ
evq2oYOPOVcBsH+46UEe2gApWjpEFBc1YUcQPjdOqzKZoRrHPYYMjVQQ3YM6ZkTD
NFbnYNWFZ7Ly1JPOtw63UU8f5l0iTlg+cB5cUJIgAOaYUu8JYEn978cx4uM/nnu+
SNvkgzoMgIefUaBV7uBaBIJaeeRXX3ZSnE+RT2DSw3o5tzcpLXkAgRSBLJNCih9P
XckC3Luf6+GzsyThH0oiuMQVHuD0OMEK3ESarfJNxsWvIn4SOzJ2FDXFX8Zlq4ai
tOAG5228wo0GBVxWO/QAsn3Mcn8RFck6TTwCSQvbnqA1h1Vc77fpPGIr6GlShzgJ
1a3kxunynqQ5hy+hwuWi5jZVKKrFxVnYtVBTMQs6JG3nyTVfIEqIyuGyeBxgbAlS
84otxb257IAMLsMYHhfbWrQ2VVaDO5OSV9Tebln3jpxZbb5KH3YXoFEShBfyxBru
RdViIuxcB0/md2VLN1Z/Tp/TzirP5rDF6MxXUuD5PfDxFyWWICU6qupC1sjeCI6r
+hRCrQlapeBVI97C/ZE4n5IamM9UFz3uNPvqcGuki31o7mwqqVanYod8BjF83/bF
7AlI3Ey/wiu/+7hGuUhpXaJ8sXH6xzyIff6QZlAUY17tcFxAYgvs4ddjhqGFnjCJ
2qu6v1JsiVchcwtluC6lwO3nbkhAFDTe4jYteWMHxf7pUgUmB6DWOPtt2CGUUY6Z
XKjCcAN7j/Xq/9Z2nUs0OA==
`protect END_PROTECTED
