`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gP7gcFq++nhD2dH0UQPieuw7V6wvw2qUxxOO78C4Nsa0LsQ79kHXalfSS2QpTJVW
oaUB5TAXYS/j5klUUE2FPYJTOc7TMy5GLXWjESXpRbvVH6dsVNc+v/yOyYOE8Pxw
91vuIlZ52meSznsTlCN2+2uz0w+NSPzrslbVeMXQ4HNk7faSQQPZC7nOR2r6iy4O
eu29AsVv1q7+umtNA9BynZUAe0WbVFNKggIhTG+dvJ/zVIxyvQee6nWc0yq2YwGD
7AKpMlRVXx9PJDKeGhsLDKFXvWejYgiPtpyQ4WrpD6FAFYYxXTEI9S2SO4/B61Vv
eLPXHMVqNz2me9bPzGZ2fioMPwJDFVDesgZePB27AdPARONmmKuNJ+MNAL2t8WiV
+zkE96dPs2oQ56ZH59+ZctcYkBj8HDR99UGE5sQb/9lMoxecADBvSmYN9RKlGqPP
+TAhPMrGxSM6Fwc3phYDJBREDqjyhVc3Xx90Dn3YHcGHdsPYdrmlinABIJFMyHAQ
OtDN61zGkpfPZFei9ZuiyJWy4LMVNPOgTz8u6l4XND6hy8Oi+WTrs8DTpt/Guzv0
ZmfXEC1t4bmt8Dj2wyv9ZbNRlqzcfWZq9iHC/f8fJNCVJcAH/3aYULlp5Obfhnet
lcFpDHm2mWdLnLBGTsA0bHbWlwEHRilX3FSrzYo7wC2QNeqh88igBl490MgQ5f5w
XXLKYwuBpjAf3K4zNxbnEmJbJ724pL7arPW3VlVAE558KaC4TE2L8h+TqZmNaWuC
TNsC8lUAe171+5tyIXGvcpaOEx7D2SCHibreX29Tk1M6DyPlnMQFtvHJTtWFg4j6
0WqZkja27xRryLMwFGZ+Z+5Ca1L0RVfMvNEmrACLlx/dx80IRFGFkncaSbOzWy8v
FeXboqWq4pfuSFhbioE7lEDXaAfqbTC6wYKjh+9NZEIluA7VICjFoxPrkX5UdLt3
oGtOsNHbTd7J+3jTBLbI2DyEks6p1BBD+vx7FI7ewE02FnoLPlBViVOxv0eMe1gw
nRtrgtMVU67O4rQVdSERQT8K8hNeiWnBMfJlcgpqO9/+WurGXWrqn6DTT2o/f3Rv
57PnUXVlSNWv6ExhsKRN7zX/cmPHVshHPTM9TlKrJmhrp+vHCnogcx4FaJxNW5N8
zUZDYV4VgODBkLDGSwpzLRmIm6RVkNNMO8PK6l80tyufaUz0i9ZR/yIHWMzsmsmc
tryNdNErYrAJsvOM1Ni7i8DK1zu3HgLO98eCl+cOZS6G9pusCP+C2qxA+qD4xLR5
AECmIlHzsRHVVIYOMQ0P0EnVrY9GEKAUR0lWmbO8QBwoPDKWHm1Cb6uosXT6DK+e
SLTdgo4M7IUU49Tex6+0q9mN/oD3k0gtuU2xCAupGeZAhX9j5ivI6Zjc+2se1wpe
VfzI6VnVnZ2iI1RNqhMQZt/CtdewRWhuipznoygS6b6PzPDQaYw8Mmjiypg/XtZd
j8mOixr0k/w8P86U8pddNfJYV0VyF+IAXo+n30BbUWyowEdeI8LiKngphG0E7BkS
2SyFa/tW+cqFHDNyMdtXUUCggGTUEa4k58Vkz0k02Smg14y/+bb2oXyz9l9PxQOS
1NppvSEZYnvtQ2xveOWF2bJcO3Ow+QI/RnmWV2BMfVrmXWaA2MhLYkH9PBcXvX4Y
AxRwv9IEUUTinO/0FzgB4J8SRvB0vVgKGtHWfDQ/0tV5cYtrGM6KuINZe9oiKbir
CDzifLblrJQe04k5QZyhw1L8rsIqTLwOh7jLgpQqqfhNYjke+aZXltZ8zqinR0ke
D3lhiADYtn2kW78uhBCLJzjJEcKyMOx3NVMCULC5dtfsWODprDmTAXk3K3jP+qJV
6RPn1ZKnMO89kluGDnyoTkbPzEk9bAPH0KhvxYNhn0+/0aPLxL0U94/hr7DFK8gF
oN4NpdmaBMY5AEHSuO2C28gkqpZtBbEkF2vl0ClSC6J1GnozHHMBpkSMeRNEiH/e
6SN/P2FN2Rp3yj6tdCvwTMY1mHIpyBT3JkGCK7s/ZME3NlXs/Hea02azSTYZafFl
Qr1zuwbstpnB+OyI+ag1QPHdXbaK5jUpena2tm0M490Qxv+9hA/7aBLkZy4o5cnk
BZrz6uKQqqokkgFfAMHMJkY1HgJZYe16ONTO0CXVEZwFQXDuwC3tXIzWtZgyR9+Y
PcZCTPQh/ViYeeP8zBF787PkrzJI7IfcLrdgpuKXWZUbvS1OPgyXa95LeGaJDl+T
Ap9IP7DZZ2TX4U+98P8Cu/ajef7G6Nv6AcODiLWVI/iaWTYS0KEYHVzAH03Pgf7U
4rgD/54ttt5zvAoywz4j2FjRP2W3TyR5YNgf0Fx9FRIHkf6auZhyIGf8CaX+4/iZ
7mBPcRgQWbzDC9vBdO6D/Y2KlCvTjXqHRwgvJMEBxjllvMwCuyaKIQkGXGy7kpOT
IhXaYBgV9umoPUXKX1F2rsU/UTKLr+i8NinuIc0qjbwzOc1DgzHTAYwGyN3ufGY0
ctrhdPLwo2K/wzPtv5SUja6ildcs/jNc1ZK7BFj2/8jZtXVDudXoL+qRMEYubBHJ
oYuL0Op3vVcDIRz8l9Cp9JdqV4MRb9dXoT3cRdQAFWo=
`protect END_PROTECTED
