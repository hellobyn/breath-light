`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJVHTBHk1ZhezuyzWtTqkpE1acbgZ14RI5TaQqIPq3vE+7jYS66BWIaMlO298Fh7
QjxQnAAAK68qwgm1gH7G0j6pU4eKAPE2BhAsnIFniVGhUIUAe6RrRJ90kNfpnI2G
/PiTmcaXikTyeja4VqLrZG6f5bLctSFbuFQhSHEI/POlFdWSm2M77ylB6djFcGXb
whpJNxVtnGxiUI7p1NjywvZBpShTmuYnXhUJUTcgRNtrV52PqoIKTZGCLS/J3Imb
B8JPy8ELBmTPU2f0/8jy5T1V886OlKELp5T9IVseJsAyDeszFQvNmu00YbDK3yhr
QSmRccS/IVSZO5ap4IGbw3Jc43Jr2dlX0IOkn2bx8QElAnGeZzioBKsG3ouxHfxy
83IU3ZwHgGwXmIN0exiBzqNwLtSd8UDNG5i5qxGX5XZK0o1zWmyAyCL5gCNUr8TI
2VOcWzqIs8Wfz1GZSXHAJ3h8F0Hu6trqKZYdPRnpo0ExbhcQXQL/+7e9jppjfSJq
LRBhNkUeWsMpKSbykIbOFrfJ2em2KZglqfsiTEcJrnjYfesuQ4Da/oe1d6EN2K87
v8twsmV55lpEoP7+05CTA/pOY9wXl5k7Ib3/kva26qOXMoXwJiHHVGT3XaFoe67L
YYzrQL33El8FvO0eE4g8hSJFX2YOj9WUcCDaPqFSfME8Wz6wL2OSG3wFHapty0Ox
uEpmtuY07WWozntH2lcpRMfrNhKTlm65e4PlIF3UHOTHzPbntPcfDuf/3YbPle+n
vH16s0YbnVgO6GRm702zGkrdXMhqof0eXgB10k1MmWQAdgxU1rBtFKlpCzgPDwoI
9esh4bM0vi8uqUbyCo6IuKmeB9xIIP0wMRYIARvrb7tVf/z0oo569J7Sxu6IbX2i
eVn6TddCbBcVTX7BUYfhRee0b1SZ0uPZH1bvQ6dofS+Bz4gcaH4AtuHo5rsvwpp/
OSqiD9c5fSFHdpN+UNuHHzldKslDDGarNTR1vc8oOcEiNm2SJizh2dRbiCVtCPAy
zIfJQ9t0vEh1xGZ2nXNx2jh6ZqEDowWddxLJOCjFdckLNCQyxXo9HfiMWP0WsPC/
iyMcrxfc2SPf256NJ7/li0UnbMedg4n+rmqLc33XutKxPfl+JIynt9+3DhO4e0lA
XZpjSEaXi7tj39KoAejYfExxTEuNOTdtzq0xB49x1xzB1T9kZfOIKRcXbXT3AKAc
jQ3EyFYsLwPsX8kboIt6hkTupIi/dN9xa2KuzMcb/OZvMMRev4r5lyxAydunmPM3
5C5SPM2/YQIVjfPXBP8affxAeqih0MdihMil3NLOLPr8ZqfSZl9KeuZFLigHvLhT
1iXKEyribU+MYZFXNq77nYR6NWTJPhfuvpUuFOjPujFxBnRedAV8WKEy0FiAq8Kf
xXxeztXs7iJiNfN+rLGwqBRDAFek4PKTyUY8fnSEXyunBZ2yvEWpyAn2wMJ7Buuc
ZHr1KFhII3JEgI0y0avBstEy192p1jaigAm4gNXXr8u2aeZmRq1PywKPYXrv/uSQ
7p/kiYqVBXPe2Ebxyq9awJ/8GEbCutPuAceX9NpCe8g1ud8Cz2GlmcIn98pAUgr4
NFUmNr8ALByoEbGneeXSLfbPTk0Pxu0kWi3tRy4fzcxR4qT89TfmHy7QFMgG53Ii
sGDfHAjo5icZjzb2mzZ5RwVYvoyjS83QJkyF7Laij4gz1/EsmodRnw7JUsmhR9C/
PBfL4JIubR7NtxsF7wpF2SAzBcbeMzF9izzOeGCMieEH2H9EHeDGludNx/RYC0Lg
7GyuwCkbTxLvMzubevJRRLiwv1UyK9uy2W4a4m216AVeFqMgMvMXQg4PFfhpq1Go
U5toqFUlxnIDrQuyqGtcxg==
`protect END_PROTECTED
