`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vi2lsMDyGKvWnaE/RgwOfkJ04ix4g6wOPVFYt5q7an2ZffF5EkbVd2N4TmSEL/uq
2vSpeQe5HOkPzewRvmmCzH2jZzXZ6vbGOBPZC/KC36dOD/TN4Z2tsyBlsVMxLJdI
8wKptenM3+J5LA4klI/MuQq9jSumU27PFOb1G4L5e/IhcCkTr0n4RwkIAElSwESz
m7o4BYfogTMaINq7ZCt2UpoYihJ4Z1hjxc5GDgY/t1Ry0Tu3hke4Scw51WTJfDeO
cSij4LgalpY+oVCgtBAdIWhrNlehEaatFIj6kWHl09d/d/waYxIlEzf+GJev8Ec4
vt/ghWhU8t03+TOQXnH4mDGZa6aiNq60U/L0ODxhK5RD4CYdb8v1/jA4/6cgiOE5
UtNM/ZUNO5TvQG0IlIfsTsHGEPNdsZ3Puoxn5CKyu7IsgI3ze2jtGfVenneHXEHY
J7SvnBupqvTAos6W5t318kecakqzvD6Z5J/TVyaeoM0fv9gxIFaiZzD5ThMbaBPa
q3fyTynZP5boQqC40rVI3YBECYxg+Bv3EwIL4vr7pSjh0z6ssaS8xXAkHdgRiOzU
ySMzQpoX1Q7m8byw/NrTTCsK8dsWSMf0yDsABJ7Sc9sNfe30Nnhxn4iWNLrhOdsp
BwXoS9Q9BvkCFkCRMroT6WGRzLgSGc/S2YPfbVuSZ6P2e1UcIqW8USY0r4ONtbOt
eYLHO3+P1UTLqkTLBfliHmDAHMYa9+U5flDVk106N0StfoqkG+A6NCdhQH22pYlX
kSoNzgwCvZINQzVwn2/6o7weQAkQDGMBPVoG7jy9h8M4NmfeSdBmptXWk20NMBUu
BM9+aozftRZk1/yezopQnR/EJffRCgJCsw1Y0wOxwZxc4EMGQvwiYGDo4V4gHuyI
2MGkIEVA5mq6eE38/t2Jq4kxPIGbMKEXRRUCvKGc0JejAzCY/ntooNsGpS7mnNKr
Z2cK5sZVAPqHvQHmdQZXZ126bdM3qwkoOrMS5L99V1+3Al0v2Gy60Mm4LP9Qi4S3
Je/pJy38x5Gj5brd2csb/9nn2eCtWBDYZfZmaIrlzX+0wyK1XYSXefSV8u4emtZ6
TYRbddObR2sZyQwXwi3uyXX8lavXtNQXqTKJS2DZKhHrn7S7xoHgVLCKIAnRdrPe
77EUI30o2XXqpUFMRFmj+xp0sKg3gTh8mXX+pVhVJPMFRSRTxHQzFQWmHXWFJOqS
`protect END_PROTECTED
