`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iA1R5f09AYhFPOshBblTqudm5Smr9kWgrSDON+81hcWD5ab37GM1ZvgkkcawFR+
Az5p5qoNBXhZo6RfwAegsXWJywL97/FuAdF7WzIC9AGLCxrDkrWJaknq36MJ9QjU
rcJFzDaQ42lZUJWcSST999LWjiXmqqmkC6yCAFa2UTaFIgKxnhNb+skfRY0arAr3
1Kfi0L68Dq9TOSfK8M6n0XRztYO6VcZLzu9EBggrQQsiFU6EFLadSFEcL0PBzRWD
n8aVevZjbp92NYBM6Utq3ahvJacHA+s8cbefCEJIfcNFM5WglYsKjpMEulej8bll
dwHNx6Yx99FKjs4HnHg66Xj3JOLAhRMlItpv070X9grdA4tUUxVVicI4XbDrx1Sz
FoKeijGp/BYwMGhBT1mzZ6Olf+2qSR5q/CZ/mMfwtu30TCJtLxXZPe6NzTuexAQ9
YgsJF75lOKGJAZjpU3Fu20V6+6hYF3YbChVNG0epxNz0aEoZJl8VtbwsNRACSePP
Urb+TdEMgfBBGyeUf/m8WK6KZHD2itrGQ41OzGv8sIqjTR3kyuOj+caVDhemL1b/
xxllhaxscUtEaxnsHeBBKYBqtClkyZKXNVYErBffSRwi9ntsDqiLLrliP4wz5yju
gzNN9s7kaWUxAk8KgClibQKfp4QqdTUWiWGwMqRQqFFkbwamjqE7Xkq0/XdtKF3S
Cy+Go39FP0y1/d3sgvR6L/yRRzrOuRJDJ9NhA5C1/2pIIGVtjYLmmUUkN2qYPOUT
PDW7ker+vupcm72lf4BJsftwGXjlbhR9CuyARWydO5Hx5VFlUFPGBR52wH+30XRw
1rK4bgqsEmi4EIgmMJJBBnby0dZEq1LSRDRUKqLdKHfQ4as8684zZng5hbk4ZgmZ
mANQ9G2I8I0iWnxAxoStV6+AXesGzcPUMtAONOf201bQrUixziGfJW7W02+0wZxm
5Rb++gfIwcguhYBOlH7PSxa/pzyD/JFwhsG7LeIyuLVWLGSRBl7j1ojwKhoKXacQ
hJLIyxUjTb1WOJmNkitFqp/j9nzFFD28yF/f39evYvdmtcztwPBps5uRt84ETkog
wsQZkqQj3cFLKhPNsyZW4K1Lx10+hwwuLTint95GS2zsgGiWeBE6wrnmQu34HItT
3mW9+edT38EkvxyVf1RyYgvxZzX3OQ/biPc4Xf/bee8Fmm5yBsvaI/jyRlM9qt9A
uPigB0/CRXiI3DVQzf7Iel5eTlTNjMd4MTpjZ03aHRsr8i/UNa6W0AuqrUhnr4lf
a85F/Up1AtoUyiGiIN9rvQ82GYtX65dso3CfVmrV4UByGxsbYfrmXEdhO4jGv8GR
uwUqM6sZP3q45do8GFrGCPq9eym9x/Fo+V/6kEvdEG7E/4krFqLdrqulh9V6J4+s
sOkb+xSsJQF3z4QxrbrJXPQMQHDX+mKy1WfS77g+eecaCk6o+Xa06V1kd/nfXD4p
lWqOCsGk3/B8eEZ8ziYJn4MfDhzG6hUUoISIDi7Btplm0UeHrQykffrEDIm8aGWy
pFM/Ct0km54a2nL0cBH0nol3B2Hs3t1woMq/1l27aX/w9t86qrkkHuXp/hKbgA/w
uHHrnLwgim7tzRYPIyNIx5tZ/U2/JVRicUWzO9Iyh2FVZfcI0SDilE+KEdKDpNpx
8TD0j050ghnIPQSCS8wVnKorVvAqMCxq/HhOvlFJiWntwQL2mXxEmCuyyq13ayPp
b9ZFXlO0wTj9K757CSSgpoe7Nu63o7SiZKiDMPx9BbktWgUf5fnHAk5h5ayFDusE
sH48EhrfeqvmrDI8k142zN5aN0jHBZqRAWRinJbDMMwEn0kbzcoBkk7i19G0XZeK
yVd/OAbHpn9Vh+rEjaBtY6qCAaHUQw3Io+5p6JMcqVOhWm2RgSeXfT1IezGcPtPS
Eg5TD6lW12qjEeL3pqU9duO/MUjDZENbWOM/tVG7OQOcghzxzRNyTJQCKSZ0a/uy
BTR+JswPaZARrxOltE1G7c2Dp4j+OjEECKcG9lAllpR2sfGSIBidvfSEdZ8g8TiO
UT0QNU1hbQ1b79VVnGaIDRT+X78Or7Pw5jR9uZsrEj4U4WlBFRpZqZ9Q4C+dOvxB
hs6cCctqq7d0UNC8Gfzdsr1txLz1PMsa5yF9V6K3qUAtK58U2DsOfY5mCLO0CQjm
buL1zNrJVQ8c3E+dBaEKqGTWRCzYjKO47fb4dbBSFnWupEone96JNpFcqupoDBQ8
t3e9vkAbh5Ze7Y4QNYs48Lw6ef+u5vW8stVBFWaMjKlj1/4ZAsMVfDYg9V2TLC7u
YibTyfaEvyJaO6Jto1Gbs0JKHT4NhMH9ypfodo+DWHbLQi0mHjg8myt+aobn6cOC
pQhzvGAm2ueL8BMVoTS+g+1L8LbHp6MqL84dlBfXUgOPJg836ViBiimW7C2Liy8Q
Uen9XNsN2RoGiq9QwZD/N6dIKvdAfxPGXBGJWM/NvAMD/TsTf3BoaAPva447RwE6
Sxl/DT5uZ9lJlgJG4oRnvyGitKpBqkxED6BzuyRmT0xLRnXPQc5vZEH/fqaL+Jq6
XH/5EShOmJlQUPzLgji3rVMJ6YiwhIjib+QqF3DGzaJCBMQeup2QMdStpxeTDyZp
GPF5t0i21GtN5Z4WMGG1YKbBdg1D9S/eSGtucSdGvAZ0epi9NfIrzHUSyLgUD2k9
nBD7Um8eCjvMpilPZkBjOOfFAkM0lvQKDUMX6QHeQbaHsOjE+JHs7Paloie57WG3
vCm660pTvfkC/mDpCQCA68NTQBOFr86Zwa9R9+/lddEfU7fgmdK4uNGgsSu8dT64
G3Qa826d4rjlRXtkZmHNWHqf9d/SMtLEAG3YM7JjcLeOL/SHbKJ2z9PHwQnWud7h
R4X8L9XRbcNYvJ2q2mokBdulnyC3CwKc7f86DJIw56G44ewq5ccJuiyTajCBK4Oz
dq0+PsJCxuwTvzZQaU2+WgK5Wcd3ref3+uXT5C2Yyo9q0WSehYROzlBXpV/QSgDN
8BfKsR0CztFqCSjl6K4bQ9uV7lK6tpgI4NILTtjVwq4XU7NsExzWGfGWD4DhdqLX
LTynyEyK90EKzqAp03Toyj9QZGUeFNhuP/J5zn0CUikk+TQPNFY4zv+SWrxdyL0O
11ojAWKzyd5XJPQyzpKz8WKpFd7JkIw2XfoVAFyuc1BldB6uogdUbH8QuL2YoMU/
yz3LwvkWKsH4rERd//dEEcSzVvHMQNZCowlnnYkGzyyC2pezMyIiH0BSCiPx63Zf
kqVf/Xn9+zeQQoMmD2sch9ff5K1yQjWyQjA+c/Tqf+426AM5nxOEew1MzbZwTYR7
H9Qyx5cFeAfyhHwYoyVtkQE4StTuv1PteuPAqVvH372PHAcxaozBpROHzGyATabd
8CHD3S9w7jdNdEJngMP68ZMjWwyFzrRoxR6idBOIEPVw8VJkpSwstbnUIU3DUoAS
LZFVHSBo5HNmoJ4LoAe12j4hECDftDbNwl+oMdBgpjYntDxBdkLjboLbG+xCPyMK
/4SGCyHS+rJVG0U61T5oRv6HsBxzX1DkAuE/gt0tpKhiZOzP/s2OMukMfSufxc9d
gPhcsMA4upNqxpoE3+4cYj8EBMgZwabHxJkS5jDcV2eAMwhKvEE0+ZmWux/RU0MF
AqdYF7dAK+fGkmRNWlBbmVGfOdcteJMir4lFc4kEFPcdhDUQZnpSw1Oosj3RJ7XP
ngQl5fDjQyADPfbo0P8yAS8l96uy/ZE40G8utRB4/e3sUPIMnboaoRr1DCdYOv+Z
7Bp42P1ARxLX0In+BxkM9bcPi15Cj4mIkCwG8i2eYaWr5OBZXfPMzmtAjX4/8DtM
iveUC9QQlPpG/Z1WoQ9zAfpqoN+q6jkE74F1EVAck+tCrIUMYfGWSp2y+oz4Th78
TaIxNV/jD30SOYYUwg9flBeVJ+URo3BkdTpNeJaxd1dYBNTw82PHlHfhNs8jMfqp
Mnn6Bsem8Gr5jUwqaZj5wQnOh2CJgUFzHtQz11a26UXWYKeopFtHJmTL7RAgNccw
OY/kqQAd7IFYyZqxQ03Vnrd6lTfOEKxKWM1Es6aC0lg23HhMGxu/vQRvYaF9Pw4n
roeAcbnYpV6vQ+fgnlU2g7j25h2T4NhEq/8Xpnx0MUMBPcf2HtkQAznY9sByG2el
tna3iJTLpz/JL119Ij9W6bI/yds2udWuIBokMjGONOPScObAdQxA6VQDViB/QKQZ
GuHLEq94iwkcxjIe+alH0qjB3ums1VspbsX7gFVvEtpHzxNz75VhLIWIr0jOo1Q0
2QInE9RyQ9NhGmj+55PEOIEOFa9stcTf7Rs0d72iZoGuZpwmliiw/Y9eI5Ph4KIv
wI7HF6eI47FysGbHt1cDC9ttpm1BN0/BaQJU1fsfSMPpYGQ0SNqUBP1WpoZG+kik
OqRXh3s/iJds8mvh15o8pNGPXET9cgqYTK1R7zqVYOUHs8FgqlWOssvw6cYhvAU4
55ZkJqXrATvpFZxCzEvb7brtd+LFL5SeYOdzsSU6rGd1M2GCR/pvprYXt8KrVve0
A4H3yjtvyMo3/zA2XpulU4V2LeNwCGehXjEyXN5qHr9PATQm+wdFc5dlEscZSlD7
8awSP8D4CSJ3/sGxb/xLQt51MBIw/Ii164ccxA/NnZ2/MIQQYGUH/URcmSfKQHGB
RvPU2Ta+vk5Dpl4N4C3/Xob/46Vh/jStltE6nJpUXHBn1OQEp4KQVJk383ZZtECz
bgxPoUEcSDjcWW7ycIh3t2/3e4s7BwNTEeGYH821qBfvfHd+xpaqI/CprPg29ApR
4526bMYFtntP0hm4OrwZ1lZLDMR0BGgDmCBbDgsSml7ZrqtoqwDlPyiSO9czu1fJ
+NK9U8MWM+kn+rN0e6ibGKyNy1bmW43l5pn/DLAfBcFjdfihIEp4sYAiJpp3irCi
ni97f+oNbKWo9nbLs7VRHxNpe0kbmZGAQpfG+xZln7yxUjqQhMsb2dmr7hkOOMPp
6lapW/Jtks4k78MEeqd7LEvKez2KV5j5lKzb8hx670YR59jY6CTHOvJvKM1+k+B9
BsNJN/JfEQvqEmv0uc1PlCEsyxJME3+8TiZfnMRwoj+Ise6uXsduxY3TF6Z8mJoF
QiAVMMqkFvLBIw1pWlJwKNpBrwKk8DOQQmuLBdwD8/stc8jXiZcJmzzskmWCEx/N
303Tlm+eOWg6zwhn3aNlYDUZLpIxE5qFTeFlPUmxonIdMLiWvumu/YWn9eQy02pm
XeBNm9KO2kG2oSguRZxMUTWJnkd6j3DXLylCXJUQMOkC8/DSlzGYZu8y8fUSEzqt
WwVHfyxgvjAU76fRb+BI1rIs60Uj5RVTCH+MM3epfnOqxG6Cg7mMbEjASSNgt/7U
6qj6BbrR9tg44a804VwYQJ5PPJ8nIRPfWHEK6wFAx8YV1QK1VUq5HQHxIuIBsARN
E3+Peiw3KzokMRIW5sRYbNoazYnWx7hq4/vlhoc007k5LDPRXyoPjiPbr0oy/B+X
F2+Qr87mFjYSLNy5yWrsob7PAEUevVrQOpAQTPRc9/w=
`protect END_PROTECTED
