`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lF1+kv7eyfqaY5iRELE75BWEIIFIP6s72tZDf/tRO4Q8jXWkit0iS/1YAfsC+suQ
uUD7gN1sfP9u/TIJejvKTNjfoUK0ikDP4if2+LI+5KuCl+CdQIg6uxw/NcexFxIy
VzpFUCtpJJjAC0VKCK+nlSxhoXFD2kVWjeRJCoZJvSRTf33KJP/cqeKR6D3m6v5q
mDyvLleMLqxA3KNBhnI8yTQGPRwYNbW5pORKh+ewV7gNfaE13zKaGPFjcFZHNuZA
wVGyeDcLtYV+IwkMAuSrhTMNwZh2cVCjW9y+qxY4rwLdoSjfrw8ffF0ZnL8adUGb
rd6KpQZLbVhpisrM1Oc6Wdzs4ubC0UXxuVIGahy4nrl2P3t1FIHW6h4w7YKJh5ta
Q3r91qGLzXK2WlQEKX4EDKSV7yrnfNFFS5X8cfuSkwM=
`protect END_PROTECTED
