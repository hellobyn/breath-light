`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4s57QpIDQobtww24Yk2O9y2dzoSUK70cL7rnrkcga3Yyysuw9u/2in1hveL9t/g9
KXy/sgF89gCOqjYprzeL5Nr+nN2Giy5boEvehk9eHwDgAn4JDO74KU0pXuKMrDQK
k+MEf/Ic40JOs6zzn1iKzWv5cIHH5pb8+sQAy8DMWQcIG7Ux8MrtIFXFHb5EEgzl
LU0vL2l92qIh52Nhn0eOpHXtSRR92z16qiqAIwnuQBI/xT5/Qbu2J5f/a0SjodxJ
bCz/BuByDZ6lJL6m4WAia+lkYMWsZutlHd+4SrLh+Pl6sIOJDLjusWi2G8BAKY0x
BFKHENVnRDDmZ0X4rO+hvoFt2QPfPiVOVV5tvZucUBYwzTjuxbhOgWvHKGcbBf8a
SqNvqCehjaploDxj8tclQdgaye5Yo9g9juVPNaZlQnjWQqJIDDmcBMM+19C6wsGN
X5d3iS69J0tsb85RLt/cdARA33TPS2YrOCV9jvRsiA0Pkunk4eW2qKos/IynxhYy
NSzWhCuIN1diZy66E6a2Tccn17wLoFBIC8JL9G8cqCCSnkWKxVuvJ7Lh7fsylS9M
FYK/HckCYJS+7+UUc8/cZGO7I8iH8RYNT8HfwxkXhoXAZdDS51imeOqw5nqQ2Ffn
Q56lqHgQhqKo0g1FmC0FvygivqrwKdu1Qv99OCzmSPaY3/MvjK8HmXhWBqiMMY1m
OvGiNCp7JVcdF9Tdb/mpzOdLNd4DMmcm1489luBaUZV6WWiwYf7oQ5WEaChcMEW8
oc9EdlgH/cIxPqYDWDIv0CtTW5EzDNK4v2clTmyjJ31NEdcuHdjHPCQekrwb16we
dCfJP3smCYCk2TCEsDVumk0w2dlrH/ysPZrhnDODXkbZkvtDAFqWYH9qAcWG1yzF
pS2+vwkXHYeE+NoT6bJ6NIkcvRk+BoxpZuOEWfzI/MyhlF/k1ne+4AELkUiz3RGU
7qNQ5KumTMhwuBCJdTt0Fqc7fHzAdpmm4NiIkygPaHMdWVfPhZwxKZ4/V0hlY3Mq
ybRxWXy+tz7rjTNHJOvO9/Xcf001aaS5WAFCKjX3xLk6iL8JEwy57bPtwytReYVh
s1MjWa7ko36Pciop7chlHZo7szo8mMQTZFPwVqa9N0TO6y96yN0EDMlUf6emEf/R
mND7IC68KO2DwIuM4WmcGhncm2Uxa/SlcZJJneYYU7ZwOHa3PBRvzvhswapidiGE
0z0B+O0OtLUi2RgdJvMltpf1jj+RwW1waB4hEIaec6hjREujOfLyZs0jKDluXo1j
KVPiESQ0sNP0VY2FpPuTs+m09nxPMVJ0MTcTpOg7Ko3KBdZPUSmpP/jUKOhDtu7k
CN7EJNzqM2JKgsZP8Lv3HFJU1HBHY5r17adf8kfDxgKg5g74AWxf/XLZhSnxmZ1E
ARgYhFpb5X8KB3e+Zpw+e2EKnDeLMSSNDjJRMX9R84I7pCjVUc7NklYbXVjwJPWQ
Dkegxs8ySMsZWaLhT0NJNanTFvkdLzHr8Xcoiw74cXhVCA00NAgFfQ09CelR0nEL
`protect END_PROTECTED
