`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtPw+GAGI9y+j2LX1jzbCc7kBHloOUPBJZtxbsFndoS+97q/TzmaLUNeETItGluP
nAckHxs4HwDBG0C841H13QD8tyLjhRlhdxaovSysVqly6rYXPDnVZxUMbd8/o87V
6YUMNmBjhsAhmiTgOcPE0MBARMndWL6fRymrSmimZyjaS5HLfgjupiyBuGmCXr6G
civrbXp/8AqF5nlh5f4AlX9YO3AscOo2qdjbtl8wshnMz/4dGCOpJaTgpTbBBdeJ
ep8ODq64fIAp66+j+HKv6/YVPSQSlkssYXqlFO7+elXP0ARAnHtE3oEPC6+pWIMs
ShLYu6CYCO6A+niywHk8kPjQm+xGhOdwZBZh1paGgKM3MtYU9Q2o7cWUwlCdEgtQ
PHN3V9sjPQ/X26OzDiu189Jh9EteusDwNZPLz1hQ0aPQLocV+xanYkX90R4Kf8zL
YJUsSClt0kv5YqZt0vci9oNfxPaEk6NZB8O5fR9QAsbgZMEO9xaMoJAYIG6XWpk2
vJDGABr8Fm4C3jWu+LS5/Nzb1N/OIVpQpLrmLjjElDljt0g7P34vv08GyuFkCNsa
AJ0XmGzTb4GCpPSMjIS+oePZCxdc7Khwd/M27S7Phmt+zaT9KUY3RitXn7ifdHiz
W8Sb92YJS1bFcWYQqHS3paKcdyAgZKz2rV7/3N5OW2v02ttijKh51j9cWcnFgCyv
FVe1x4130Q5VMamzet5JpwogBADxOjhiEz+ZapZiHdp3jQaVrRuPEL8letFxxUG6
VYevZHyXpwo+U/G6OvMWyp/Fl1Zg/jBMWJSl0DWpwZzpahcjhMImnfdZyYtWjyfe
eGk9hBK/aosZEzR1F8rwueGBJbMk+h5n9ZrO5ioN3heD7n5MmmnP/Vy1ZkeDFQlV
RHxZxtap72XCpKW4FY/95L6RypChIQXc/gkn5a+colLkPFHbdJ66DeZpqDjIwJrq
h2KO7lfQh6z7FpKUk86eAmoCnYi27/dCZWQNsNwId86GTY5EAx4uaL9knxBZakof
ibql5O8GF5se7CJqBey0Xx03mHTfyfp8NppUuLzTEYRhr/brurIYCFDnyOrvZGok
cU/BV5U58BJAjQn/Wj3wqWDRUTd4ItnCYtY4Gx5Hrd0dj3L0LLmdeavi7dyts5ew
mrQmG5Wvp5qz8Yt+KrNwjJDs1hGiqPf4KaQRVIsV63L7rJscm7mj0+NLio7ciUHA
eO+fEJuT336zJ43CZqD9YCM405rgeJCTdaFSB/h4EtMXjG/ly3m9FUsk0Jwb67tM
hGrQjG9MHZXp6rJhS6tZTIfYpTiY6PM0r0yI8OCN6Q9fKsESX8buV9/auRQSIBf2
hQsSviYFVh4PDz8nwmSBnFXf3pwIN1ULny/l4fa+Qa27a+5bd44hwg7YHwidTj/m
L2cQVlBr5pjDvw+kes42c2k7TZLiu7HSgZPScPo9qEOQhzWoqTOWDd0Ram5iAABY
xLPKvAXjM73FHYmkX6WbR+3ttaUa58sAQcS4+0lUagpauR4msKKMB2lypOS/TdTX
sEtnqQLAZh3bPl3VGVaLbm91OAsRZuR90C8PApxaComnB3ID5L+3NXQIBlUXKXIT
+p8FJN3DTp6AMwsdI2HHSszLpfeQrfNmBmMaygQkvVksER+2XnVUax9HcADMtUqI
l6CYgLByYS+BfdmpO8iHtwvcVSznhkdBhgeXxoU4gLXQoXIKeR1OSS8yZXZVBaEo
+OlDHNKZNBOc3hHIHLpenEpTlHhkZt2T3b0mO//BwWTMPXhdv2XTlLWK47AQNGfb
CViiigQx5aCkBZlkL7yC4TcTWs4oepyBhEf+8oUKYLorPDhy+V8+0LBVCW6qGZ+7
96fgOgnQmOhc0YYl6y4hLGjcyI0jwRU0yEaamrDEqaeRBt4Od6pPxEaM4h2KVwYf
F0Dtqm3FV/k7WhSh5H3D1LiB/eyqcfNNEOrTm6akCbBmdUP60bFGWYNhZxP40T5M
L/VXe8hdLAg5Q07c/4mdzSneIsachzf1J3qcyvyI0YX/gaFnRyHVZWavFJ6sD2/y
IvB/J7tyNRkmYCo3/Cx5E2TigMP/GgGRW0jlfo2jLubnffdXAF9YE+WIbMMQKYrS
2/mdnZIk6PPhJbsEzPhGAA6Ntk2CuNv0TqcxiZdOoSncrbc3crImnBFU6ifY7Y2I
oHUbOl+qZNXWM+wEMg8+iahRVoCPHJcujTBS/HOskuY=
`protect END_PROTECTED
