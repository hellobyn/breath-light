`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSA0UPXho/wDyeCiKFNBS1AP4eSPzgIa/vFAQ9yH8/WuwmiCN+PdrNz8PNpacek+
ZKSbCBluxsz8bBI2BikQnJLQ+p4hd8g/2+cRvwss9amuE0ItULFZSLNSHoRcH/Dv
e+exdCJ8mz2y2WITEw2NNsBv8adTVvhs2Y5C9X4P/lG6HK3ASqiLZkVqtdVuLjBA
tmHKeYNWwe6Kj5RXfQrfc8fbAjcI76QVO9NB4s7t7ZAx2zbXS7uk/W5gYBjP20JI
9ekVuS/oW/00AnI3A4+fVfz5sV45LObQ5qDbpNhQ8wfStiJHKeNQOB006s/QO4cH
3FqZRPZw7+XFlgqMejJMsSAIlArxXrCnWmsXvMvFfx3jAabb2IPM4jvrhdoDkCMo
QTYuGtG4lbcofuDv3iOUIaHP1QV+IlhWUSRgpccdenpkW4e+i9AcI10c0M5Oqz1l
7uVwDPgXEv5Ej+I3EPraWQtYTLN68EqhDgL0PFRiIHDWBJSr2eE3FySKuAe13ZHi
/29P9soduaDIza6K/fWJ+x3j8OOJj+xMJ3HIUaQum43v/AE5Dd1UWb7cQFunTIPm
vL8JmX7bYCMKdt/PdpegqvGHQJN6qhdr3IFN//i2awRYYicHr42R5rdOIJ1G8No/
u6+CROkdosodk/a9BHlBetUdXkyZ+a94OPx15l/4QrQPv7oHxgtznTd+lnopaTQ+
ZkvVTMJMOWvXA0tUP7SNxUca79XuPzTsi2i3J0Yslmo=
`protect END_PROTECTED
