`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pqyrjuoxg9TOOqQ+gbwcyJ9kKiig+V7/wySvWFbuBQo/OSlpK/uzQuforsR+0huX
YFKeutvZXG1O56DngUtkCAh6Y7f9LxALWGpg+110ZzoBoi3zTIYcDzSUEn5CnBu3
QdWRCwx6EjG2FB7Y6waOJvgMnSLh+liIxlBN1ACZU53+BfhzjM9Qj7ZyC7fXs5k9
lKI4Xez/jWC+cJtSbwPWRKg4OvuR1hc+Mo3qpHlxVoiR/dL0ALSjUhHuUdxStSKZ
XR4B+IWXSJviTAGWD0fkJX7szHhCot9EpleCFIZ9KCG1bpTES/WLDN7aE+fpE/lc
60w3/n9/it9lM1PnfDdyoVhp0MCcIyacVNZrmCTi+Qk5qgZ0iuq7WZuBtyhRxsNg
npdh9sqsWyx3fzCEc/zo+MM4S8eIV0e7GCp/0WkRWaifHTcofZbvnfk9c1LAIVbn
ogT+fMrt4uXHZcCeMHroVTUvIuCOXwYW3C5CLh2CIEkoBtRRiM8FrmPbwSkNmMY8
YDzR8xKYSfW1lrBO9uUZsKNu3YoHva6zJsZsS/Zcx5CCU50A9hxik8anjj/ctR9G
iqBM6Wa20vEks5OYfXvPK09ihc6npc4y+Qq3q6/hRPLplpbvu56iUyGYuj9cD3U4
Q+cF+cOZMhmI7Szo0H8eiSQfKuJQwfYM1UCyaE/JcDvi5vTHHuzWGqAPOPPq7r/m
kwxbp2chIvPMN1BHH/aYMmmsBPs0oFlWxPuk5BwiXTpJPDCH5pAm1JUHWVDsyJkM
OJhgifPqZWlAIKeLJ/Jk0YQDogo+p7CCRamB35yJZcSzBG14wVtLPMnup4QaSCRb
5WZRXiZonDhJvB4jFxCsmgSSQ1JkcPs8EIfJiZqMf5b/07o5DH6dUzQcRO9jX/XM
bUHdC99uzaTm+LrxTAws8pBDWC4eJFa4UuBc9Fdr2f+GriY85XRu+evSndAT7vLx
wgdRnIwx4usDMb09AXEMy0EJ7v6k/wPz5yX3BQJY15xAN0FCtiDo4eMGdNgU8/vq
X1EJUs6xqF7O+f6sTadwSvi56XHW0ep/XAMx7JTfYzC9xGvP+4ZWgKMQvOHcgz+h
11MzC5H+XioALbOr72Js2Qkd5w3jI8aHEFgpMKZDf3humZEL/u667WNNISEckl0j
Mo3JhTFWINy5xUNsdL+NUWmsazG8f8GmPliJnxMVzwTysoDktMIy7PYFaH4HXhJn
y+TZaBgcJMq+NZ7kyzZh5co0T/Xm4litOfUFD01/Forfo1L6j8nULB7umGxPD9av
nK0xWGhMosBmrttfmC7ZQ+9q7IaBdWxdYdrkITrGC5tFqU2Z6XtRcehiyhLN+LmW
LOZjOEotPRcP3Gb+2+bCVKRxX2QzM6usp28i3nkkGm0=
`protect END_PROTECTED
