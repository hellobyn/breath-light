`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7RzMeXW39L00g/mh5J79BEGHN7c/q1Sboex4clJxTu3q6dttR0Yqs4wu9XID4xq
3koltCuBga5luHKv+74BvcZ+PDAsUxKDl1Ya68ojKIfMft3L83oKu0v+mMz+KqFk
WVFdHNFpwuNxikOl5EuHCiS86TRP3yhnVRQU/eFxNObkAHtg3c/3VEhLhXW5uE2G
Bjj064TWMhf/hqqGZnCtzbpXS3oRqxZh6rexaICBzWB5BSFgTHNdTeNh96QjvnVV
lzgx1qe66IR2gWkr3mLdNu0xLK3wwGSY330Bku/8JrlFeK8pvjJF3nrMurvvpMx6
6djWUziFG5dtd36IIUDGrQJAg7Fk2F5gY38s3y0uEFaVUi8lG80gCduTh/SZKN1C
cYq6agrEsVyq4mmQdKO5PBtmEUNNqxjZNjDvQeO6bSHxVLZpiaEfRMc0BVJB2PUw
rSCAGZh/VpbZ0avMNmJG/FxXfHXMR7AGBEzEzNBy5o94JPgEYJjmcZQW+gQrN4YO
9fOqY0pYHYB3AEdr1N3vfwtD/+A/t4+IZfQ6xlFIzi5V+pWOWFLtJdQcJYhvoRFb
npx0WYeaMCRzrGCODlDmxp/ucTansjrFqoNWXmh1atQNh1kRJvVqWWcqu5OwjS8I
xoWX01l5oPuXwOFaUOfuuS8e387LlLFs8MnM9XEaSu2efP6zy4DVOM/xFU/41uuM
4bRgBtefbNEaMv4Pl6XLKqQszCegtktpAXzOyv0FWsZQ5djg3a2j3e2HfJKCVhtQ
k+Y1Fi+iogxHnm3b3neDJluzvPu3hY/f609TrSxj0yX+Cfz8RgbGGsKKipRmRiEv
alnIp14FjOIxA2cEFR1l+U6drckhkuXY+FjBmAFiQ0dgd+cGcEBCkLiflqn3I9UF
D9h1seTOmT3a4vDZFFyrLBgHSRQN9weYhu61ZlkTUNE=
`protect END_PROTECTED
