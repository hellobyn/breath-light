`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
blNdY/Z+dKZk1e1gwXWHCNO1yzohpknFRb7Wm7S2SukGBMUmXv5EKOObZBFdmHcj
FURfoE17EJckeFXyruTJKBwgOIEMRLX7Ty58IAqYVznaYN6s9LH5pyqVYc8pZDN3
9A2PaAuT4M+29BGzj3JztkrCyohIyb+l42aTDoc/hbe+sayjI0JNFW6JG7aAiNvd
5dilFTakiT0zl33iRkWmbFSmCqU/8r4/3YssoKuXEDoW6VXv9SDB/IGEbANFnkSZ
50KFAU2gaas5ZMQ2ovY6bZ9/MKpCSvrwu1OkzDhdySsEgawtYvk1MZ7M1N+vaocX
mNWLtQ1AoppERR3EChC5Jq7jZphPwmc+3EzyTtbUR2v/4+5nMM8NfJvFnCPZSx2f
KuoNPJCdmI3VQZkXhQ4E5g+RImu6c6BOVSCI/xd9onV0POUNp6wB8llGrnR2yssa
g/OXFFilFIMTQHVGBqGArEAMPkUmB8Ko9X5jRjA3O/WD7WkL0PvVPMIbquoFPnxb
bCNd7llhSXlX9enyWIybG8xNSjpGqk77AEC3FEb3NBJy3G+zTYCR+QZHOVgNco2Y
Sh1whDSiTBSXHjjwlmfOVucsyODkg08gOWfGtpLJDYFNYJ9WUxwHfztl2fDPXsXT
IdSg+WOfAiT0BU5qN5tonOYUFrJ0vfLQ6GvtQVUr3oiRfaD/WuArtoTzjr2hB8nj
4u6I7gJK57VDHA0j1aeHQ20n9ZX2si9eTLmQn/kLyxl2T9iOcBaQDxnqKLLriq1m
xyW8O7kXgX5a7UMBEUxFnMi0s2Fn8NAPxpJYSOQumB6McijQlc/cBRWJ8n+cdvxo
n/Cl6YG7/zYM17Qo27HxTfCUrq3q0fnJ6goXJBxQQfFyzoJ2U1wl4fnWZTqP/x4q
uTFTJI0QmodOG8hx7uTXkdE7lQPEv6dxGHGV7OmuLO10SSysZ8+Sg+8onkSaaeB1
xHuLAa0YNJjySp3ftlyfnpSNZ0dwzP68ejaAMFeIR6nPmjbChx3r/iaTtMPMWM5H
eVCaB9gj002DulANq8CQtSjt7f5s82vyZ7N6sqVQ93JALxHkrsHtk5HGI0uFgCJH
U3I8oTrlQ83XrL/KleGUcni3rY7E5Pn1ndNUFHwDvX7mhcNvxAJbb94qoQcLiJd7
4+LuqcmhhLLRHCcKU0EzIKnAEJ5ifVXloa1UjefBJgsq85xUg8WgEAswu/IA5S1A
9rG3nCJtLOdxgqAzc9DdA04Uton3g0NgZGiwQjZilY9YAa18/deNUMXxOHWbnMyM
`protect END_PROTECTED
