`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQOQryEFj2qy+ASnzNKQf5ppahMdgHmP+j8dNwM6OqAlvEVriXhglD9urYCBBnGq
Td2nM0H14cgBGHyoPjVUk9qFhwGPp6gOXzG1RPaF9lMUcZCh0piJOZ/jDbWUISJ9
WVLtbdheMOtHtp6qVEwX5Bi9245QjhAS+SkbSG/TK7ZWeIpak9vQ5RcZbWpFGnm3
VVyg5JYT7te2zfuC4yHxFSUvX/l/+OFr7KfpdEdjdtSl9XY4GzE7pOeGMLdOW9Dr
M6wZpm7Bv8pK1Y8MlTbOc2ZDyAfjFckGNPxcbqTRZ+TCQWSyCVqQwFtMJSD1JRDD
r3JGeBIL4OUyXsEoc1xPhaWQ083WPO1UtGF36GAIJ4EYvFyU/7Z6NG3edeXgxuUL
Scx02i+J8iYIlE+/1P5de8pJd/zx955YOG5Jbo73LcLiMnWV77ZwncFPUC+bi1hh
pAnTDSrB8l7AOswtP8/mV3LXko+moUm9pL5/fI1BNNDf9KZCVOG0vcqp5L5/vGZD
Zv8C8nhPk9bSLsRmj6WiyABGS3Sqs2VCMVZMS4wdpmfSjH9AL8FAdCNsAMteWTwL
YCPGjCT/Pt8wESQyAeJnz0TCgvkdCgLsf0ErsIhtiFW9l1ulW0qVD2QU7u0ZhjKU
/S3c2LatftHiYdRWmZWR3+VdG6mKX9VjvaKbwsSmVCAp9xG5uccgAtmUUq0GP9Du
WvflySlQAtHpsHoMIqP3DzVOZDrkQdLVTf1XZTlOlomWrV2/PMm/HwLqjX0HL0ye
PAUwmXx7AWZE6CNTjzoNvTG3ieTPSVHUGk1K2pXTLlHznBMBmRWDqB6gCas7g2Fl
3g7bnyrOd0TZj1Axq08lnTgRBuVgxnw8X2fkFzSofW6xzLXQxXXMe5jAXnjw1fKF
CRFk4pBH9LHOqA2xXJdCHMDt3nUXGdI37SkTRsbbXWn3mvDY/5pj0K5yPzFVNf3v
RDH8rUiNx7oRWgehame+Iy3eaGz/bOiM+22BTp18UBiPapUPNTiULhNJKIlOu1bV
id+8Z97e6j8BCy1ERmuKYFWXaU1ZuJpTOmkTc7bAdXnDkEGcrVRItEMlOmV3Axm6
/mJPjPojMuzvVShE+hp0dDVHCQy9qQ3qv6V+pvPpyKWjFL7pG3nUaJ/S4BokmAba
H2vZ/GxKq107b99wUU/JClfapefEjEo4MpO3M4qHORXE9bJ4gWbgBee5jrEpkD/j
wCVA7UnNfkKqPZCKBp3qVFRemnT8x4sn4J3nGzqHfPKrXeRa73pAeggCfsYhv4u+
AiaNRWWYs+T0QZvYgYh1yQJD/4zu4/WY6sqgXfUgJDiNvwm0n/rpCNj2+YBX29Q7
bwOb1R2UXXMFRe63U42pDQteKYZ0s6BrbZIV4/sHEFmL/ogHK5Y7aSz2Kc0OJ0Gy
iVXhJ6b2OjutLtUVTlRqCI2atldVsNklYFFPjEJH3yKTMk8rRaVHRBs1qsQ8PsQn
YLyqKTQUIVbMlPa+7MM9YSF1hWfoRCl/w0LomsOs0Oh3vBEEweQiZ2cUdjHTFwd0
G6hxXFUltHIUuM4V/CpXcv/GjQBT8FX+adlOYABnnvTGZezcISpTQtxfLP+nvMiH
O6NT1qkDarKX7wtfuEER+1BPDP32pwh3rJAJ5bl4uQIMbd9XgqHmqj9Jk8l6HA5c
JDXQLm83HKjgofYMcPVVu5RNLlmrr25z3zgIBuHc9bbe4d+GJlH3XQHQa+ER9VkR
kGTQa9L5QQ4xD9+4E5RMLIlHNYnuzmGkkUi2T157ichiNN2cr13vscv+3GRoeJYu
WuVY8kf9qMe7Nn+CBlmkoKu26Z/WPxFbM1x2kUtQ1iRw/LZV3ePRMaYi7NX/iKLW
MkJxAmQDsBXkZCncOlxAPXkiZb21CbvcaJzinym2aV+hnVZkD/f2W2CW9zc8K4Ee
sBzGVlbLtpLGPZ3rQTZEBF76P2KZXKrZ60wHGcpZtkp93CNss3Rf9YxIkTyJ5mlO
rR+TspJ0TED9yvfCYyq1kjBxDp0Bo92NpN12fWq9PkM/lTeEiCXtk3K7vIvf/YX8
LlDN0+cMQkOtO7RffR1hXA3wRsuFoCOtoTM7gp9ZCuvpFRJxJpVT41CDBdeil0mm
YQYbM6OzvWZNmED30JYl96Wmz66D7GCc36T4F4EFlponb9Z5xX8BMI+/+dS7p7jt
97i6v9EaU+ms93ZvMNWHrv2esPho1/PktVCVQzMAe/rkn/BZEjWTuG3jZLmSxEUr
hryZrmW6aBsBccXvPF51Tw0W9y6qUbXXKdi1g4mPy1fmYiJCBUA57P7MMHPraxe/
FkeKdB+dAgVyv3Ba1IHRs7TDmVocTb0URg6N6+Xt1pGR4iS8G8fGs8WU1OOJ4Bwu
Ivc+LrW2srwzii4oZse+JFf1yzSRUp+5YpL0/r6llwYw0bLo099Eag9DdnRWk0+s
BV1JqGoTmR506aMtlJsM9I16gxVxpv+s4d8+hhuOjEpVANrt3rmOMxa5xZZq0uSm
MUGw7s8kcn8M1qIGdwjLHmZydbAsaLIfPWYcVFo7duBfoscVOYkfAMHVBqdOayWH
YbUNp+IHLiMFwdlrCo4YWrkigqApCBT2aFqaatZ0T6yAXKelWIjExElCGrWfnEBg
+eRxDs9XmBOakSXKSjRPJW1st7LkPp+p17BY9Sy3ayBUqGc8eUv90N4B1HIrd4DS
9X6B1wh4imSlzSj+w/32fvOjozMNeFP9NUSIoO/iBFX5Wpz9cUaW6SbUjo6WpBJx
RZJXM6V97DEPBiTbrFfPetiQllD4LIgeeO1eoW9DHBdzJqJIX+uWxCnmOkpTfGBL
mLKJyYL7kZwvt9wBQr07SrFwftlB5bAF95PdC00Cg3XB8L3gaVMESp0StrDrIrxb
B3M0p9VgHS8201+OM9+FjGOHWN2Lqnz9hNmyxsSateYdtJcpZBYA1/wgWnkabetR
kaFbhniXrAk6oonlRJuUQN3LJXhY42giGvkte9hSZmulX+gjBSZZSt9ThgZ2D4qQ
Ak1WfJBaR/i54iR6rBIQwVOi+smhqJZATrlBI1u4qs/2/4X4WOI2ZOxnHW0R1CSr
RV5b685Y1h47bi/k/MaMLfQHA/eyff3oDBa4FrSqCoGTYqx2YyD2ba5aeRAbVR7g
UKX7jzJiaXBo0Nk0ODFrghQMo0C2+hAQrMMQBV9jQQqkPFPMc56DAaUYUJQe/WFq
W0oKBNL/lGaishe7KDSiuowlolpg3DUSKSbZ8EsMgei19zwQ6imibogmoMlB6V1S
dXwir6/A/PZM7MBaqWko+Z2MtFsvl/8PEQDGvocxJ7noR0Fuqc/N2m6otdCWZ1aJ
HOaY5H6nc5sL+YbDBVScejpTHHszxKyQ3DNrAEkamNZeRfIBIw32TgqFLvNYX5G1
b/ExmYYPH9QUrV4cHxYhpZ2/N+w5WiCnF9SXsQwVUyRQFB651CYxvFWEb6iHafjs
/c8Ii6JDLFlvj6YqO8pjbIA8EJLrEdvZuMDZFM5Wd24ynYaVWXBPsnXta7mn6S1H
ale0DnNweqtlZ2p0K5Ln0t8p0qs5jmN1oCrXBfsh0fE9RBxjhNvJrk8AbjOv3Tfc
2jnJRrx7wVzBtdKzf0HPXE4p0WywUnuYqMHAD3oURDvQOuAmiSsEfg5NueXTE2tm
cRGKbOA67pkX7afjofwIKFhoDV7HefS1T8UzoJkrKBV9Ac9nE5UZnf1M+eCB7Cvh
XPcvYOp3R6f3xT3BsoaT8NHOWfIXKAFISHZuuIpTDOYgtCRuaIHH/WKs6bLnGw90
WctHNrmo/AXOtiix1j10cG1IgyINgdb2fkGthxfqR1oavX8msVjuZPLino/S6HZD
dwakNUhViWfJvaTy83eMSJeyay9mc5UfbmtSJebDUBVb+YRM/lWN2jJaXrElg1dC
7Ic27GfPuFDQk/pNPKLQ/cfEGiVBPy4OaFYGU2p9SncsPkzJlubSZEsH+rYxqxaS
S1HQ39OH0FKX3Qq0RvDoB6csE3FfWigDCvU26N8JfMrBdCeQajpnU3zxRE1XjWiu
LCs9ycXL79qBkuvlmpqYLpeIGMF3ie8WM/OEsiS8LvJ2BbW05SDUuchrsOgo30Xx
n7KMQvmFLygfWPUNKfNfsmn8G9gGqYB+//VLc1U1LEGyQZ+n4N3duoDtKeks+QF7
vv6WVbmUNTjriaUMGfq18QueIVGDCEJG00UrSWYuPv3uC1ew49xWubFk6pHEKx00
nEqbIzBjhh0sHUnNg7ti+eTN8dg5BFSDX2cNxUSWeJwXr3jKZ1gYrV9QhIXHXSOn
XIxIkHScSdJdtB+T0AIpKiO6TQQS0Ghb+twO6Efb4wywcuwlwR9UrZNPvrjzkG7o
hDl0p0xUTuURrkVOaMCOzV5MlU31lnz8VaKasBmvu351wqVhdA1TlJiQISv7YMxx
p8KgASBgrT+FXBquXxjxxXVvoORilzScvfXZhHV5JsJEUSOWZSXatAaRJSHA5R2M
VHMUHp7U0lWpqxSWQ/yV22m8HeopUiAWFIPwAzfHT9V9Ts5jIBcVE1SPArOcbdrk
gsaKoSdvAj7LbH02L6FymecpOCgxZkDq0cy3fwupblACXvcYnTm/68jJiXmdx071
VmiwE9FnNjdDdU0NToNNmEphOLYa6TsyHSV0YMMxwFzcwVbNGH7DP2LFFj5fDRoT
lfhHNdbuJK8foQQS9UqcMJcexpiQDpzBUK43lrcA9ZDCEihQCFSImFhIOqf9NvfR
x2Oy+6lvyeDR1GDOarn3ii4Rqozg2kEr7OOqhhgV9RkKsizlYYJWaSr/gUxsAs5C
dFUMzibSPQolPDSH8Le7TxnRRhEbDjs+pPmWFf/gZMBgi6b6w1mAii5yn/oz7GW3
qJMSrQFUbaKAb2Esl6unqy1T64pXJD42W8gNOhtqT0QcvxANnWgBMbl6QZWvTTi5
2HPB4OxPEiIOdqRl4S11Siw/jH6oZDUeFXKAFRddhGYoIdwpPCl5jAi8qCIkimGD
ZB6V9S/bo9XwUt8bDUraZM/gTLQfIb9Cg2Es+nleee1+1N46fPr2iybH/2KWoOAK
nARGYjr+gBPscT720W0jPPB9451vC0dzJyOs26qaKi7HBSwCKl47Z2jGPHhCFAnv
`protect END_PROTECTED
