`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxaaf+ohDTyUbzEx2CxHypbNfPy+9yNSBMyhxV0NpaATlKRKrXf5GmA7VCVyddhE
PBxw5lz6hx26Mwcfsmv8EDVMcXP/6RGZJZapGbXmdf0fVBM9o6j+IqS5mYBHLYv+
yJnJJ71j3aXt36LplQGd3+uQLcCVl5Mve2gjxQpBh7RV/e6JFpkIGBMLyQ7Pf/I2
CNMu9xpmllG+PoSJ+ZHJIUzLuNfDRM9ra/ehhPRbui2e+VPlUHRA8G/sMZgWJjUh
x4E+OI0Sovasz79i38S9UgmH2K0KgGTgbvCb9PbzRpVHmkm6TYp8XuHa6dJX47+n
TE79Quo64iNu2vJNiMYniLHxXlxrCMEgfMoOGdXx+XiNFqLbQjmRzb+RodCaT3UC
VUkT5cMBcmxXeljNuDKH8edOtVxDxrqrT8RKpPKPtyxxRRxC18gs0VS+OzaULUmB
+IWxGpi5Qh27ByfHVgKA4VnGcVm7KtQjlP+KhUj3xv4H6tjhIPfGUlFbQGlRGk1x
g/r5TRBv0W20cj2bWrpeydc1IRQuhNdGtPqkgAEiWkgjubeRsSI2JHeyo0Qkqo+a
LPjvW3K5LowFc3nIroSFbrfmida0GjlWLRaCuktfvgzfldy0BZyVqKGPMoFHOG41
uexzruMuHdvhOfi2TLaz04nbPsNDzoL67Dhga+Rnkmky2tnKiLg1hb7+K6qn/ei/
MT0uKucVHBZLylXIF6PwU+1WNvl7Jyisg/8CpL/zlzET5qMFEKtGwf2WY98ihk21
8rLKYT4Qb0cZHH0iKvhVHdLaXmNbq1KrREUkA3M9eveB3+Czb9y3IGGxsFewik3Y
OA4NWZBdiM6YU4WZahQlLmqP6k79msHwKgp+qyZd+0OF+uJUMPNxDWDAOuON76ND
3Xg2zkfv2d+TrVsrKY612WIwHwp+NbomDqXj52IzKkdEtQLvQqhVHDP4NVw/lnHh
ecIB7C58apWwBETEqy+NkGFJDU35vtddWroLSDFmSF7jRI+TTQgYcJ5xmmMVjEzi
XiwcgeTTqeP8rApHmHuUEyimAXxQwGA+TlQZzb+gaTS7I7TQ7Ln/DXFV7kmzXTuB
9pxtb5bnjNNhmrcmQYNMcwA+GDwSCrxZgEzdRZJEezneh9gDw+XTq0iZsbM8NAKB
6kwcNHtkoP/PnI4Uokr16EslZ6v93fhlBMwSK5pxEiv0QzT5Eo78rk/61kV4ALIW
oF6G3hHbwKNhG16yWT6NLmvoVgRlduYAT75MObtBSvE1sgX7NHY+6r0s7OLrfImh
W5Mm98TLiYWwu0URepvUq4yefYOrjHhT9CoCgpUWX/OydvXgUhWRMDPYzIMdhIQc
DNtG6U5LCye65eOsETUsbp4xzh4nnELgOMHArVIKFLleGTRmtZlgG7l/ISY0ZA+R
2pTGLtcng2Ne64UIHcI3NhasX1K3RwpzUkHkRKdDuDs3trh1RxxGAIp8EaAu0xHg
LCpbIr/dVngfPXOiNSjy23PyqZAXWKmbbtySTWjd3TkJfB3kEXz2UWHLA2/wYinW
zQeHV9csMlCFqjUjihSGkIVeTnBbeQdVGDE1BM7WrvP7XZY5R20Sgld8D0Vf9Xx0
38u9VhHMMWcGyjxcyuOh15U8iHwkoGrIfsQgeFDiHAB0fg36LaYeP8DydZDQow7f
XzI1SdAsF5zClfcstAYx5bfI/NtQHoi6SBD8VkOiMSTQf8IHzd/pcyPZ35hxX0AJ
NxJ/59OW+5W4VOiz/uQDAgJG5lwWvY6Yw9aoKm/iFLxQN6qYaDi7lEGoDqvhpyp0
JQzS2Is1uB92p8/ucuqAahUXjwem+0ZKh35SDSEJBjAh1kxNLXyKQ3EFbzLgPj8q
MjBu5C8HjcuMxoRRyrC05T8Dy7c85ZG9felfcPJeuwg2VL64NwTi1vN+TzoWTywa
sMHOK6TiJ2tT8XqgDMhovXBtw7JaUI46esQ5ki0HsV+1Dxha7rLkxLMgLBxxvKTC
vGzLGHfSYdcZ6uTP3Cq0q6bF3iBxnRr+EkF7szHppzaux+aEzIj461Tdpj9clrQy
9nzLi8wY5kGClv174KTZlNffo3MDHnheyrjcbNCOZvOVHCFkodUeCM2UPlIbKKKu
uU8Yak4j79NvD3rWPFMVzp8OSsqcWfF6/VZjXkvCraI2kkFGwnv4/Fl8hWFTWg+3
kh9wHG5RHQDQPWdOf2GSGs7vBOdOkT0cCrpozEz6YH9QcWvHBeqEPshnuQq73JdO
TGx1HpHMn+rO+k3mGps+k/Yw2H8kf+BnhpDX0DfQ+VcETtkN3qmbR5mVEkQEp2Fi
3minjRH/EuUdSm1JRKKgrvbJToRrkgGqKOGgkgXExM5e75EFQhtY6xO/2csenfun
hwOp3gei7wLHrzTPDOOofuI/N0jjZr/Z30nqeZ/nkt5Q4SjV1fjy8LrpKy512Gxf
I1OsXT33ieEJUpUHuf0sCqsDCrYwKGS5im/4El+a2F5ygaPK613J9Be0tblSeBoz
hgTvIkSTdC5fXwqOigVRx9p+ZMf5AKNYVViFYnOauahYiBRmeDnT+fj/weI6zDXm
Q5pj7bf19mQEctRauJHJE9rtwwz1ELTMgSZ7CnXExwckWsV8HE+6yhyr1owOkX5T
auFc41HUyTDk3YwTa1oUqp+9yMWbneSgUc31AIEe9OP+1eH/ZmcV22NpHMYV8xU0
qS7Yvj5mlHDqtwROB4Zx5ztFssDwOuIHlwhRG8WfMQBvNIEvrPoJ2Pndkd63I+7u
9SN1cDlwcqPVgEagiiIUfbRXLiQHbs3HIXVfhP5Rm1D/gFNc9o7fO8hJ4otB42LV
+EqOnGOt5hOVyjj2nHP5fkpBcWlQH5xB59GzL2kaCnjcZzmMt3OA6zqFkvJ8dSpd
vdus/2EvMKAltPqyelTxqWXjiFn5kV827L1tgE8wU7ug/nSlJ8maog6ltaDpU3ZC
+Pf0V9tM6lZLiMsA9LEGSIQIs02UKeFVTSvwhN9rV+EPlDIoy03yMJ2guWiJ4s0p
iVC4t9fdZIpxRcsHrpqSfyYwqoO9H7Uyi/IGnkj+bBlC0fyL+Ulx1VEellVdNJXq
rcC7VqmduIaevb37XBafAKp+EtfJKrW56ODRms7rE5mAekPoW6pqn8Jij2RO3CIu
PobnoeZFy3pnJML5FdtrBXM2aW3KjXpUnBJsaje3Kt51NRi0wdPk83j1s0SzpLYp
iNJSCHGdHMyBarJeeXPXStHkujHbl30aCADwaDf5KAZOIW1NV15iGiuCJmNHB0lS
rxmH60qPD1IKH3/apAfUy9BOV0Fk7VAn2qz6akSS1wNz8d0wXIwRV6sCf/21ahmO
yP3lkENp6V1ITvGrVX77CJYzDv5tiogofzGobt9LmKzxG8ZTJ8PWrzQW9u0I10Tt
8cGWjX8TL720P/NO4mR1GERA8CuS++ghm12jm4blqlg0gjnUlYFBNoa/glRBY2Po
qO54erMDSycl4lEt99Q3Rt3KXS2gCKGXqtA0a757OyOj3/uXBt28/ZEgBp+FsW7e
8aXWB54I8hkg6GLt5+/Uw7wmBh0ykUTp2YtuuHCOGT9Wdvfc5i6WnSgXy9He6uzq
tnJtJRIXkZWZedP5swvZUG8ZkhLVdJ/Or4xPY5slsg+4VS+73y6rj0b0/IayQVqr
2zM4skVIQx3nDeb+PBRd5aO19Ilgwm6QZ6WTKSgCA3XX1bVn1neKwLAUmnDFNoUO
f7Y3uV2JnflP1DDfTJIcxREmDWTBvDBCSYt6l4xSU+S/HDTDTCSqUoZE94xT+n31
kW5UnawwNeXSa4VMZzlPEv+e3gjyr+F4VzDUxv+wpcYtupf000kK7sg4JmPDKE1R
y8ncpQzIIfyaoVtGshWR8uFKdh1WMFFGpMz+dlgmyAmKSDHhNlo84DQIpuo7iP8u
uQAPDQrYO5e2IYxxAY/ofGwJStteQf5491s7OSrPMtGmxz53Aeo12rXiSVt0VVTT
PTptZVCjavoG29T0gjdyzLqO+w05uiOdo/2vIePqrdkNCbrhlTaqn/TzM5YlbuC3
MQaRISQvqx1Gcb/NQHa+m1j/n+zBkZJSwWCx5B8Gslm8txNtpqgCWk8A4LydZLan
nct+LVEHBkLzKoSxVBK8YzcKvQ3A+5DDyzPv04UUZpsfBGxns1fRfT49P0t65arV
X4XImC15kwznWW+qqPXi4Y34koWIgz/6AG46wzFYzSTBe0cobgjHxrNYZIqAqepH
b9KdhcwPU4zTxWyHEbmmccodvHGs1SgWvSL6+qnI+vlBuWz2p20JzipGzEBVka+u
dxYny52ouTE6t4UEAx859PQRR6E75oCyrops9jp+AlPvjA1yo9SBGTgaRdE0h73a
VFLSYyrfi627L2yucHY0iVQ2QgAS8HWK/wNfRPNKAG7DRiFF+cARM2cOj3NGwpde
T7lukcsiWpi5NKu2zaS6O9Dq8WkmfvNvU6W20vVMbFFNVFsT5HAmf4QvhQoiQXWz
0aTRL4Vw21+nGlCJhuoyToN3jxc+3bMN0Wm+H0qHBVJ9IzY09oyYABOn/jJtorhF
MZBbTDwDwEGV5G0hbr9GzUO/TjDnNDIWaG8B8nF9f830LBpujyuJiLS1bLYq/ZS2
8VWIm8usR94ooroDW8CyTB2rxeduazGXKDrEz1/nPoou7LuhUViiV6bK8Q3vP+xt
ZPyzKtwLV5Xgx86xgaYYmu79/EmdgvqqUvsagn5De3aSHCxSmE1svCtgCYnE2ilQ
Xc9cm/IARq2idg7eTQm1JEKzITk+JKOTQjZ1/Yy0tMu/VkczGXtfAcXb6oStkuu+
vH6H40XCVWKaNJf++vgC3peapENun4dv0cj8QHrZzuvwRVK84xhZhilCqJoL/6Ew
Z16mdoxTNwI7IYZFP7GsVoxCCI37MGDgW2cqojmlfQwXxGrv5UBMd1t2qJk4bB68
VBoMGsJQoRL0lV87uAfAmLHYhuoq23Vmc+5hSjK/iq2nvweSET6LAzJN6Of6ue/i
VWqNw82Ks9FguBRbHuZgROkTUPpC8lpg/rS2sCvzSasm7BOxDAekg7kDliJWhrqp
TKfjnti1EQXvvjoTgsCIBHSVkwPg77veOwP65FLY/5T4jCU7rP22zQxrkAlfzUrb
+pd/H0oltKmvQ+OOAgARkKNmENS1KApljsOeYtlDst+S768tZj7I9wR/MwDle/Ql
sL6Glx1pXKkmplcP1JCaaNcLmdMQPALkxhCuvSt+FS6yxn2HMnZU0ORDFhFtNhvM
OWmK/+/Nr9YuBLSkwNbX3JIh0ufBoRooKc7pA7bNucBaweAeA2RfDZ5Iua5gDefm
7xd6qwXzNAB8esHe2thQi2R5xogJPxbWIFSeWu21KKTBqnggBQ/1naim3yRYMSFf
NnGDYTaz/oEXu7MrwcIEO7JKyYBSgZ7Tx4z2psRtUyKkFkDvW9kPacDAJn6K199Q
Ac5ibflwWRu0SIqXL8r5Exxr6CR2wxu2V5JS5MLGP+21iAhqhSwg2VG4nPseg1pl
/Jo5AZL+4M/2Qiu28iPspX5EmEcmrQcoi7MLbau1oPMoTwgQvP5BAuI9QpPoLm85
lqzxIehC5Zjxai7q/L1GNplxZOyVmRyD1hjAyU9QUEokKnBEkXKDrYHFDu4LS6W8
f7D0dYAdgcOzbj9ATyeft/AfkYQUNiTCY22/9qxzfWG/o6kBNcry4J8iRGKMipPh
Oq+pC0gFIuuQUfMhyvAlBSi33aS3nerNQjaUeeZrx6CHR/GNYj/lzCkfXq9BFRH2
7L8Dmy+/WWVlAk4YcHGQ6q2ZJ5m92LrPrdOe9CBwc6P+dHzUrQRRtXeCsLKty4n7
m0dBrO6wd6c4gMeY1BOtRAMFhBZhOfxUiasf9MzlkenUlURnOjpQKnHSYfwETECz
mC52NalpGIyFtayngU9nKgEfXAVdDMkbPSWrmmZlZ2QVRyNRLFTaUbhlJJqcFfwn
XWB/u8Rz32ZByl9BPSIfQGmQ8mUkQs1VrsbSobvLi6t5YhGkLPETbi/+4Ih4a6y/
lp0hc47O6tZXfdXphDE1v2wvTo5Zuy+CK5sCmuRh3lYRuR3buZSMxzW4viROHAsr
6aIkvrPS7dvdJgKmaOQhqPoYvWoi59WmvGtKLtXV00+NzIg16duSH5awGNaxhF6w
Uk6iDXZDvve0UyQqIjd0DAlCOjQRExHt7Fh/JQBf3LffUj3APJBAR1xr8MdUI7Xc
zqvMNNpx6j/q4LwnFpoEkFBwblumRV48VINS9TS942LQh1PaRC838gzJSqmMSe/8
yDE19MejfWhXAC8cjyc7gW3diSEA4w5hRjxcQjhmw3xs8wOWe9M4xTo3tMCWj+MD
AlEeJ8Yta/WjAsrN8C3T6AeC+Z6rtFr473sqsCXYvqyxuvbKw7LL2sE0La/J9qqg
D2P8pv7GCxSGn/bYgSJNxPRZDGOwDr9Zm8VOh9mgXj5vGzDMU400peg0iTIY2xvO
lTL6D1U1vkUM/G1WtnXdhdo2Wv/BQrUU7lNnq7DpQ+X1LiCOnBFNBG7gicKGu1VE
1oMCgpKgUY8NK8aqYvZ3i7vOSHey/NCfef0oRLASLEpeWoDveFwAwskLB3k95Pes
qd66X9cs6UqouJxQ9oPFTOn4Y/ze4zkSG2N8aUArxF76i1IFbvDezMMt+O86m+Ht
`protect END_PROTECTED
