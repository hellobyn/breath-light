`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PsHOfHD3xYiZEsUGe6HQu8M1XWQvs5d01daYNVcoNfnQzl/pWLPt2Vi9cBL6trEN
xJtqUxlVbNZczYu6Cc7R8L2v5Uk0JhMacCX4FUI9PFW3gIDLhFqGaGI/Pb0agHNa
ira+UV0uYfrLgDs3u9LcG/TMt3VCX/MJzH3ILsnZtpO42+VnIdoEjWYFqrBW8F7f
Y9QjIAzHcnTBct+nj8734epLgGn0afEehZ56kz7d6r38WqLzOuF6EAbjv6yGEIT1
cua+OYxERTmst+Ttl28hT1dlF4PdbWmcbMeWj+fVc2TLD7eBrebvFzbGsKtvAvrP
cFM4zbfqA9QCTI3AU7wykLD4Oufq7c3Tu/m/1K60Sp8GSyQIo6kPUW7hDrW2iKC8
oL2BQb959/uqfIrOs1gChax85uET/qjqCNW4o4Uz/YSNcfTc2r0NTLZiSjPeLPg1
bdMOQ/R95d88dPOg61aXlsTMk0OY1yk7in7fOLB+WTSsUGY0S8eCcDUI6feZRaF1
sjHnQscB/RkNvn704uX6/RHQTrdQqoePMebQxbOBoqtmINkvsZKQ1z2UiNSCUExu
KrkVLr4JKGHlVJusS2Bgqoy2DnyYzIKpY2qETBAVSDtzOVb+8rdw8h01CsNeqWGi
Bne2Ck+2Ic3qjFTJgE1ngGS0u6ZjebufdjkxU2Muh2jllhMrKy6K07MIymbITj8G
`protect END_PROTECTED
