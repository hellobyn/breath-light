`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0x80aGm3oljyZDSyA7T6H03MvOnnFEeIxb46C9L/B0EL3Dun2iT45oCJtzJrbfo
8c7TMBozvRN3jn7ypaoRdogPjMDhol3UVw1JVtQd82QJ/3q8czQdWn0PrGYSjAP0
71VQ1v6pQ0bXPo91l7ovX6ZdwIaoscntQuglzM4SZz9Yda16jRohCWPvu/6CHlND
GEQxq91ySyG1XXkREtbn4lnmCSkboQV9x4kA4XszBxZZn9A2GFKPf3gCk6Vg45v3
AifxiiiOXSAqlxNiT1N5Kh9fmv9aPaqMSCT3R3vsXT1Lkp9rJwAr9EbEb3xa3N0W
K6ZdNrDvb1yWbnXdMyWP+rWxdNTncMLamLh99VIFLeHC9Pctff5bT4WbJ4w79ud+
P5IjecQaq6HHNdmQzOqcQw7hBSrrNbjnaM/2J9UlvQ2LdejTderO1slnJiJ5hXIy
w63WMlxBr/h04AFVcJOzKZ7yJMQ2jnGEQRuWeELbaNSkRGTcLJEsyT5OzWpvBrbC
6xrwz0H17qsTDezGWnqNa1+fFSUW8Sf+jrEn9evmWbueuvOZc67sKktEIaJ4jvX4
OsiXl80ObKZEkyUPulmMM2kLO09VhPB/rLJcQ/CibFbRMFe7+LK51q9LwjMYjIjT
BO0PIj9/rXiakowul1a2Jpe3wpU+QrKcR99dacJfyPkrnqRl7Z9IuKvmPkXuvXiO
8BQcp6sY/nRJ3YX7NpfWOVxh+CGDvvN7uf84uDxkLLSsFMzy81fmDPNvKpABp8h4
pRPztFn1faGG1l3VomWy61WbjzbLwiEn6e4LM3MN7KqIQu9zFSUsiGZgmHgP3ofS
IUsNrOfOK4PO33W1tlcigruz2YDDFa+SCBoqkIjPRMC2VXTj/9oOHwVik8C1rPK9
fHCeTHPW/LbaeSqqY74ifTptEo8CLlC2jcoCK3OO58EFHIUk9qhBBOg9xcXP5KJc
D4T+GnpialBej4GrBK5vMesSug6mxkhek8EPEsa5Kb07QgzdpqnXN9fJVjeMSd0k
5/hfgUzyqm95eN/uckmz1Q0Ca5Z1561TvOcJ2bFxlYuIPQmGQ7WvOr3mEkHwJb3l
M2xY0bmOFeih9yAebrJ4u1JJZMglb6DNQjqCgZxPtVSds62kNVTuP6CYq+T55dsL
4g9lVMHIGe+1i0tG+90BgOw6mfm67V7oavaofUOQD5GLhqF/EK9zt6h1vKhYvAAJ
mDwR4H/Y7qXtZEgckx14en6+qF2vfGWEo+3RLU5OJFCeziB6m0I46a1EJXc8yTOG
+RKfDd6S37FAhB98ahD76oPSoJHAAdr6o3zQTcAbbQCCytKNtd7Y/JYuPMBU2DUT
1OXEdjgGY764nk+lGAzTcdiSFuiBtFyZZyjFaJkj7TCbHaYduhCWxYKbm9jk34J1
IMatfgVad7MLP1VH1709YOfiFw1bV6gyx0xx4A6TRGSFejbF5/uV6OIehmyBqxb5
r02fzE2kEyEZgZjWQB+HnyMOmS8DNiAWwPU1icwr4AYzzp1SZ7uanONVFIcxqfK1
jbrQ9G61j8JpD5K9HflLdbmgxcKfcZ0q2ZBv6lk/EPFif3qH1VNQUtmNPkX7zFr6
Xn75RmMatLUhapRfx5FP/xUiGehYCe6UpI+0kK9xW1RSufhmEQ43ZBH6LHq7l4ts
uLzi02VXKyxtFnJ4bEuaQlfl/zv7uMKNacjaMDGvTv8k3LQ86JvctpdqWLvRXPo+
4/WYIPL93o/W1p1l9+4NI1qPgvt5GYtrUfQ3Fk7TsouEBWTGGRcwRoY6fnixi2pj
7CpqxmipR2U11lhr4Fter88WWdoxSdEPTAunppUEV3rKEytqMZoT5RW1VX94ZehP
r0oIPkrr5vXiPygUcFqD00i987uazV0UTiIIw/oFMbVeFM8/rx68o/TvyJ9Py0Y1
rDsruy9e8vzTG8I7u98X+enMNPrrVv8Th4/6Ht2+bs7jPdHoC5D1zEZo1+9+tzyG
FxsDTdMWTKbUp10AQ1PhFC3Did9KToOUuLo8rRC5ULKDUVLBXckpjbk9H8Mvxd+m
skN9r8Dj2SDgZv8qmGQodUcj48NeVKWcqHiVjFNWg8EaNaXfjIPz3ZJXJpzUO7cj
Dnx4/QeqZTSNo331r342zb5kbyKk+8+x2niH22kzw9uheg8JoGfrE0GU6Skb58Dn
IGMBwIeY/34TJ5Run+fpKQdwHJZUK9KymT2ao5aImF9R0qhWrPbBwB+/3ovRk0JO
xONGW8dOU/GDzab7WiRuZJrDZe9v0EYk7xZhEeMEO8H3X6BMARkRiLbfS6419Nxx
CoC+LDsk389JV4n0IuOnOusOv5Woi+v4lkuGH/HLVqOChIFJCcvuDIiCrfBUi9WM
ygdD3ttWggV2OX0n7mEtOoJFy5GnXGDPKda3PPuWSBfApUGE+amtewEPUl+sUTlZ
SH6H+aRdkA8mW7IQvFqUs6Tthc4ZuDlIhL+IWM1QclF2bCIO1CtEGDNl3/W4QBjH
dolhCV9owSDm8nlYn7mNwr7mTm7LkZtufbKMundxNxrltddLCWvkuKN1CdpQSZJX
2/sxUUsBSRI9yFw3tl99xRogp2ncuewO2iqwQxUlntYgCTO7weucLphrCejA85fn
g8ZCDuYyOwgInTX5R8aWVWZr2KRulCjI7SRdQjBYWZMkn1gdubWMo75rdWTZFZL7
YjBbpHtYsKgmy9Bf7vExTIOjJZcPfnpcmHbWk31lKfKYGRccw1corJbM2ECi35A/
Sga1UhcQTTzOoHuYVm9RGhIJ9Ns8eJLiYJkocSsfoFF8KSyuyCDWKSKg/dRYkIa5
BuGzPfPFtrklA1nvzzUng9VwZ2dUNk+pOoywzTRZHW7DubvWIisHhw9PTXPMG3G6
T2oeWGj259eR7HDExdfHaMX8xG3bAKuKhBYRhvRRSf8t27PxPakOpI4vh+3ef7SC
IrWXsZoWLkhOSjSjSWEnQK/2ZOgMpeMLDt7me3HuyHt4Y2QATDezKxZawLZqbFJ9
Wtnku3VMWUYI13j562nyazd1ZFjsr9grJX7WTx+JOSNw/Xw9qnTkmYxsKwH4NqJ4
s510EF7o0O6QnfAy2aVmYlQ4556ZNoOSTQCxtf/IHlQqCb1qwvXsrabf4v0rMRnV
k+tCUWocnbFYUJhJ5OvuOJ56SjOvVkiJ5O6T0wFllQ3HTC4SmeXN6qMh/qPfjCoE
zUuHwiPxFLyx+kUyF54KfTr/9VRPeAUOG+CoJbMBgpw5czuurKcmb3FGpOYnAiD9
APJJbAMfFQENIVVYpbJPnuZzk+uDU3tDToj5Zar9GSLNpRZ2DVz8c/HLfst1xmer
mZWNVymun+3OabskpZ2gv2XMOHjjR2YYqdPq+Vut/vWzf0fS335TAKOYwr2+kPaP
pIFQprfcZujZ1hhDAjfEiYtMn3sPOknCH1Xy+OM93wcK48/IAGqRMl0NLM/pyXRg
DS8qjvLbcEe6GbQQZahbc3kxvo20+efDB2pEY30Riki37mT1oh2hG26PCJcS4keW
LJlH89xydDXWT8G2bl25qFtfURhgOFCyekFtOSY1qzX7KEl8Q600KtgvyJilqPnv
+Iwh8+gN+zPnPoNYgl7YC1fWnUG1+Li6TFftu4+gRNxXqf+Y10iq+kjljj7L7M/o
cVKOY/yfnDdn7dBHF/9rkdFDNXnjuzkthlPDfQAplziLhhR43XEWUZJ2Q1KV67p9
1zJginKkquIojRt3x1AQVeFgcIyp41qH3yjpodDz7OcyQ991g4gdJDxYidIDdHqo
QypvfpKCzl0LEzHGkaTG2y6jvRbM70Ub10ZAL+y/oFH7jM4/RSCFYXU0/dJwIcYT
2GlQPqtNrML6xtNFHtGmvH5g8Tg/6TwzmTmGuwQUn9NKY44kk1QitSZcfPJvwEiG
ZcrKpZ3XP9+LKMxmWPYwWgSreII5gKvGQLVyhROGUtwbQkQHi1btO4e0iZly4kaM
wMC6M21fHXppyIwmoikZuDbBMnq3dRvDAC3iLW19tNUIqWC09dh+3WrjkfrWIgPl
uWSLCJe4u+KzhnH+Xh5O/U6ixfvfRFVL3kxYuHs05tiX5exLkeOzySNGR9QVnzoj
6xR4bF0+r94D/xRkPMvuK0V5c0RvIZonwQzhOTXI7oulfbdtLg/XLfAseyhTBW5U
8jUWZELCSgpHroZCjuBE4s1bpvjgBzGVIMeM+Qy8JbNFKl4+iUX6vwkdcFwAYj2K
vhlVbHPL5jwN1CY4UTqunpfPLfFyarAxi39RgiIJBdGjQbuvwcJcJzKpQgvUb8zO
yBvYH9z02PXoDDNhrgOA5rbuk+rZiBYOVXGdNwqc5kQu5Ve9wmclqqK7nAkBkuQU
lH0HWouCVXuNeI7u0IvhgznkKCnx5QSu/trc9Fw0bZcYyDnuXRdaZh7AyfxjaPpd
KPxxpzXUhbG8RKd9FJtisaakv2AkJYuTspNqiuz8tBUl/jyD5OqI9R5msrylEnPX
JjGLZQ9xfdFlvhRno6hYd1MekvFGg/+yfC7J6icnxvXqnymk2qZcjwHcR4mJo1Iy
uNC2JN0rptzbSlrqrIhjwu9nLXT+lWATi45yX6Y9XjhmJkr/FCsalQpkDSzL73vZ
FKspRyto9eu+J/2lRQK/tv4aTlbvl40WUOcpJF5i3wSRZgIVEjOXbRxO5zZwoRea
TdDVLXRv+nBo8Lp1jES/DgnHh4rC1oZQizb+FJK061aIfi6n2m5h2nVkO6oQPpCj
t/9AbLccVIYc9kbOiw+a4lSj5JuX34fp6T9PLZQ9xRVePpaC78KgduBr2jUfCNfv
3FwxtpAidTfob+CdDtgyFSuCSVSBewW3OEm5aIZfQv27JQlMr6apJ8dFgd8u6WCR
7FJKUhtijX6DGlnh0bBRpqILGZV80acCMjBWb4XiDdNO2p39wLDqPTtEv6rCdul7
iitw5VRgeubW0ADMxMU1Vqg8m/bdyR90uIJgZAd5/d2poemBLBYYtbhM3Eu9lshK
YkcoY3oQszy2irDVroiiVfekoksJQKlqVt7dPn78V+POigoqYflY1dUstXsZupu/
VKDHsFkgLsrHnbmqj/d0/U/GJm8Bc7Co1DJV5ISSOH8eQJlwYFtiJWi0Aa1/eQ5w
/r1/kKN8ECA89v5JQHLobYNcytyD0kRlMZcN1fmkKtNEO5IF/XNhhKje0DH8RUFY
uj6CklPbCyxOWH0nDl+reVie9eAvkVn9WmgkXqe9SRyjto5MzQJUEvtxt5N5Cr17
JMyKbFkecDgIsMlBnieXccPIdDhe1coz9Sy+AncW/e61/AHf/Ox4fwQw+pGwzCPM
WlccxJloYMdPEjvlVszo7GokR0K4py2V17BoMJ0WORx2KZAGhEYAmRB7FZkj+k6N
BscBqw2acCclBg5Bnb80M1Tr4TuwxOhB7YVR0oWVTt2SuqefIi+/eMoVs2Y+AASj
I1p5rbIiaZn9mvcmL/R1nNpdT13hLwRWWrJVpvSWcmbzChJ2BDiwiFbj+EeQHmX1
Z8CNhuwScNNlcH+HgHd606y7WRmgOuup9mzRVOb+gZ2PCV0PcUi77RbQtJbdLr6i
55RRxQIE1ehIIncaM6Y7heUGQJwaoI/01+D6RpAi39kgECFIpYMA42AyMItAOcCx
Kpguxeoqqy5VGEDVR3QOPmpPosEt43m+2xvcPF+emn1BRRmLlhCWmKFRKzOFPPCw
QOqqvNCiBmQX0birFcOIytT7c7dx+PHp6VvtRePMj8MKMXoWWv4tOt4dseh9YhBn
2q2Y6b6K0BkAqbgy+nx9f44QOoBKO11BEtsTouF8KEGu4LVrSZDsItshPH/N+yba
KN6FJPuqU7efYKzKb5kqgLUlbBr79FGRsThg7IEXEpHZSvHM1guPCOOTjdNI96gh
Tna6gFdwDR0Kgb1Erl1iWQsDBCEYgg9MW+b+MpMcPEes11gDRm1PdhxfHwjrftpB
`protect END_PROTECTED
