`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPVGMqW+P0KIvw1LqiTqCsejfy6nY9JsTUK+MVaaqLf/6H0thlCuP4ZaNQsiXFtt
+laqWz4IgRC8D0Aly34WkBe9UgVLQ8fT2lmMxaHZfXvtxqGEjKKEYKfUuUeRfJ1Z
Ik5eiot+I75ohvnX2SEQQlWVD3zdz/0yUbYqFORGjgLZZ+BF4A12aJP1eE5Kozmg
NLmBfnh3XvhPPPtC4fqMy+moTVKWNTQ/PzFtd+HXr+l4tq/FIaOAaeKfavZKdDLW
xCZeAy9EPRNilh2G+smLWbbCKtxb/HfEZ77pIjMOtvtXkIC1nkofZJG/tCOZcJUq
TZ9huCXJBUYJwNDvjjM46fbUsHZu75OJJJ8G8KdlK1DOtbvewsD1u4jxGzJM8Iei
PhlfEWILlP6TWvTkXTpMvpPICzBUfyoLHkM8bBX92ppRDid0mC1LXFTFGACIvGTq
NTRi7lEcYNomlEGY5h31i3hUeQy/tCphtz0IZ45+VAu1kM/3O31sp1YwfAMLCNKB
FnIqWrH2st6JET7dwpt42VUcqrCkMjfI4qdf/6XV5B2miFuHWJY6uzTXSPcJr0qC
0icFtG/cbhmTGLrp2YW8EZrdFU1lYPFXHYDbDAE/PYVGHqGBFG7l/8TGKBEkXXOm
bgZiYbA9dbAsyUPZpI40Hw==
`protect END_PROTECTED
