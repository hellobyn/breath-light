`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rDPHcwdUKg+AmJQK9h1YW1AzgweBsMP38qzf+WO+kiKs101exWbXQ61eZUD5VP39
QiYspSx+kiZaN1mdrEosgDFJIPnIK3aiz+gfLENCPMEr3iNezxb2+o+rVg6DiE4J
yuqQoh35myFSKr3bM541rw0qySe+cY7jd7UjT37x1iKB7pGTJMc7AGr5b7RsSkyC
5BT6+7Sgp4Z6qupslOwVt+31Gqr3tDijS05hmywiT9zTAqPcNVCLh5Ap49DgclWH
lKUWCEKrvHZCMM1qcoqfnmE/NGx7T1xeYygIx7I9srOwSNK/IgHmrl6WDWdwKBX9
2EGGset1zXqYF/pwqhlKsdA4X5TutWs/K/7fgS2eUUSKvdz5kqTCFFxArYdbAnag
LBRNbaNU2hOmt0nkqgxegg3tIsH/vlC+EcR0WgOnyI5k3r51M9bbQf1/Muw1bqzh
3DBnZiZkdZPmylUwxFI6sDHy5h4AXhs6ofj+dOmx/q9+8rmzVZVenIZtOzSZ+HNd
Ih0r56hmcyoU+/1a4mysdGaWA4Vwy+9RMUZF/+F3e6819NNlGINKIQ/8dM9LHae7
bbqFsAJv7ypTNpnB4Pczlcx/tKF12rXiYfJlqUfaKybv0VApzoKte0DvYtPPboVs
4+BBweLzLMIRrQsDJz/a9p21R9ZyTFa+k1kcwswk0XkzBVplPMiuiirliuAOVOSw
wUkI3AljAoGQlYhflhYglrw29ZUFK1zzF15DywQCBfIgXY6zmLrVbQZeTrC4fTpm
V/SL6jsPV+MNfEmHzxB93cXqhcsMF4rZYB7r0B0wZsSwjsJgVcGrJZcLDTrvBuaw
4DobTllWtiuLsNsTVXhrfawQYxXXNG0KovEA7mlwFD3dkBod12z908cwqalQgBZx
h+KYbu49RBrLP3F+IeHRWnaTfDas+UXFlfi/1FR95vDIfV/U8PesKG7fvVer3SXF
M37Z0A0dKRhABr7tQzuIRd3B4Ns2OOmYhlykQ3Ue4DmX4gpN5oHXLAiwIqyb02pJ
FXdo5HcDgfAitTf94DzZvMX+WQY+XmPBJmc+u2t26UfTJV1dKHpuN9sItJymClwm
zODmGVr1lFn0oD2puq9l1aRu8evXLILzU4RHyJFEtQsAWSBp4ZEwORVvtHNYJF+j
MBuflyQWIVHIkBKEWTosvZgUx+NOhvGDBxjIY0C9yBgWDTTNHSqbti8YcJ04xZqX
IDGT75Ko9fuxgJCjMwaXmwNcfSPxT5Cn6RxYIMdY65ZxWB3zv39VOAyO9EWoNFZ0
myVL/fo7V8+eeR4+kuih8y7rPoPrSWJjs6fHScb6jfVn4PSwjRvmKJ0ZDMm9lgeN
Ms1sQD+Ca7PfDyCDDWNLL1LchpPGINz0HYzDMLqPmF9egbsRHMSX50ES5kNHGb8t
tH55XYHApQTc6KodP1dWiaUW5ibGl6llTRgLAeBiJAF8AEA2FIqT2NyNLgg54Nwi
hK3fluzjWnDeylKMl47dTQVig1uSke/M3ONLQYscWQd63ctGmap5kc0VXGy9WxIr
GuwZmFPS5WpX/MQwMsgmyPLz1sMhpGAK1F6lC3mEHof3BDxD+XMsLt6iJCCwpJlP
IqhHTi2jLVcfkj8IyjURuUcNYcYilEeUlVnIkAvSWNbNtLnHeOcYHYXWYLb81BW4
XAWsdJxx6azhtClhL4aN9ie0RpLR4fKaXm3mNKgY5fh0zBWX7+2zz5fwDE2EUhhK
Hdq2UCBnnn4NBf1K/1RnyZs19NAciJVkbmHoAzpQKl3BwQzYodTXXLjbC7vl28ll
SWk6WOC31Y691UlZaR4JX5Htf+et3DoguT871LH9ecCY7XKb0fcbzQARPnZTi9cp
yi1450aelxRgs0ALa+ADf3d9geXu1Zo+WZepg/Xl8KLMpdovKIPrplThZ1drDy3i
Oa405wSDcq75E1A6992r2TWGIZ2ll5yWONU40UzfdoEgWAkpiyOmtAuZRa0wtTzx
5cpf2uN7v0Ak/69gMvoitGyj1orxBAFaxiM5ZroqoUIKdmuCdpjvPc2qBpeuEEsD
RXIeQULEyTpitb3g0oFdhJLceePh4pjaRGoYcnwFQ7rc/pohcA6bwQWqp4aRk56u
EDRUd1T7vetZcJXVMQsU5tIMlm6mLPVQ0vOOtuQmUQG232YWY5lzb0bDZ319au0W
8YOiJRxl2qiK5Xs/6vU3jSReOM8N3T+m5kmnhK98v0oJZxs03WjevHxSVca/+nF0
G6nyXaSLrzU570QkQ7h34kRE4yPQk5SBWXty2pfZr6uzmcE7DZmRQ3u4tbSuCUf0
xaMgiNNvP/02MvThJX+h37B6GZjRUxsRWRiAzTmJ5DMZlxcKfJQy+SObIVJk87fl
U2nHfPPK+8gDiHKGF6zr13WvFhVy3Kgaag08s6URXzkth50dUtw7yzOe7+PWWjHy
wJSVuAhZiDLYyOP1pS5XTVrS+ItAgyOxaU8dBF4EBA7sFl97cz+7RnrLIXG2IAXp
iRiJV62pxo75jpwcWe/Uc+axghnEYtYdHDaOFcXWxhKBx716AsnV/7EVo9X23Jcj
`protect END_PROTECTED
