`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V53RD7F8NdCrMjpjuo4dfTVuLmK77AHmjGrcGS0HXwOLlQ/psZWI/OeXboppwgLH
PotW6nZrT0l2vAZm8UYnwZmoSM0T1otoKVRQ/bc3WOXEFNUZGebm1uW4KNBb6HuV
SQReqDh81GiQDnQtLIPQk93lrHlAuu9E1gyIQsJf5YssUdPTH435SmMexpog76wK
SO2j65EyvmsF6XgroBqBlhlrcJGr952IeXdwq0lcq8ttVDEv3xQ7u77E9kEccoSi
a6flgE41a+uHbkDaLXguZkqxvskqamFcKyEY2c+b3lOE/yypjDK/RN2rlysu6Jfq
Z/dna6SS+FHywr7S/x1LY3WI0R2cQs+4s0/qmuXGZQhoEKDAvF+CkBee/FIdD21m
wBxh7tovkX++/Q7gy6kDOz6tQ5zMRjsX7VdpAF37gQvdvmstwq+BK7wpS7rvlckf
0+E5bwgiDb+NNgICfTa7yZHu4X70cBOjTZoUjEsAUm03zeG/guL7r/2NlfOlCrpr
cxPeYYFZ9Osk641G6nbJ2Brq5uM7sxa+/AfDZeH31L1y7u3SpctE42ZovF339CI5
9m3J/sbtjpNmcgLYZkd0kpy7w0RXAbEY2cVmJ6rYN+vVA9QenkmIk1u+QlanQATi
uU+QS/qY6I9v+DZaeImdmHghFrIV5jf3ukNw0cNlpQdqUrHQlKY3Gx3SFazV1hvY
teNWomfyq9wb4MXMZE4ovvelVDR1qqOKTI2N8PsD9ak=
`protect END_PROTECTED
