`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSvlhcaahROuQkMcNcTUrQH1V+2GRfiHKR+prX7A7hkw2A80/dMUnk8j2EbH04eH
TjnUPdGkWU1k7NLWmcjwjuixmnL+DBnT4ciDg0oSGGhgc7b3FL17pvMhdKsIbRhL
i/JUZ7sb6wdBj2783usHK/uAORvTgrlRra6Ki7iBQEN1XfTBb8avVze89G2zM5iP
uOkJ3n5mHgLyL+AMUZxoyiGZ/cP1ycFMWwk3Zkv01Pl+UASigXhWqOTkLDacVhLc
OYOarA+Z26gIeOa2QuAJ+XrVadTjhiRLfsDmtwUokbTqw9wO2CErIU7sa6VI25sx
wDjF2yG6MwHWkWtgntTpcijIfi31nAm7kHEurexPKLQrontMQwFcrhWv2quLxPPG
FG5a3OkPtl1rWZmk33MBMLQMZwzbKjRRzsQN4BS4Ge0nTGv3umXdAjQtPO9Jd3kV
AgTTjppe2K2guxhM9pI0Ebd76REEvtYkEyZHpbB2rffkWV9FIixDrC1Unbn4Hr6E
a9bXdDxGQvrVuT7FBtPshgRTXZsB8sCM5egX3LFUkXZHkU8il9WawqG4Lsk+gDpO
NHjLYud11eo9wnke9O/HJzs2N8j4462lsOLjcJV4v7B2OfJa6ju1KlD2tdgj560K
s0IVPyjFHTEpRrCTcz0hIO3ML/yTz0dEhrg6xZxfpLwAsaFDpdZ/aO6Gh5vD1g2i
xCIR6cUYZwhggiAzIaGrD7fuYY2a2cKaxaoznRjEjoVGToTk0Twp5qH/A7/HLHZy
yW8p7j9xfcp1OzuZ/0NgkrW8eikjlb1R4GABT0WLVdZvv6zddUfraotxDGe8lHoy
FO6dm9Og7rJVjON1OTL69vxMO+5av+S0PU+/ZhKUca50iQzbOytb32Dqf4dFuNYP
fmnff4iUYpYqdsgzwdQtRbZ48xfhldBm+jZOnJRMANzXbPcsVd9/2i+7Ulr6A7q5
zitc0sqckfhoVVJNQGnYG0uBIId6xGrgYc+jxzKd37zksAxPPAIAsxWN7eDSphT+
j2RnaFcPz0Or1qqLTFsTXkIhZviOOjXhzDcDZkmv0UpgQWPw8EbVfYNtk13yeabC
3bnzdbV3qNPzywjs7WJ9JHxSByIoCbOVURm9X0V62m1fg+7lTqFpUvjGiYug3uUY
iuXkUeAhct8vusbAtHaxXMc/N/alUhADzSsJ5BXfOx2Y/q5xOgh6sFP9xIYfJy7T
K8Q+Jwl+clz+53dioidIblqIPMfediGGJJdralJjQVV+pUaFf24XpHcuTsGPJAEV
hE6ANgUnEYzCoyn0N6XJiqr5wxE0rNifjSmdGXcEF+SEouc+mTvo+gWlQlJuuZ1L
6NTxl6ANLAzHGaZKFREqjZZAr9hRn33h0FJNq49H0uOVFpvrWJ/PQshPPoosWdix
JPwNtSnLAltTIjrcVL/pzEHlbt/UQYR6sqN76Z1KHBiDc1L0f796uLuDTgg2mKDH
m9ZM/9+45HD1qmKeKehwZjdPvvVt1W9AEAObZHdW5Tke3mvuwy4RDkryY2lsLplG
5zU3Ozzk8jBGSx+YAVUKI75pNkZSxSWKhCa/snuDvfI3QLLm9le1d4gptqNL0atO
m93NyFwAc/ztHqqgd+XC98x4W3PKLWDkPz9W3dyqRcE4S7Nh6q33Jq/pmjyuTx5y
TIvVTMudZAciuWiGnhFl1pPhOYzL/cBNIAe9psYTp0QDwXcngqfkM2mPISx26UFa
/eY7ZZHh7TapmVu1r81cEqI82Rkz1eU1lMWZs4v8NPdZhYG9Pur3sq61VKM2m+bx
DV7SDTLVid9ERzSB2t/IMttlpDTjY58niEqcpwyfkQsvkxURVs59FWE1yULHG4NN
h+koeeCR0Tl0z7nMzAB4GfYNTHeQYsYfCY+EFKwYqKNui14z3tLWTM8owyYS9X9o
BUxC793I4qHddGi3qf8xek3rG7+XOLVFSDKCxnRPNaQkIRxN3Fi6Js2bKgT+X+DU
5B+L3OXRJwuYKSir8Z2vojZV+js6HyCJD/DuAXanc7fML4xkqXoePVH+uKfmmXBV
18O+QSJbmya0rFzn2F+9HaAQaXStLcXkwe9xqGKwRSnFA4O+LomX1e80/AkldApM
t+BkEhtcLa2k9DYJKhg6HrEH+lJ6L3ds+3OXG2zzhA7lAvDHnq3c1bhJBehVlnnW
TzFfLKfZGbERzS3Ie8xd/kIamZ/dmcCI9SeBQGdv5VNNzE4hI5ZrqNurw0hyRow0
5TiPeaZi72r18/fYyXAzaZ7PsGLChxLauzs3YD6PFTS43RiMaDqjqpK4ZQv6lfxJ
hfOj2uwAMS6/ivM9zvWxh00kfsgd5CjZ+XBggDUJ2LAU5YTLky9oZqyQ5NFUuMz3
gkmPeV1ZBz+qOvYHjjX1et+M99JVBr6TD/bMsBNic4tx2ecBh6yaA7+erBB0wlO+
KXmHWlct4pCsSyO3DDM3sZl3nmvc/zk+GwJGxuxCvFTPwCXk0ns0vJ0VU10xb/zU
d2D0PkE1EL4/ZxPId7S13p7RlHw/0liBkehrbI1aHDTRc1FEG1+IiRuCZFmY71hC
hHOEIFnggvVOq0C53O9XQoYu7mZnbb245r69wPjz2d0D2JFMFxH/tFIb0UNzFbdK
fFhLS7qPARlRbzy0pSatsf9RGpoJjn5NjnMQp0GMByNuhEwVTsZP7A5Gb9XgGOpc
Wr7AOS+2FhDTR71JL4T8WhLxSKdhtjAGqa0ezckO4omOGdKmi2trC+t0JLavFNl+
lNDUUkppU2t2maHgTSvcWaY4vIujE7xTUoM0WVVql3/JCoUHWZntyC7IJh9eB7ak
naRU74Yo9LS4uAS0BikZgnzS2YdRTg2dcrLC8qtZaAJ4ep4QQnHFsl8Gf5rIfDXD
kg+E6phUTEP/uEBM7yhSmsxzWLJlXpDeBHNjtFTQ0btLwixJTvwIp7lU+U++z8mX
9B2xSJIF/goepV3ql7jwTVlzUI4SLjG7/xQOBRhkqOLVMqXnno3IRO+SOJq7n+qo
QUJmUhwVvVaKVF9tG981EFG4jX2FIFHrVMLxskdlsgYusnAlBOn6PfWQA02FSF4D
0DIClFNoXdzgTDy3Db7KPdfAJBA6hdq14ytTE17x04AQaskme38UWC/SIDDs4Eoc
8FVLbfVlwA1Yi4OfvbQFWu0COqkKwOxxid8FlPYmOAowQ0buawr2b2jr0Vi5zoi+
UMcxo6HU38mnKw6RH/Zoq7bvCsooE4HrIPixqCwAawZniDkdtEUPgs/5vsEZFnkd
wI+J05S+1vmEFM4YvFtFFx75J0QA3GjyK2TRPX9EjUG4OqXM0sRuJ9JDjmzrfBel
m1s0PvfWWoUqx4mQGhBJlvQhmdE8qFZpz4k+V2lAgAezws8waxJlB6of/AeFFzfu
oa9hHKds70c/q5DZxb0SToOfmXMJzGKRVltdgLzoVzh71E5JseS5n5z4BpDkPqOq
1xARXVjPQY+sCR22hwuIl+IFV0CiupVPoeFdJovcGDQC3GlAlJZazPZ+LwJST9uJ
HpNdiZi2ekYYhsPmkpW1j6InIeg29xg1PfrZg8o5J9F5UDM9j0/94v08RGrf+4Q0
Y5OT/nHcSca1DHBKPgr6kqlu5gEQq+Zgsi4tPnE0AntiHTyWv/aFJx3CrjTJu+YI
EE7GI40kAZaxPg8R2VTRrtAn0oN+Ksl+faBpXTiZlR8aLdQZSmJHLBBxQRywJVVc
1In2+K4R0RrMDngSLkC6DcChUooUsNmg99JvyA3yoCQkXvhjpSNo+uH3kN6hyHlN
b23a9Znydwb7UGY4AtrPR3dq+pJwpx5JnAp5XJApgBgvWekC2bzdjnkLK1rzVzNa
bd1S4aZHnCAsy8y3TW387bbwUJxiqqaMr/Ur3X6oiCLe1WA6RU/7zs1gjRah0IkX
QfQQQfrX94y/4OQQTgNVHFXqkY8TLfLmOf/v2Hg2YWCEej4C/eY8XC7sI6xiuYgK
M8wp0Xm86dUivyccbm9E0mwZL0umR82Keikaww3ZgzqllxoXkmEWFlx6KS7vE0Pu
GcnOmTNiH8qrROGaQyRkBehQhvsyoeoL6tPsgdMTKogPX5TvDhrMylLWjFeM//NY
/GWLZSxNvDJR1uus40rQ+0qR+3ZGJ9FwoH8DRgyX0VmTYt+Gnp2W27b4eAicAozZ
eXTXSSAiu0K+VSMTxlPCNtr54U756Zp2yB/T74mDYP4iI0qzS/BxpWBXsu14o+7X
vhXBKfKSoJ+J1C8KIHP8UMm474+kMX19qvOy8ra1WEAR9XYPE/3uuBnxip/ucLPs
hg/kyXk+yCm7cGloaefoFKJRM+WR09iOMS04ZrKy15w9thEZnBsc2ol2EL/n6pmw
x0lnalTth55EfsQK/160oq/5Qhm5NoNdAlnxoLqu4LJFCQ/Qh9bjd8sJ1ZmFZfOP
jk2S4p0Tk6w21IXoxmfb5GLo+1XfLgZ38FjQgdf2y1/F86AWQAagssXYkUmAu2fy
/WtRfvYw+ZURUdA0CmNRpzzmjbNqtJAEE+aYdCapyleiqugKiq+5TIJH3vk7guhK
AyELsgCv2uK6h+hkztZI4VbhC8g0g94RwUdWDYjil1krVyYeSKDcKkK4w+q3zpSJ
/aQq/MgFkTeMNebXCJdInqNQh4oGC8Up6lspKU72T5bNFlaFDTGRJVylPYejYbLR
VqY5pZjn12cdGvQeHC2RmwyHWbB3tnaVI526sb4P/+08OHATzI1+MHGoIsDfzWa9
I/Q/Ut5X87AOeylqIFHceLJQ/AQMKvrmuOnW6qdDttjlRA7MTdsiTALxWvDjBh8T
WvZDxt6eTZ9PLkG1wSwKiT3DYThwnmtF7zny0v00MgdJr8WQfCNT0eB9XnOIT0dN
DPr7ARxA7hcTW6KqjNsxZQgWicsoCTGH4qIHDCKygO8terE7i5JPhpf1D+UFD4oH
mxun5qzlv+boBQjvyYgjqjizJbBii7WDJlSf6OEGVd25wUlUILU7cJa4mETKSHbC
+lsOE8lNG1b5/APIFG3tRlcVG1Hbtyq5RNuUR9JpN9V/GVeV7yDAsHQCEbE3qBNl
YOXqQK1RXYW6uyzEPMnDcaVKzExcEQYD7ZmiRcNLW713UK9IQ48muWbBCncQojOb
b/1m6WmhPJbqSMRtb8xqeCJfY7E7cUdQKk3NJ6HL9Wyw9y5NocN3lXQtYul5rc2g
bipk9MoMwAVBXxOkDbqsZojOVbBGHmRWARedq+jISw31fNtUZAxK6Bvba+hj0kig
FVmJStn1hOaDY0mzlCuRC8DJuBbHwHtc8HeHmSV+3rOaP0NaW/JVpmvATT8sMSVW
CwUld/6ophOEbNnQzLuCUfYhSogm9Jjqr/KMk7sNNyI4GkYxRS0iq+eHp5D/5pmJ
96Mh1HRDKezpTeRGMqtiRvH1lqGxlujSGTwn16wkghudB7RQNzL3bMhR/soq8ttC
4blo4sW0LydtrfU6iUwWdP3yl2pbj8xu8sfbPEgWnwIZvcw7Y6iwNzeiJ6ecJcQp
v/O40v1XDU+B8Wq4JyM63aV1myl8YeMZJs2i+YQgZ/88DMJ45uhX3lSlSIIKgF95
Mj/2qJZFmMkf910P+XO6PrnSPapRUDdZMsCf1UIOILJG4n/wqsVqvfYcVsLzNByn
v7/xwpydrmNNxpt9gdm9FTJmucfEUMc665OXhQB+49u9fXNkYuzRbOyX5KjKFWDw
oRdqvK9svoJxEm2WZLQ6HwlIIzWkajhL9Mx13FHkoEONet3bwqELo49SWevUhQEU
pWS5KpfARITIVmFR6JxJl+VoT0QylulaaeQyNmRGzoZecHj49+SR+uvr0yIKdiwy
tTJfmEfJVNfOARb4+Rjs7YUiD/RB7p0A3Y/WscQm14NIP8hQoTQLy1TpkKSFuULQ
Ez30FOdvkKHY9jeHadEVTmhds5I49ePEwJerVRZ/ywSnz8R7MGuv5fbhehm1D/Mh
zQ0mym65K2LP8ZfsucOA/YpIhorjT8TO+KyjfdrrTU+NUCt3oYVomhSIRHbKByWQ
hph9JYEh2Sysc2FG9d5xjd+iVx5TEfq1UQmIV3yskbBxfceTUoZ8L2QcJgM2hX7E
272iNN4mmNFkGbatYPJN2AUv0kzlFi29RdUKhEG7gf/i+vw8p1nx15mYidy+Zkvz
VKaPIqaN9RnT1ldbWG23FUQQgjH5B2lwHvkVDpnv8+s8zJuQLyL3p4XrTKiXC44n
p3HOiSTg7d4UuHrAiDfus54S1Os1h+fZprezVSCyuaex436fHPvqGJ2OczQhM2Dy
seSDFAAspRgzOgspIhi/8UwIAQfrdhdaFNib5bGTvtWNWfdMQUEwHOu5faiRAa49
3o1xw7iwYixunRQ5rfk3zQ/FZgfkL3gInBfuT1ynNVPQBygRTc4faFHUA5/EZw+L
G1wTufFnnCP97/OfSx1a/5yNCSULGLUKY0hec+cTLkInW+f1JnQUNQiUPfTWhO7U
CscahjqOQ9rXJd3x/vf3dR68PQNJQK7lYQWMjvnSNDyiklfVKfTZ0CPL8vjiiL2H
2Kvg4ZNRw/xNRrKz4/XJThkwzjEw97lJz3wFTR/IPU/13zDpCRDXe1EjuE7ZRkc4
jIKScQz4GSg9qiESoeje7Xa5mnsJLVM42SXm17iBr4sF0HB/inSVM+OsKH6MfQ77
l1T8KD6lw2LOoOjSGwFKbwB675UQiestjkB0YybWA1FRQfmiKewax5cUKh3nmFhH
F78r6H4/KtmHDayoAUj941G5T9FD+EyrZmwDPHf4m+jfNmQjSqbY9GPD2rXZMYkZ
JyuvntbUndpWzro6E7GdLcwgjqT/ultacNQCCjGXgg504tt4rtBMWDdrJbGUqno4
421IJPoD3itmLU6D/w8hiRvYd1pmQA32LSa7Wh1wk9fNSwA1vDOjzD443NXDINMx
8A0uFsS2GHI/TRP1/V7cneWwOeHb4NpsmtcVJsUhNNX/ZVa2wHOv7CLXxr7vc+uU
YhsWqQUNy2Jv0lfralBGNbu7tNfNpVhTbtvc2fuB/qZa/dh4yPLorUSOUCPtC/dl
V8YEn6WkrIcn4PmjbdE8KRA7++aFYkbXtM1o8j55YRV6WsV7/SFUCO6NH04WR1hn
MC5nUCyuaK9/nKGMKug+IcpoNWJNuA3T4shO52EjpPKwRBkK6C58jrdWEz/0A4a7
03Y4DxnRdic61r8DhvU3IatS1YD8E062qN8qcV1QbPXArofvtO41Nshrp69kDmiZ
D774p5QkAWcqaZuRwyfNlndQCMU2bDFMSwhFHmmWGI4ZFL1wSnnk8tzoctotCIN6
xAcfX9MEZEXcosJVYZschY2t66mRCYhRAApCdAe7SsD3RRUlz7cfKeYd6trOr01u
rVvXjirylXZ0e3AO0qeSumq1jm/LQwx+yQ7m3reVuD/IBSDLccOJf7aGk/UiU9nh
nkB0Nng7Ym/yQgNJethAl8OK8gSCB64kTfQgG7ThteFl4IP3X6vd67iBp3aQVHy0
7m5cRIN4XGsj4KIEu3VNQgr+9sBlmrwg5wLFv1vPdruEp6IjyUai9DXX1g2K3wKR
s2Lwzs7B1oLiqCvASMV/e2gJZVlvZF8adDF42aIx1qABnDnbUmwQ4uQ8ktOuz/Ar
HiNL8q09DJm/xhEVercrDzupHrUXs8Fz2l+eJfpLR5M1aeH6AjkCCiOWwnfZIet1
5bsX2/Jap3OkEYkaW3Hqhc5YqPmegLKBkTT19mALTb+BkY9JFw5UUVThRjL6q2YV
y8zErCzDNhIyz6CxWmlCKQOHoXa6ErqIL292tcSAghmb+wd2uvPJ3P7kIA483UDx
GtT8i+zecBnmAX+GexSBqu5dOsGZhuXsIYacJxpzr83eOLgoiODabwKA5hrSyw7w
KpF4mYgzXOkdWqeK7N9VyuBfqgjmhFAoBcQtSU4KshgMtbw/eDYgHLsbdUSiUC5h
rCLos04aF9kvzvcwrmpUxY1fSSbXRhyZg9+owcfqwV11n+adsV9P+XEXrTOHCXZV
nW10eG/N7WucFIeiKpWvTSML8gugvM1mUmgypzWNydxj68QkPHQDySDls68kWVgU
Lequm2BB4OTCWv+6lRW3mju8fQ/UHyDSD/7yuYXmqRDWoyF0hlsOSPN1+UkNng0s
Zj7wxSznln50MSDjWPesYOnhcFolhzDDNMEdYWfU+8lHeJuPTZ73YiXRNuOdS3lm
L/I39j8tYDCpcRmRW2UDUkrBg/uHLtGboMVeIwc0ZNKnv0TPDYGM2hYG4nCBFY3P
anYvRI7DPc4JK6R9LHS+oDJaei0icH/dD1jaeS2zBHgqXiT9ymJxXSIemGEuQbw/
VVyg5inmDhSISeVaC04IqPvhGDWx0v7Rzvh7/ZGNqQFfa8KTK2lYMHQQ6UdaVHF2
T2t9ZjM+8aBKlmWM9vFfQ1v3grPizo4eyg1Q/wRwPORXe7nMRF9e3/o7x/Qv6jl/
S9QfwbgOdJZ1LGMghUAvBOwXcuq0C6Tctogpv0GLjYlq6xt9SlI1DhUXNfrxoRHn
gMRaQ1+vzBRJWnZC4fJ/dUTZnELHDv5zkjy6ZxtbaZvy69bRh5xoppUShcSYeuYJ
Sd4V3hGXLrJxhN02XjVQ4s/NrLLuWFUihkTbW0yDFaCv6dNl2/VREz8s4eRWQgqw
cFxQcC9bt/0PpraOc/sZl0oOlIAcmtDVWnClfwgPlCpxAgzG6MiG6T+Pb5hUGyO+
9bfFWeuThXXHSMhuyEpsJuF6n8DNyjfYmUMwNkxaPX9e6QHj8vgwnHLuyA5sznHb
WxIGhJT2XXyTNIPYavaxmw/18940yVCY83z8ITKXvVA1noH8au6WxomRPLRh3QMH
E2wjPlxM12f6hIXN9/mxXO2hDEqiN+YiNvnsHW5Ef9i6g+/XZuVCsMIdG/flFbaQ
yZ21O/ZI96Ey1qi0XtsxfKHBbiFpolVsKE7XCHsL7ODqCDz4QbqRcexKwwRV+DO6
y4LTBBjMj5WxtxgKUxiST5rxMHm6YhV145MohXYInMN4EO14XjRmjHM5sKkeveRR
N5D/RMoaPXNfKLgJ4/ezFWY1/KKo2wz3Cdo0xJM7Fqav8JkjfpIqa++40fVBKBrf
wGzB+H8//4/CLkQcyS+qrC+vn9onk5HoKBnEkzhu4z+vTU2Hj9HprhA+MXxm5nKH
D7k0+O43dlm19oXE5hK+XT4iMv2gCeknYXxLdGf6587SZYpPSXXkNvq/YMYHpTgG
HOlOmwYiS1jgU2G5D6cSyGfeIpRs1R1YxoRCcm6NYbXsVQyc1jxezaIqaWOt7Zln
oh1gEKMl0JjqMRsKKcym58KfT2IfBNmg1u+LtF1cDo/tFKrf/iu8KcDHd9nfE4Jh
JKSMREPBTzYKRtwqEhB11poDnzpvTKF4rDM9UF5gGIT6yJW7NGqT3mYOpC5oFGAc
RZaMu2I4VLW/UZjcTwGXEQZHG9RXBjaaF45SdTUmrV9tOyCcYmsfiJtwMTnXHMn1
wnxk3YMu7SrrqMP6Qs/4DjhOANWL5/Cj9OnGdSOou/wuJKEmsF6vfkN1DAesHQbK
88OQViZTB/tEfeORkRwUUPXJDyfJ0VRMZUGdsCcnP2zrUjHRY1NSvXDtEyTzFxRo
eNyLtO0P3bA1pMsoADeElzoYJaLwzmecby8dPaut5Gv2OsKYFDo2Lxl4CPkGxcxM
pGI6RufhL3DNeJYEk4NS6DOnSgHwu6dtBMeT8cEainEzsl/a998S8oKkWGFOQORH
r7jXLLjNGOHRCv/AXosk4J27c7xBwMI3Js+xGMnu22ELcFnx1ZaEqlg5HKHxOsiv
1kwOulvqeoOP7tfQ5koXi5l8L4WtuyBS8YvBOeNHqKHYdUk1Zf87HtA2nfDhL8VV
/No6tQu8jrIvXChE6vLI1c4CZzpX8b9CIXL/cgUgRKedkcM0OOKwaNhb6OZINWrT
2T2oEIw51utu1DwcaF0uz+sIIQKh+P7LpOWfoAzTnZrZ7oLcSIir0EoD/b7UrG74
I5RmHFP1keOiUxJ46+BvaBHyW5QHGktqoP4uDmG2vuvk4QHDewRdQkfBBCkZGBpS
KOnluF4HrhICgbDFMODG2ZQKH/daTzMN7nq4UZY+jyIMRNot95B98QKSZdoMyiMg
QHdU324RsjH1kX6q6E3EvJPics1uEpghSmxhDw9raz+1FlYg0bivnFRJYsndX1Vd
fy5lNrTiL0bdo2GSMZWjU6OKkMX2vIKkm3vusLvHN1yf9miVIq90BdlqCdcqeWg7
DqDEYAadYejU4zpo3GRXMwNEv2i8lIv3FAoG2RD50JyYYLmWOWIv9WALOf/m+o5h
UZEPvWrarDWgdmoXaEEg8OVPquFQv+VYJHI061Stv+wmI7EghR3jKOZDKJnI3kYc
retb4srHvhT9zUS0Nm8viLV4nZlnlMjofnRLkmmGQ8/Q21hvZ91z+ynPlIHNO4jA
ChapOQdZ313jsBRhjjvk/2DvrHPlx/aexxSGVd8mhICzReyBrLwSpGMmMkJLxXPi
XEOJcPD6aoImFCzLPfkzsYmab57s+t/qNmsoFBodbG0gvdGa/E3WDqvMme4QoNru
74vcwXAhSw9QC1L4DoObP84wo+Ae3U7uQnhFJfgpzQAE8XWT0woFodlVFswnc3MQ
k4F0c8SVY0SuXHc1/ORWR66zy0iG5meEJxWyw468xrgsBW8Wa+2BRMk8gLU2oWtv
EUx2gXK4vk7O48Uh7DnyaSi+3EsB+wvHiw1bAdLAo4qC2QML4lfSfYtkm9ejFraF
JZMACkab9YInrpiFnRfzuLiUh85BTouM9Yurg5WWvL5JPmMfthpKRHsm9Ef6ELsu
a6ioS4VM2i8c8TOnYkP4X4D7UPkZ1UGq/OKss2bT6PrEW4006tpcgA5a8cX9OCr1
Px8zs+nSVck2zNd71M6R9kSWjqsnHpp4Oz8zsNsHnLlOEk7ARXtu7LGcBUaCaZ1F
jFuVOjR8skbSFTsfs3X0DYsuz/pAaLLeNTsAoKqkIsraIA8HQAhV6X3ODMD41vl5
ZX8qBjK7y1Cu8A3YyaSHq9wyYtQpCy3LND1xUFrjb3LRVDxiJ+PrBxgkjdYfvAPy
2NnTeAbjsdgRyHCmVJiHlugKcHoimtpgGnO1SE4q1rVjet4u/rE2PnmJ/3Dq310a
ZgCjVF4ratgJMA7zVsD7cp/y7RMlEgn9y6cKj/nlP/tKzolwqOzZqx+KMGuD8B1z
pMNJGHtSqyJJnJU5fiyTRC55jP7HLxmwinam9wyZpehXX0i2ihjSbdCfBKRHfjE5
T8sAXcqwSvr9Bp6QyurBkPyd9xrTKmCEUTh2GZ7lAPhEIFly51cI2R43Ao44Expy
bftpb1nXhNCUyH4DauEV9ykAxwXouBf2C5V5BhX4COo/pzqHjikOmW40ARa5aks4
1ExSWQMuXh/iyeAwXA4hx0cYXJqM1S1SWN2lwT9BL1TEGQJgl+VkTuoisxWNEBv8
vOYiO9vQpTl57V18yokSPk98ZyItZ5AAqSK7iEYTg9vZWcHhmCjrNbb/hNmAOggi
K2+gVwTGWxrXoZMVcdDqpS3gOyzB2kderai1wVb2UJg11vdsKTMVUI1NqbbNOmF9
HctsffCPvuo9gulFFRWcowUDuhwAlR+hq8E6BP01LxgGC7IJBhuWY+GxX7GOEEpW
+wqinVhpvwvDlSJBrPdmupw9gny9YOWO4jko8/kfWe4dm1AZQMeGMWo0YBO4Clqr
L2ARxUh+a0LLxNiIE61p5zLxEKkJbbMynoUCAEpvOvvEHvnIiFzOmvPqset3Ylws
Bg10IX9dluPvnSreThdURbkWnasXrjROsJBhCf9o9wMgUOkSrIXmbV1QdAW9minr
R8iq4n9bp10IdKiYxfcGcFP5TV4WPldQroO3sDCM0EMzG3wnBAdZqlrFVwQW/Udi
kF5WkEG+w/G6z00cv7glFT12/adihxMMMbz4hGe7z2lLPZmk0tMKq+CFWUK1QPY/
uNUaQeBCWb790RxVoh8tYMm+gJhsyhQi+1seMilkmprTeUKuFC0UxGcWSyWVudld
tjWd3WEKqjhWT4P8uzftWdt4ChydY0RNPHrs5BvaOv68c3MIKD9m6kwIw6JPj9B0
S8YVFdu3VyAJ8JdHsdxMPHpUHhuXKiu4fxcHcwHy6lKFF9hN4tD3BLOT3KdUC4/u
37EYfuPWc3pvByu7SRVMJPfeM5KHylFin5oPXHtyX5jlryQ29alHXgRhc8dYXAew
NuEOcLDB3enYCLnrJ7A3Oz/ED7RMLDBNR4V+MRFJBj1lydAFJ6mYpz0R2XiZWF7X
kud+U981GIxQf8S3Q/AsXPKeTTHyqogyvuyCNbnYgICGJ9kHHHgPv37BGL+Yu1+b
IfvAgkihgUKfhwn4nmUKD3t9OcVkghVZvP2GIiK240Z5calsda3Yv0LIkwEyC8+b
ButSfXQYr+aH5wplrLOpoIg3a4+6bT3NrIuhHB3VmufqJrDp7an9p1vuH7bSgGTL
Pbv6qXvbUIx8P8ThjoyNhawMxroH6NawMof5zUyxndFkV1W5oGTZH+PU1q0zgyme
nMPWz7I/XGwQRN8RFr0w3xqVnP1uqYuMrYspNlf9M1wjI+VAxj6o0/LxnH2TTR53
hheAS9hDZoj4al/EUNWzW3AmO/vNCIiSC8gq61lyS3Qp7ONkKkzYoetsYf3PB7wh
0pm1+fRAOSfiqBEmOdkL7GKkhCY190GBMcOkU4fgLRRrUhVwkPLMcBuh2y0RtNpi
iYPe5ydEDc7mMpWi1D05TbYaWq3JTjze07uYvRnqM9SBRtLAb03bLl2f8XjDZTDT
iIuDnI1nZa6gadtP8lReq082iB+/j2tbangHet/c2HWXHIdznZVymutuFxUgJou7
iUbkb/KrEAmAZssyZwuGHBckUpxTvR5yE+HQ9Fg9JlV7wevlN7F/mTAE/0/IQM1P
sw6w3Fjk5FcLPfbBR6OovtFA3x4Y3ee2wdMWhbPVzJg2XYJg6YtShuNP4URnUAbv
In/XBy1jLz9MixWqHZyYxDSiQa31ohcYZBPCGMwtAzol5nHoMX7nzjCrucYzUK5P
tUWpmXt+pgEC4q7OMybbTBz30FIcOHqqeRGnLJt4jfeM5SWzjbRJLoF8Zb0ufSbL
8I648YauJIYQkH2kYxy8WZF6AVQ+yktyhe+CHsJvKiAygVzmm+fKbNESbJMXrKA/
Ibd3z3bSVM4Oim66hVS7ravUzGSApjgxoSGKt07sBjf4zXMR51isIwQrpTmuxjhI
p20OdL1thPb4JTUkLQZN732WJ5o9ajhzOPk846tq4S5ZyacsRscY3DUTYK3GIgBR
GSSrNX+Fa0SpMlHqO8eJ9mhRdtcOcCa5oi7NdbxFLVr8QqKJ50lu6PZDTVyONqTP
Z6lQ0ViyZuyZXRnSLz8XVQHvzFvQuhqvgGhzkYrQ2OfLsCPF8QGp7sVBOXNHlZLs
vvjXxhRaU83w+MCc98Mwx9z8VsjmoZ/wT0fNVccw1f+tmfhae0J1vzZ0UOzZom7j
D6uVg78ggISSJG5pGS/V1eIWHOv2jYS5cgVNfucAuDR1iqB2f7D+zIzhsUrh+HbZ
f054o95p5+z+CqdfebvBTaCMP+aIKGWjVyubEQhtJVFBlql1jJAX4gOqnXgXz8yq
wXBj1Jf2M5yDvao2IRkIkoVvecGX0rWuUHFqz+1vxh7rxxIjsmE6UU/L0rIeaYEb
BomAsQuRpg3XnVpXOhn71cS7BUoFabLJXYXzjNbCjpPPUaqJvHm+j6x1Dp8xXP6V
rn/Pp4VqU2x/kJdx36TWFRKjSz77ouFr4bZIzu6JYs0+ims6S5GU/C+GlzyZLqFw
ZAKK8dw1EMd54kgfu3cw3ucM34XQXLPmbIAySCPlhjRF+eo888XK7govrAJidgsy
RE+iDBX50Ei9bi//2llMtsrEYmj9hMGg9Odf/m7ftZG3EVEib8rxvfu9CwHXNN8o
fDw3ug24XJUB0lDGHPnsAKqE7x+Z0FkxFrMDsO2LwKXtn5kyLaKRDtq+Ppie4eVC
t2fuTBqC7v64/rcpaANG6fuWZO4rcTrliiuD8E9HziYvNdcnP2z1MekRuW9khZ/O
Ks0EOm3rqjHyZY6AeADH/6nM/tXCU4ij5pjSdr9kIz6SaSEfKbMyZGxfH3Xjfqbn
6aBJ/SprC+nSJqMiZSPY/Va7ehi3O7oIR2HZ03fcNNiYT3fgPUqhK6drQEf97+9c
1WxYIDu1zM+5ezaBSUXluwEVJKu/HrGZ20ksCy6FRc7nfpTaLlsUTV7GlVDhMdpF
9VZJ3eD37LA/rTJj9WH00vHvENj4HDPlu3ckwcYrUn+1HQ+XfYJP0uAthpaBRFkn
oEXX9PsLyOqufPwdy1/wbZkl6amTgmyUT6OlWh3oOh5FoFU8i77iy1ugN3XNypUb
P7GYaAIUtwgoskhNjxPzBFuTeqFKAHwZ06VYudiAOTwJgUd7tSTOkILnaMfGLjUA
H48i+gM7VcIq+qkKvCThC4JsBbAOfy+q+c0C5VwMrECZNzLnMoOovl9BNGnh5kle
z4Wzqrwe92r8vwKjdR3aPRiogPbL0E4G6qE4b8Si3zC8miSQAiVtJUSTb5iIxi5R
mEqHBjaVfA8sJq/lKpbamVg7u4syoaRW1F8P1Y4UK2Gpx75R6V3IJdG0jxSJsuN+
Lbxs19DoAMizE5m0NJd371QhJY8cMJ2u2ujG5in8ubcFX6lWhL/7bQ0qFsLmOUFI
k+K1OJbOulN7eJFCovKDLOwNwPa3HogE9CIpJT1sEPhXkItTzpi2krGcQKOhCLhA
121lzrmCk1mvHtSUK7oJgOaAWAfVw83adsDG1y7mMFQ9pvFMClAkKHKhqFZcrCts
0PHz41WdPjZ0BuEtDvoqRBQFZAHYLk1eL/ySyJP6fA/ritFMu0PYMAQQVmS2RF2k
CI5xwzHhb6RcNK5DIdeLX4Rm4m9dziaH1M6u8rZ9lYdQBT/jOneSTw1IkHLYxnoY
PQWz6tL56VyLq6QPBeNjRcteI1VOOI9nMUQt83Uf8lQpE3AsdBZvSCQzK4P00vDv
9D+3L6vnekRty9wwGgxJBqj+2qUI9DX8NDGDGskYtgd9xoDXixwL3CLRvKCnHZwa
e50DBuXsXRV9v8ybY+NAZFzRrI6HWrOrG0lKQo1UWU/NmeiWC1gl0iNYlDIfJvRv
Gqcpvo7VD22VtpLRkRYZyO9BameUA3sx4LAjky970oT+IEE9EC6A0xGnuFEq6ZVw
cYo5gts5dZ7j0Ri1ktaIK7HXlr0OUgbpdAZUDspl845QDb5Vi4zh09voPm1C3oBf
qJVJ7PZ//28rSnbWKJn/qip6BrjxCPaToSVvmSq1tw/bGHcLexRP3IWFirAE6Mk4
ePexTNrxmbR36mR456F3HvQadwsBC3dwFb4Knv+G+TLebs+yamDbYlXkiJDRFejq
4y7h0+oqaWDBeUXuCcwOQgkCIETgcNtmd8MBaoEFj98nGMQ8sE79Lde4bfmHSVmK
9yX9EarftMf5lomc4HTH9Esa28JyYfHntgt33cI0jzBG5rsh2lL3G8aTsemrxLoH
RI9AUHOZrWesrDh5X6Mmu2CNM5vV3D7bTniSNW+rYD5lRFneQYkyhseEoi+SBvDS
jwaOSN8JGtSZvlHyKInN86SqXEMPVWOkz3OKafQJ8aJxwGSxjH4M1utywCsp+NVB
olZBt7XOCWAcjYQBncsFN5paRmVPNYJ8RDzxi9XE5DfgNPLCOEIqeHmDbrNP2qVs
Kb+UDewIBb4EmWuGBOk5BxcFNZbGS+56LL/7g3peaO9IvSyn3CsfxiZW81De8EEu
xMXOM6W34X2FaZWK0rwEvx8ZprJFmYHEWN6bFwJj/HxlXH8JyIYdM4/naPhm9gyK
eZYT8Ek4LT3RtIMMmMALMXEOoSX7CyYjrXUOZGRpsusvlh4H1NcfEnAkjZMiweOi
T0VMbe2pESlOXC7UjeeYT8ot8pu1oUk+Z4xM4I2PbV6gn8dchY+o59BG0O0wD+C8
HD+gv6IXw367uWhPC1QDZRh0JNKflTojNEUBOcWSHP+DIzU+1197ItlvOFfTBSdk
6+F6tfpS+9Nqxo3teSCyy/auevYLRWhh9pMS9vLxogmvvLSs9nKjH47rgaMNrZXE
yT4B/JZQAsLdBOorwSPDl5+1J+UGH9mn5g4GJp11KkLxyl2MKQ7xM2pYyG069aYy
qb5RCe/77nFSFFU62ka7OAiKAQacSJeM064VIFprJxRIqEbuukCKzdAiNAFIXJGV
rDfJKO/F64xLo6/4KOjoWSglnDD3rkPdugZ+R8HaxFzXeFRWw3pu9eJ8CAoPZnsK
tlymif2d5ZOgHEpS1aUjuQ0GPh4J7YW6uYGaXCPJ2brdX9XJkU52/DdtqYX8NZi3
b9frWuwHR0jBfKLoj2XQjLpx3hSRGnRgaUZUnfjSWG+nrErGkEbfSlsB1CuudLeg
bpomwj+iYxz3mK2SzgC5srVCxxRGoID2pRG9dgdx8mwcCqCEnmC9EKUta6xmVmaV
H3xQgdiUAn2gqW0llwxwztjRtypWGC71p57kxCPYvWQrJqpuhYzjHb8EXXGwtl+2
LtYMofW40ZLtKYO8SvhTfkckz0kRh/lreJneWvHtwQNN8BRZYIoDet8M61Wv6B/a
OamK+5rVoPKFCbaWoq8r9I3I7k+e4pEjoXqdVMmdK27v4UbWbUVm+st1xE1xOroV
u5EIown2wWDhmXlRQLC01fUBDGwlw+0ut8C7oBY+DQwTqFaliqbMUu+RUGqt34Zp
bukjHxFlpzTCa/yWLiqaBFieXmYSO9VhOTIdrb8YvQFAyG73/Xjz2xNt5ps8rM2b
QE9t8Vgx90KHibm/rbVLYZun1eXPTtux0n9W5Yql9YQHajJHBlfS//9JedVsXKk9
ADlT2s9qqT0ZeeA8QqLlB6/9qwnBZuJMVt9wtQDPkicu9StkChbtfPRmbqzExEe3
yc5atxAfwAXC2UsBC1deVakEMAe31enfjFX2S6YD66HNaj5uFvWmxLInp2KEsL3s
B0h2dlbK7svz9TkNv574IMdQQ6WB8twnaVn1zCAh2u0m/m1mDEaVFYEWBKj7hdoz
KbxJv9fF+V+5zwOAdWKdwyZ02iazD06SYlXW2EbcNd85TzHPeEf56Z3iTSOc7Scf
Ybcki0WkF9Tle991JVsXnCzU82oXcEWhMbuuv0i5rUDFffpwl0x3jZLX3Pikrbul
Tkr1nqkSMzWNzFzA7JtEyl5znGhUlRWsMwVp85szuQbSMCCtKWRt1LZfnbXWK8bQ
NBQ3Zy7nRtKRSU7qd0ag8Ar+gytahEobxwWiJoXdHkoL00gRot22rCYqxWiLoT5o
jiI8tr4c3fxDVj4MPNMlhCkzLKCdabetppemjaEiB9MqXKheka+iWFQuUEJgYnQe
PsUUp91Ild2JLn+raJ5QSA1VU3DnBwdLVIprlWcWcByeXSZtO688naR+MQkw+VQW
UJHvvTxsf4PedKjqt2GFk9rxPwR9l0ik8JMt91bjVEFqxbhkhveEyvK+TfSP3cvI
G8oLfxzpEb63fMGYswk21g1A8pswN/cVvyyzEpkb8W6TPZeErymz8BrmRMIsIK8+
obwYxyl4F/xvWR0jzl5u2QuDHfjermtO/ROkZG9GR4ZrEd3cx087DwrUQFQmSZjn
9Io6GI7wMiezSUsuDGFuFh6e+JOVaOw4z+1jCOtf+2aeIYtgRaBZ3OYOVdxTFP96
qkozmlolTzKyk+t3sVGGD1c58/M6mFW61O9agGjPFsO0HAdcVtrVUZT8jK79NeTG
IC3vciBjIxEO4iqYaS62WcyuHvusnnvk3IQQ9kPYzqmCl/rfjkHX2D10B+VeUA8c
mQ+lK6zBo+udCAhazGDFvIL5pHA/3noQc1iYjxp4N7nnVrRIRc82GfgQ6Omosg39
yj4kPskyuKZ9GAB9XNMQ/Vc0J/nV/nclqryeaggZJeDo7DQdDFW+RKD7FxmCYd26
lrZumZTIIZN+FZB8oVvVssih3f/7k2wQi+nWLBPfydgStwJlszCbEv3Ef4/NzVtQ
EVt57UnyYd8o0uVyjHIIaFEBZuSuWNx7ZkgV7yG0vTzr/awq/b5vWsE7WJ05QhI9
3DDtwq/BUoBvPenzVLS9BgPLoLJYMxkvBHe5dM6Mdh3hYJcW9RZcrRirwK/UrUjd
zI7C2ODqL/5UCToPLbldI6bgLedsBn4sQS6i0DImNjY4IXGb4aGs4q6SMexPk/ks
m9hGw8lSJjlTcJDQhLs4d1lDcQgLeP2d7IubVat7ufMGoEk0S3oU/GHb0b4eJNrq
0YTpIUahYQDKxae8/UxImd3cuEml9N6PjRoh48rY8Q0K+OwnA+RRY4OrRpJUs64H
nvjIEO5ChNcz6AgUFjl1fm2uzUVA0vR/I4EkRx+ICmtuA5y2L+/6Xa+A79LDHXjB
FlxP7Yxr2y0FZAIYpRqOiHJUtR4+nT6AQIRrykN0STw0ZO42bwhUJLy0mPySJ/X7
E9NkQKI/tdnbJ+8A2BDodDN1+Thc8KJqu+0bysOwVneLnKNJLJa6W9EMF+ikw9qI
USx9o4sujTRmN5hqJCMUrWE5+oEBRZCmT9W/FyZnDV3XxZ6YiwBcB4t5ko7Op/R2
YBnO2QvPONZ5uQ9PadBsbYg06y1sRt1HsN7LvfMQUF7plIdkFO42wKwM4Dlw5K1d
Kly3Jv0/XAtn4tTqzsL8LQ0udhAJRfnUAglcMOHHXY0qZ3jTVR7NTP3WCJqxvSIF
QYf/0k5SYy9t3krM+1X9SmQJsJwfCiKVleSPWAVLides5YQvv8lyuzypftS2R6zS
YCqeaGkXMa/6UdwhH+ox7+1ih8NGpS9QbPwR1WR1VwwQYKfR0YwuadquQY7ZIs1J
kI3rY0+5Bpb5HGEP9iXyeQyxaHmUmjFhPiyeI8a+fxEzPJI/QlqG4GYz32uUKgRj
hLH/BZpY05iyKzwIjCeSZ9qvkeLAONwhhjA6j6F2tN1PmDUEeJ1ttHbSHV6nAHpf
V9+5+b/+LfokcAXv9lBPGRamyp8+f+pMli8T0/fXpO/TVY0kwcj2euRqgmJshA+K
EgigxWeJIk4tmh8rlZ0ee0ubVNfVWZz31AW6Q7gy7MJrpHen6U8b5E1dxzNVnq9/
i+zyZVxIlWOtGbxXMUxDSWOXTda8HIzHDeezmlN8+dyOHUgFAqnv/pwxPb0BBMlN
VPErsx5zWZPGT533vO/6NMofWLroBetiIsnoeIFSV806I9kpzfq6A+5ONHzhtTu+
eoZCj/4tHj93w1Mcz1bbLEQfbmnCUKFflDqAH0qmbFVLL4MVbhFSNcdQTnVL1/35
ns9pU5OrVBQn9zs+6uutIHuvILAt+uO9kOIffGxPnpB+MNcAxRtsXUVi7hOnHAlL
io2o6RAXhXezrtZXNjM0kK6UiQ6fGjx+nBe834QFB6vnPGq9dIi0btsoBHVkk6FQ
3oU2fLO+i4QAnKCzzVF9Ish2LqegKCyhwznlMZXZSOVRNavnSq4UHBDOrxHSpybO
jADAgY0q0+f44UFgMrESGk92/TLHwG3mHUamivx5gVyOmnX4zpVJ3Pi08YE5uv+t
yKPZTt/WHt2Zmpa+fc2JAAa5Vxf4pzVtAWdRqCr0S+pYiYL4XSqFcJW2t/i5FluX
rl9h1g2RIxfDWrSmNFElEdZ1rWgtic8ZtzueBaULHFmlUuuOhUp8Iw+l3I03XMln
DwP1vioMjUB0LugccfoJyOxKKGJvpfiDKxGBudjkUxt/h3iGLKjs9CDO2zh2/F+d
feCqzxlrjr8Oy1hkqLtzLsgEED+3bMyWMqHjOiiOWRPBmYL8OLrKJaQUopysdRxf
O9GvK64f7Vnj/cMqExxgyaYyKkloUVtpuzjZLM/5zXfSJMV5cOqBb6hbHUP44Jhv
ZaSMsnbbBOxgNNRv6VOHSXrrH7a8VAZ0NwJBzipkOiyMgVHvT4eN+0Babm/8/gmL
q//voiyaZZGA0bT2I0WWHnCJ3jUXt1bi1Eb0dh41K0H+J6OkakhHQPVaxzOAnjCj
sg57kYZIiOvUNxlQIOt6nIcqtgcJkNl+GMTpA7ym7uwvH2CF+r8ZpobdKhr551dR
48tIjL67mCmdiLW/zoY7Lj6Y6E6PyThe0Sq/D4vQkbOMhr0BhQ4vFRVI1/js/l7S
SDrwrViSx4+z5UIX5wzuKSJJgVEAMbE7/klImFHuxixkEr8GCNHHeW0iW3eo+7/K
qN8DCAcc0HXoyCbCagxfbygwoemdKRNOKWqHZwc/k1QhBWvWjs7RjyNdvdvmNbL8
KWY2I/9mo3tRu7W6Pu0BKBSTeSM/UyoDc5MEG2JSW2V0+o+28fL1mOhlXrkSm1Ub
V9FnK+19+RhcPxAtMguf+3zZC5pLL9wZ0ossW5XVf6fF+zG35Zklb2PHvzDu/imX
XainDe+Az/Juw0wK18W57UMXV4xCBTYZ5KvF3fuNtqESc9dRGK6a0D174hhmdaa1
0XX/qJbm0Nxn5Us5xdDYZQlh4jMjse2przAJg392kgzTzb00c4JL3TCvkQ177q9R
x3oHHAN7a+EUCwklx0EwiUbgu8gnOypJd7RYgAxeArtRHmxtSixmCBQ/i9siv7mB
jChEBlhHpmLUOoM10VZN3gKKM/kH2/Xm2vphahXAOCmpPIS96E9hVtknMTR12R3r
eDZGVUbFyLjoZz/b2SaKXr0A9AidRJBeyVEi9Zxkm8mjdQFM+IiEsXZy8TX74oXB
2zmSKAUGUMUYByxJx/62+WhzhMOuMnF7UuzviqBwV37bvgsWhkHwf3UV1FYGP3Ng
Ru0aP9bMxIXwkMQNwlMq3zW+PV71Y0kQhvvUUIig1rDZ01NLxe4TN1PFLg7+m+a9
YNJyWK7lPfSH1YSCQ9wOryjFfIsfUdcekbApgNzKtNmbXJ72Jgb0qo/H7/D/KoLq
cBPaKPUDOEAqZKc1ONVjpKuTamOsF8xB9qw/kjo97yUsK4/hNaAEoiPzTvmTXpry
Vi5l3sNwVElhQTVfT2Iz5TixJ890bo7+5ZWnf/GUgMqeESzEAlhMmFyLgFnvXHL/
4f33NDLC/UtxiIGBSQJX/+LraMeJ/n/CgMhfnTvKvDQsyGjzgPof83J3JZXhqPAC
iaErSOrzF2I1QQLYfLZwPPWyyYoeoAfKTaxmEOu3IzMR4GTXD2Kod5ny2wZeIGly
Ib6hAlL62VCAsG3e5hHLZ1z37IafWHHHMd+S2dlAJI6z4JS5GVyf4W4ITwzStyFu
IVWMYQAoiD+BG+FBZYJ3Zj2N9nRT0ZhNvCAMp0uo/j5/HVOjf6O/TllC5g7KK2Ra
OdUPMoqcZujpqj/sTDrQvwts/22jdX2RhYybDvPkuGM2QKvIULBYgD2QI7tkHFpd
osDCQvGOYs5vXK4mzLz/ECPWhV1dhovxb5OLaBWf/Ufy0lHkSoYVR9osgAK5b9Fe
eoLpXPtEsFuKwGFw7avzlbZ4TjX/gXHIOT5L2PFzOCjk5NUEptKiirloaRoTCEpC
GaqkbQwNqMNOjewsr0EYjkmZEaTyZuCDTxHSFEYupbWq3Bg2BTudxHByoRBSt2oY
oyjiHeJXBc1e28p0G8dycdMUGawJtEAEJvrFiuXJZ0iIoM2JAioEeIAdSdvaImZK
wF5Osfy4zuQgMd0Y5YAnqiJph9N6d1ToGuqy/vNoSqQRbgw9uWZiqqq0HYVK8ods
9WlVpEWNlj4h7Mkq2JuUxTlMzRsqYzOshJgiEXK9rS8aTn/7omdI9BQBMNiM/OXd
wV9nqzwNKMIRtakYX5C2F3mPLCDDlfFhPLbHd5HOXUz+BI10OLRpbNWjdDkk/RzX
PsZXbUi5Kd0GtKXpAyXHi0X425eUMQ3sQwkNeTl7UeJYyJGAynlr3JsM4UfIeRQt
AAjdnB8pAeTcm+05siDaZNboAig1LzPy8b4OcjgC03oa7IXulBC/pgL/DbnthuVu
NiZ0xwZTpd9ydtiGtMmJ5y+gohGWQb9qY8vHgQwT8tKk3kYXFucAA5v/QEtqnjlT
EtVOC/w67bNpJLpUuzI852pYVZafXn2OOhcThJ1HgisMU3IwILKRF0GbhnQvd2Pk
QaCFkvZ736D/Y6CvEl9xgAiiMFaxrA3m8kIhgOBlGQRQxuBPvb6U6svvvtwAXAYL
MAD5YqdcLwl4J2mgBKdcpo5aXNwjxUbFLYOF+QSKAr1cb61xZU2ECtl1T8YsGbGq
G8xbERGwbn5jdQCZgw4PsXsshKDYQuZ/dfOd44ZrBkl1O6gE5gpttREGP8o1bXOg
yd8dpdU60yJnqlVdDA10H9MWMXr4G6LEq0nsR3gZKgp4u+6Aa+Wpf4ciQL70c7C6
5WLaX544wxYqrY7xrWIqUyobtUvO9wHBLUpslC7ydru+xpDwFeSDOuM1nMGIQwwq
vDxP1s00qvFaO45cN9hF0I3GRy742QQrz95E5cRgt7LjhhBz5bFRkS+t8eIYrv3p
gK7g4pCNQAq2hkSH+zky767Lzd8TvNvxy44qi2pRnxUcldiNkFNQ/iP99zCWJmYN
7pB3o4zPQZZwgFuaOr51IUP5LsFext5b/RfBAaFx6kpEKbzktw51OFCnpZTnv8Jz
4a0u/IX7WZeb0VGVMFNRwnMb41nByxo9e9aerLqVz+Ehl1wNtCif+ilPuVjYqsaz
hEGns7Fit4ZHBODeDEtAyz1UweQthrh6k+1WmG5a6GzUau+LWBwqSrs+1CySkcj9
DrO7QEqqOLLD02QN+n8G3hbUCwS+hVclfRDVe2fP19fHDjA+9Ta7iX8W8XRvpk2j
UozrNwrGmfXjY1JMYwN2qC66pmUlH3aNVHUtzAhkGkS3BfYn3LunRTcS1zV+tPTO
5iqlW5+9kFcPIZLGi+Nu/0KqP9/3a+KD7o0/4xg9ZXPGdJkT4o7zqofdGCWh/5Le
61IxRN7LC2DY80IJpYT1ph/L5QvYnmHTgCPIwML5s9360JZyl4vV5Mp+CZ3FSe/v
DpWorbsHPvhIzviTbzKbGJNIIrXuEyb1SkwTKaRvoBHWMMvWupoXVCAG1RpzXu/w
BCWiczAYaUkIdMH34QSua/QGdYf//5cvHzHJNTJTqKJIyqiYUEuNJA9ZpyN1cl5M
N0aUMagB4/v/7Xp3n8yN0R+yX9EJe/AEt/SbmOCQn2TavHvNKVipSA2FqPz385v9
bff2XjQcEN74VP269Po8/LpHx0vIomtHWqXNcVti6/g0Rg41fVAIARRG4KT7rSxy
Lc7YAlbjLKp9SwBeHESR8s0CPyWyg49FzdsDH8uZMnnDjLY0aYUGI7HXJq4DBIpU
uAmS07Vmwn9up6hTz7i0r0hqwJzQvG+LpfzoQj2GYZUyoDSvUq/4QWBRE7WXjiGG
e2T5RpnjxU7PN7V0p05IVdnzyMuwDpLk2tZLGR5qR+Mc9TjeI9YB1K7jetIFOGuT
oU8+eC/ieGyumIxJDkWRCzIa1zTKTuiyKMsv87N6JESa7T4zMPWBbQiQnNSNXY5X
S9jNYc1xvytuxfJrEslZRPQW1BESRsWFesx1kPxgi01XEqjIzftqEz7lRf/hUdhk
ZsXghFmNEMvLH+3fHqqrUxpdMmx7JzmqtDFWx4WA8WvSYyFOlmYJ3AfLQnO3Wu+g
0Ks6HMxugQT06z/DzkaIXOgu4yi1dsPtA060nfZdq8c/v/ofjTUZ8l5AVqEOgNDV
sZSeGVcDKbk3lvGKvpuzKfYD7F/qMv2JRBrUJjfWD5JKLxvnJECa5PX8qw8M5vDm
nDe8Pe1H+41ouyoNge7jQNh6CbJH19+2umsithqMQ3i9adO0sj3OOHfgBSz8jDch
HWZbC7lqQjuTVoISQood/sTYI5/RaQ6D/DedzUEexsnsjK7eY00gTa810MiLGyY6
A9Uzq6K0zo9FH5ns0XoTOloqu8Cj70ghCj1jtwfSpWrhT2jPzeFFUCQJVm8kAMv5
m8Pnc+kS59Q2wPSFJj+asoZgxZCm5ZnyhNRMKpVuOrGdUsPX4oqhlQ5ZkswLIh3T
xXSixtCAwWxf2HpxtKU7CfEXnGcDuv6xkJIUpK8vOa4T1xYNXGmUMwLuS6i7dSlO
JvILUYUsfOj/czM3RFv4BNEw99Zeg1sFyqBVBqdYs9Zc2JEBUssirCWRyREGrSNu
VqA9qduUQMuCLmzGRZ2iemNOHU7gbmHatAwpA5l1rULZ+L/eU7JcrtBNFMRNI53K
LfDIeVYioJqfwVMKE2qalecD4lMkdKm4hKiZlHpBqyTCBzpfLh08W+yQBOr/+1jf
uk+zcjMdaHZ/8Ijbx0xSpn6NrjnEin2sIUtQi24h4xv6Qew0m6yvYeHSzv1vmZMC
V3uuDU8A50y9m7Jdjuadz5SxVIQ/D8Dg34zTVGoNAkJznYGQW6gShz2oMiqkhr5i
1u1gb6oLT1a2XS2LfbxETp0XiEoFhR5DuMy9fndYTJiFlK0dOZuORXcY+76sgrqY
aVHI9ZnVDs54zYzu0niB0dIPU7kQrD+qzRoKmmC1LobO6O8EL5g6tfL/re6CUb5N
RE9ZkMEgEgoPhq81sTT2PC6Lxqmp1HLrmnO2XfNmqLcqJm4hRPa3x5ynKQ6nQJkH
lYI7Uj1h1FWJobMd//QyQ6NYRRbzzfn+2rI10snpH4uChqcMVHw+tsPDegfJU3xs
8KFozvTn4teLgq1kD3izIBeqk5PepclEH8HX8CBzarrhTp6yb+UgNHX2RXbPrbWc
7bR9RLjta9lw7OwTzSSCfjaccwuhdrG/t+z0un5qLsJzk0DG9EHKEfIFR52FA3R4
E1D9XL+ljHX4hCnOnyvIMUVdmKriFGNR4tsoGwcW3GVX8oJDGDyKOotfMsSBUpYl
KGGeRFwZ4iydw9qRLjK3smW9lwHmE0R8qH2KNmjtD1UXzVSpzjRHkrUaq788+IQT
TAAdFtL7M8/yNTxa2vdfnlN1vsfkGIyUyAHGNUgkKGEQz0I0N67m5/K8WZOufYg6
4A+O9Gvs3C3XG3BZcf3zezwIbTLdt8Nne5ALsEYnSheCHEkFXdx1vILOfILM4N4I
Si2EkOsfXm5cCwf6/7Sg1KCx9Qvq+p5uxKh0nKF60ngXuuZuQcanttMV4pRz4Lq/
rLOS/SeFf36nHKppqt1KyUx96HNaIiS/KFATCx8hvUeETKcPn8H6BwK9KKRMD4rK
A9zxhm/4hlSP6h/0mgH9dYqIXS+gbwAvO+e9yTMyNGS4d7AspyE9swSMAbzx81hb
9ZN9VH/GvE5eSnzluPJPvf9C33CFmVVVWRG5VlYakwFA3S3Pt13FtNjEGg/GOODW
XzYrJUzN/DwhFkJucKH5v1d3Ps96JF+m7m+UrRVuulU9kzr9PPH3VN23kbM+ZF25
goJghOnJz48nFq0YkjFTtCDwd+5efdd7tDohwFlL9FR9MbEiHrn7uLQXD/bQlGy6
KVpR24IY1H3AFxAR3m0MMbOOroc7aS2XL1i457TVkMW/MAceYpQGnorolvD7u20G
PlL11qHTg9oeBGRQpXZ5s/Gcdr+g4nj4nJfUub8Lu+jWBhNkj82jsro39+46fJ8h
T3A5dcsMTcEdzIHrgvNV+rfYaJ8x2cV096NER+3zu6NaSdJ+iHs+JgAixSNilzTW
eHeDdSI1ikvw7gWXvlBMiixxFYAG8qO15xws326iJjIZ7YVql2R13iG56DqPAqXH
77KbrToD7+uRw8iZLPg6xkXdBB7weIPRU5twgVsbcJbeL18OVE+6P7N3jvrb20/0
tTNs/GV+zBjWthOpInv6c724Wlb/P89sg3N63NJ1wUCkveVkHxeuwuQPvP1L18e5
Ka1CKH/kGaVHFEGr3dr9jI2hYjK6J02MBdfOEchp20AOUr3TBobpfwm1yXH3lUDl
RB2U6LQ77UHCZatXBNMHH85r1ZHikWfUk7tMeOXujz5+Ar2WW6zstDeAuMEgeOnJ
eyDc3EHK91i+ffZjlt2J8c22uqg2lQ8CKFhs2l+hDUg3WVY6KBixTSXRY4v0KgjD
ACxBzqn2FKAhW9kieUcmwaaJn+Ifl12z4QeCyS43uMg7F1ee2DzvVEa3miCgjxAI
TfOZ8Xy8qsZjnS5ODRq41YU1RNnrU/gj1xLrFPwWerUROxRKcimH1I5BrxWOJ46R
rCmUiajQCas45dcsTVW8kM+FEQTf9uQoj00P+6BbU9GCIf89r2fZu4Y5IZUhD3Ci
27dhR1ts41nGibaSFovJjzMaIS93KdZ6BlErK/tpabufDlj+t9mlY4N8kV7TOeQz
B1PeQKOTrzhuc+//2hBgBm3b4QGw3fk/FkpV3gXENosYMcBfekphFHaskE6wGFGT
oCXOlXbG9PRZylTOx5rdTntPHYejTvpTWWs1rrejeKyP5fkPUAsNJ8k0L4r+xOxF
llnUxCVgqHbXuZgQ5qvPsFB+kl8jyJ6v3CHDZWganVeGv01EOm52eBXft6SkFgou
kdGTSeE2z8QwThESC+xN8l6okRRQ9WTHTUfB6YVmq4E0Ki8skB4DXVJg8RkpGNTt
vSowMSnOqV3YrcHHBMvJKXxNDKSFLLt9oSUud+PFqAEoPh+67tIDqgaPjXNF/P4s
VNghBhejM2hiOtCwa860+cRf4CUMShZkwJG9Uju2TxUT4ev6Rgc/j/WYIJf6gsvh
ax+KWIyVZFWdtqfmr9MiuKB/91Q/4hiSRYRykXCDVcNUWiK6ZP9Vdn4ZT4FXZ/Qg
qv3qKhD6NdiP0mh21kUq7oPIKHE9U99TFXn1IDSWmgVR8lclnVww3QxfQal7W8Tp
3KRv+K2MtZsWFMOspIVPtIr69eGciId+bzOe2FcP45peYlFD1QWzHvR2wI0DKyt7
/XENSYmV6KIguiuK3nPAVs4jnHurvYe2BjRxUbbMuUip1SKcMO1tjq5rHkreG06R
GHOQ373KS76LokqXPvErIHxTqUpzGWXDDck2xxsjk3s/F9QNChYjKm575G2UwBvc
Ko5CC4R/aJyksmBK5eMaj/6wp2zV/hrkwd75CUiEgx5PCJ9wyLXdW9QjqxvP9S1v
wRvWq/qkj1IlxGMsbYC3210j8kVGCSu8UysIUEMHn9Hf4xVmCwZZiboOgVFH+mha
T3MzWm/3pa5phbtbYu9UhL/pFsFOWAGmsavPCRDJvt+rhBc2Prb3hxFMPqR5RAik
2aTJ5SyeQvB6vL7WueivXgp/+2u1oMblkwmlllPso1yniiPAoXwb9ZdlkPd7AFCS
YKmbCfEcl4qdhenWcwS6ZO5PzINBFIOZxv94c6NZJNIbYdEzS8laIaCbthrJ1OQB
RR7Jeg0ZspLajWqO5jBN+uk4O6hGe7NOTT3XC96z2TWudQeM4Qs/LVllYkRw82Mp
WAR3i5cdzTI0OJj4GXRKrhp0OYdmpynP5pEMcQKAoYuLjoSLT58Pf4NcqvhhgVLp
YGpPL0bkV2XuSr9Y9sn4pcj4SwLoSlCZj6EQieURlQVEf8fzFx1Abtnzjby27MsE
QcgzO2D1jjjv9JehWyFux8yVmCH+GkYVJ3yMXpW6f03d6olNwbCiFE/1Ko+AXoW2
xSohGoZC3jZmm7cCbkX7l0Gu3JW9VevVi/2+H0WLP0x0XY/p0UgooSRAea2WvaF9
Q+OMXjXPs48N+au/kh4zJpKI8IW0lJcTdZW6C93nE6UcQAxZaldon7YEXNCJ2qG1
B3crX8uY0P4aXxywimiiQfvsn/NO78c5v0lOANBofsFeJMpxjwamPdEcxEbNHV0K
9xouc99xczHV38MFupnqIbMXvgfdoO/VHn2h3csarytz195q78m0C42U58ChKgNa
ftBk44M9rLN5HMSd/K3/TXGpIS2io1JGL+0BY+2UK3l7nIr0V1Mxilwqr5FRlBt0
5X8VcWOeuCwsLqDqeahOZHcBJALW+tzshPbt4QF4HroukGQR5lZDAS5CsBdUq+PD
kuWEfeClSlB7fPKmBav6kiLL5z0myFhvTDhniAPzICuLYYubsYmHJgQ37jnRAce8
0rem8gIjwKmi4ylwCrG8NMlTKkFPCV4ZXjG1q4Dux0f8HBVDTMZgZG+IuMLrf7/3
j4vgVgZWG+uTlMPs2qVPqEVOz1sKrVKhGeNe5nC7yTHPdXq5/5W/ser3AKTpelo/
Fqa+jQsbtdxFr9bPFOq3mnhTMqqtBUOYrk6PEH3+aQww3j7kjkZ1gRQDA0BLPAp1
GUITj+Y0clFkDXDAx/68S0G4ERoagtOKTBaMaKS2Gi3uBOSfdXlr9CEQ9ZehYJpA
Mjm4a8iqFC/evu8NhdSJuySnZXJFDHQhKEZ1HhWAdLo/Fa9oj9+Hlv+41RqAC8H1
upc0U3TCcLPLlwnw4lu1rbw8nZBrWCoRUfi++qC+1Pd6N4AuCx2gii7nVbK+QRMi
fdxyB+Ogvd7vUCUK7YClwuY8g+R5QpPrG39pmgW/rE8IVhF1A4M9t3WLEmEWG8Xi
vvXX4i5iVvIvRn/Mmrkyve8BSP7cGfL4a9ObtwWudD0Oq807b1R0nlhwNbdnxgLv
VgrZjSDT/FVzyeL6O7Rzq7oP1qB/pyrk7msLQrswuc96FdF+Kpu2PlxLTojQLCc7
4BVWFK6iSp1tpiXMYCQPI8Uws9Kq14t684ONoGYvlWIktdeXjDwSHrX5YL9hFK7/
tGcxQvwNArJnXyi+QvKEb+7T1rdQcDKYErQUVImRzm3azKciP8Ixe4PhKByce6b0
RLo7N6CWHp1tConxACmjRkqgn0KYI1frfUlvCVoDuUrtgcLGStsQ2poMKeVpyFEg
xaVGVzGga1OrSjb5Mzp2+X2FCj9PWAS+JSI2WwBrUUBoSPXdjw5FPDwVEWr78SAD
2SPn05sBNEBOaLkn/LVpblydawzQXjKXocr09ug/YPqUZmTKd/YCOtJpQdUgdxjk
7NlabaUNee5ukvC3/u6GpGhFGKPDnmpGxf/chcM0dxzzsuImFDvdeRbmiLERymi5
r07a6Um2VpM5ZgsCsuVQ3/zHLj2xc1S10e+IiYLqnPm3+z5q3cEaW8W6ciXOQ+NV
aZ1T0E1xz2RzEw8CGfSWJEWtRBTHpCa/9rcuo7LyDzOB0ktwmmIf7C1quhdlRzBF
xOpHpdqmCOQMOFInjjeZJIa45NHcxiUbNtfUHVl7TF/Rr7RC8BcuN1WEU9T6g3FX
UqAZiMAdbX60qx5Q041bwvNAXJz2RZU8xHyy68cf+o7o1B2z0tyiHdlV+VnBw6Rb
zBL36MtE6x0EPByh66+uW3nIGFLupnVc+kwoxhDYfuKbWFnrF7ybOGwPYDvFCpp8
NAvpWiP6u9rhAqeERA3NM4p4orcZcX2MELPwf9AysII/HtXV1UUFJk3lg6+SkFsr
nHSzZDzRudzEkF/h1LM6HyS1sx8CNS/L6e2NJuiGSpJuq6UMkodlatywvcOsxbH5
+k10UrRcMjwTTqmkCqYM0KfCRUP6srTuWpuKMjl4p+NAqaJzE5i1MPTKouOzlmxy
h7D9FpIPFCHFPhFjeM1+dfs6pYbUFh7KmXrA7yXCOHVMchGj3PKWxC7bA/4zIjsM
MCAHLs+OL8RnmT/XshLUzuaevqWBJ2+QQmQeGS4PdARrebXlHLuHaAX02EswYHTr
j/5XwJZiGPxRy2hyoaS3xodzPz1uV88sih/UZvZ+BBUe1rsg2L7K4wscSpaeNSvr
4q8NunFsqkt17FbatgI07X6BI4VOTIix5kmi4cX2t4Ua4YSjoTAGHtk2v32grUDU
Kb33KBemOmL/DVfvjkbrQOwcKdXfHci0vGa09NPVKRtzAHiQZBYXMt3j5J+cVwPy
2vfQwAhFzq/u312lBsILGO/lbVnKyTTfSc+b7fri9YtVQYwZdpV7lS0DWNn/xrf3
6AdCcmemuteKQcD1Clr4PKNL/KhHDQreCCOzetddzy6DnsWHo3brgsp4apqIsgjj
HnOqLQV9Jth3gPNgZ3sYBczJ6oorcUZ4Wy4LR2TAjs9RjooleIO3Y6zf8OZpaKZ8
NVTK+R0TDiBvU1IwF4kA0s23BZqSbTEWtfAHT2dxahjBHM1HTAZtYpf8nQwOQKkS
aRVb+ceoGHy6AM8m5RyLf8Is7f1x+AIHMO1J8rxRNnG+f6Hpmr/MHnC4lDKzg1WD
sEdbQFvKCLHejtIj0nU8ZqINdCn8FPjvP+sK9kye/YrEtq1KyY8FvtI9L3836Fkq
bS79NKz5Px59epiCADekToTIE6HLKp7zekXC1SWPELgDXH39B9d1O74OvAZTBTVa
0ajM8UCUT0b9yNOgdBsULRfoDwzjaSvdbJwednJqtQ6cCIMzZxoGjzF7fBfzaSPD
rgyihNi99fe8VyhCP9kHnehZSVKChieasSC3tAaYt/DuIxXNABHNG6m2gFjm+kcg
KlAyBL2iq0S2vpCY79vtqIeOs1VaHa02ON6kMBbr9Cw4aDN7isTYJapdu+kiKLJl
sF3OpuXVw1eULYLWXXJWIzbI57J0npbIDVPozSW7bt47J/U+zwy5F8CTt1upbO3w
0L7tOQN5ATcXb90n4hvD6xL/iBCpKLBX6/tF3LwWUF3fIFC4BKvQDGPFlrn+GqMi
QFmd64CurfecohbGt5CjTe2rkiBPJXNMsj+3uMqffwjIptycZSwwjXmrGD3st6U0
tKJE/++V6SKTV1V1a8Kg9A4oqIZUsmAP2s1Dpe5T50k5vGFQJmsEkAPO5IkKPw44
85666FCWTqut3BxlsJGO6iXLpZ9xVy6TIIZxoDlYy0Md8zg2WXdFEh/vCMsdSCQ/
WLWgWUUjDpfagCLyt6ZtKPh4PiTx1eN1pcYdvL1zj/1BpqD4N6FGLEYn1webEi2r
vRXHUuj4OUkj/FT24zTuYL64X7WWUvyTqoO1IbWLZdM5gQp4M0Vg+aGHP54WUghs
AH7TIqV00pwJTBbGVJ65DzxduuHCRxe0k+uBkyUUowkfzC5PGqxlG2nUqypiZJnq
EtjryDdeJ1keUQzQ3BpYWeEf5R/7O1bJaseJeBywW6Fn7IRnihhrFPcSHce+bydj
z4MAM7rVcuxFzLcvFGdmFYtCg0Oevw36uG1DyCwdFytR71wS1kWSGZxZ4yDi3SpA
L/zfRxP4d58RZ8O37njs3gy0hsGpcoMWDdw2UGQiScrnKI9c6AW3G5760pu66Ak3
fdLxXvmFIeePw0Lh40zT1/pVVwY9WyXdNFS1Hm5W86v1OYnZiV9kPIvGHBgewgm7
c4KuV0QY2KyahWXL0aYW7TjIjhb1E6uOHn/TWPd4ED9e/+s4qL5s4VMwjkwF4vqJ
/DS7OLbIUs/ZQqorTtj2nfuToGkqilM3aF1AzsKFlk7x2hlhF62qEAh+QAIQ7CjL
TpLIvQd5f+VbaqA8nua9k3zqGr1g+epJmjoumjbIX0GbRIDGYwQoUbJusVUXaiPE
ReyjNqJaqPMI7IfpykizdwmBVIGbtWbB3wpY3EDZBuLam4saGoqU4bl6S7uavxvx
4Azw9kioaShNDshkgiGlbRku59CRJnivHctwZ6w4Y092yJ4F4sNOzZOYP4KPGLdJ
4HWetJ69C2+3oodtiNW2ohOsSKXweGsr95p1lVEexXVRCHPLRnwCrbxGwg0kS2KA
gpqImSc/AZxJEgkBl+srQjNydT0OiEWTRBt/oqKQT+QtIMEBNgOm499S3xbbMWRJ
YMsGMP6iwslrw8XPNQR46mGqJdr//Z9ebw2cepuuNZF+lX6t3NDSSjKTSQUzM2Ht
NqG25oK4zueOC8c5EXNVzueo06eQqDSgVbHAUFJadkT2iITtu9D3r50PLNmvkZTk
SpkoS/3sBSUpfDbZHPfV1OSF0Jgqb+S3Q1j+qiZ2faED9/Y+0EPV42OPH1AAR3Aj
b3G81BujAzsNWMZWgnQTeJ2P4B+61wGiwiSHsMW0ohE7kBRVkhy0NLk9RZlQFvFD
QewpWoypdvqwC1fY/Wv8o3Y//eoW6RIq++xndBPiMfMBeE0vViqis1BSrcGYgcB1
4fSo8K9EyQ97HEebqGX4q30VFOPP7pRgmy50Gd4FUA+ewP8ZKj9nD/OQOECsqHRx
6pQl/fUQqz1KCyIqofKwdjRWMNJLFBrc2X6jB/Aywc6lu9sSYWT0iQC98FZn0w7/
gV2d82D1CcFJsRzM1NMsbO/p3mCOa4uC7Dloyfmo+ZpDW4DMWr6HHPZkfjBKuA3m
ODjf1CzBF9XZqWBiJ0/qp4WiA7vYdgXkYGSMtEMVa6VXGR5FKBbXmjh2eVt7qvJ0
LSts+Vn0b3EmobDb821XBWIqCzMGxwriXO+M3T2Sue8meCDsnIs2KxX8bn5EJduH
gPyK9IA141aJo+cYg7Ck7zgZn40UdWM3e5wqXbrlhW4AOXBlvGkqtOsHXVTrbLnL
tXdTuIS561o/tMUL7lyTBfgyqs+tOKkMxZdrtz7neHDGBFGo1JQB4UEuQG87R808
0HTEQK4AYLNaWIjZETLFxUAc1/6DJ64R0yo9alyyuCaGpPaWv/w7G63cKBF0CP0y
HkViaYzxoNJTHiiRScVu8V9zDbLK3UlpmqgGpPwyM3/D3Oi/Y4B+h3as1fRD8QjJ
md5NlV/5o/zpcHONpZTSuWE923gBeYqkdaqBu7n/4ncI7EDwRX0WbZ6eOwngz1vk
uPDQSl+DVixb85aCycTb0Y1J7lb8+31INtfvYRt3XQFTMBVDy9DuRwGhDomr1esL
Nq0oES3kgPQ/CrdT2Y9fN4x4aL/+egoLhB95TOJ4Gx8lptKdeprjhYDELxhL6hqA
O0q2tF/eX1BqbGVASs8PLGiN2bpLgCtMs5SfZvXf7fF5CQcF0giTiSmPMz54ITx/
k09aZNhdQ4jQf7izwemJlM/bMD6LWOynFhVA65f1c97cYuA9gi+2JnY23ID2O8iw
6Z7ZawUB20RHsEvJ3J+En6YEDl9chuPbM0xK9/HcQEXtZMaZc5YUokrNE49mkSE5
EmhbO5i8MV2zgoujYMG+cT0KiDE62K+AFUSlnKFEik9fvgqrgCGdJBGZn3G+BvtC
vv/qhkOFKUCgXzRnCBfbFGCvg145X7onVtwyU6fmkVx+7oQI+rj6oHScdGjIBfpk
+4w1FprWU1uLki3BRRh0PmVTEfjVu51GshmOMERHL7S+pRdavb8J7M+Oo36kbMzO
6kI7wBriRuSfyHuXBB8g+1fAycVQG8i3C8YuErB8KJgPafX9taRGy/0aOXooeVHY
yuse03693QpCwYz79p/aCorjeFYnRw02qsTgKttVswZfpcqf/dSA1NNn8X1B+QYk
df/m9tIp37jeLecwvW3Ktzbd1YRYPbH9HtymD6uZ+QTgQ17U4hBFAKf/jWGTNv67
SlidxPQ0Q5F4D8WC3u8OAXnKToJ1aIcW31OV1uMdMJ+0hhX1Nwq+UUrvZRAhKWq8
F7+16C7W0gu9umRhTdFUCjvXfshZDtmMRO37lBmJ0vHwsoBDdLVfhLeQzOxlQ0Q/
LSJyDjEE8XqqAfZlBPEJ97GCSgBt14D5sOeUSmFUa/D3zQ7p5QaB7ivPj9VGmCEA
rbcykFNGUsjDK9Q5uVN2/Gq5eNUNoFJmOrY+RnFaiCRjje9sHkZ277hitfj9EipS
5TYYenxraj81VbjUfCEfiDp+1AkLrOimYpaZqQPg4W3hGi0qWp5vDSFvH5VWjPLG
KRnvelhxzcBXbG6t290KJmuK8WD+VHg0lV1X/1K/5eCjP9m6L8CXih2XXoaQU8vc
VPcuy6WOG8PYk/18eHtE+FU0MUmoItMH2E98R626g+xBYw9BaYzAwXkRvQ8myOPz
b1AZI3WLZuqTI6IawFu8YUIc+Qruznn3SdpQbMgywb44DiDr8MOWtceuBK5Sp6og
CQCGC3VANmMJfb7aIp8lDDpXvI/+I77nA0mMRjkEmawXV13jTdZNz6OuPdFkoBS1
taXX1m8nanc1GZZ85HOsTgrBFCAjn0Ei0rUb7ZoRMDP6JkZ8LUBgHHycM5LTUCah
3yHw71FV3FXw/jg1IyaKbmRmDDpyomv1QBiQSJ52zml79c5bQZ/sWcUkEoFoLPrH
1sZS/xbshcWHH7sKMYp6+wDUBqreS5EMeztli1CpqWQEGhu0OmJ39Kne3Ff1bwSf
hdhyV2dWJb8+LAl/oiTQKsgmWT6ulGjvuMTCeiYEEISydE1MtbItm402W94zBfkn
aHPlXm0dUwsbzNm751whk2MKilSslG5V9NV52RMD6kiWc0bi3sbDb2YD9psdNZiq
JIc+H0txowQ1oU8hn1BNkD/Nm4BEz3GnrKuMXSf4eu3rfjvvPkU4ZegUyRO3kL1Q
IQY8cct+7r6+ArFjaQ7HKWP5JToE1FigC5n9N57qJTSTDjnIfXTnsn9CTMsC/Psk
T6b7uZiLxBTSyAnRjcnHuhrYDfT+sSKAGyKWyB1or07DKRiXPuOf7MJv3yZ2bj5v
MLtHBHuBoKDnIc4AcBMINFK0weqzEzYoCGqUUYDpNRDsACov+w+x5OEAYUcivA2B
6wwEup2Rqcjiobd/tTqRoy0HlHDnYadBaTV2WqddSvuA/FHFPXSqRrtcPRGgb6ch
+yc5jhkivOVc1sFO+9s+9ldEJADCvv2dciyadP9KQn5Buo7TQBCPfjnDAbwzAN0M
mQZmKWPg+jTwUSTnf8rjQelJHMJV5ebmeADbdediLfKJP+ciuCirPSd906342g3s
WSWy4AQmfGEdpnb5GeNhGdJjbWwv+KwGOPTj999KuKrYpDvs9If7KbR4w9CSV723
wz81TfYQ+S5nyQOrN8ufakfeodFzkPFCKCO+3NDnrH9Ck9vfluK+1INK9vaWMwh0
BePhh3k7dHUCGmcc5MByTb75TojUNnfD4NDjBaizCAO7wSgAJt8Q5P99ihoaEpTy
JHo6/8PpSKKdgnVu68KVIL5lDgytR4hvxK2nD5dKS99921OAF9o1LbabCLnPM1y+
6vVZTIx83vM7Qur4wGiOUe1FzL3GUhFNTXp6+UV6r6OwXXa0MhU1jHehPSJa0Qix
+WkIfN00jubs8jnAmZyvzGmL5FuYG7FbB9vDjV4J8pU5ciEoIpoxa6LY2GHm6cBM
sOuCM//wehRtUQZ6QGtFsQZQ8oR/0vjNWCmMg/qVwHFVEPQX5mANi6kEAcuJwXsy
bzfxAOBecHfbKdpFT6ZV/ReS2b7P+tExonzC8BXrM8ytpoZA0Q4zd0F4YZtDbZxC
CL0Vgw+aYWdfjmXcUol/rXqXsjjTqN/fjGyhezLTdtsYm8NvlVrxw1yItE7ieFmM
CU4a/xE4oryWFvJsA9gq20h9Z0YOKnA1LHha8xd8+Mkm0vE8m3p4bj1YnXRimBHS
kulgU5Cq88sR4vCyUyoMB5OXTnmYIVN6758p99RPpgHyQlNwLiS0M3dTkv046wwH
TAt7GjPCBqNnZtUXWN1xJXScRpv+Ke+UNr/anq3FNs4mSSFJxz6VotfeilzWfRjz
jC+e8B0qOdtm2GBAskY6gKjs5kvfp4tINODIW9CMmq3b2lYxRHiFyD66EW5xXPhU
0PDnob6xfA79JL/3lQdMvngFpxjcqJDwsCUrJMbzHpC3uniJ/9hYjBnKO38GzzOG
s0vFXRrmYFu729nQOOPgctohvQe81AZid32mLARyDjjuPJoK4fZUrIBK8CslqsSq
qRdiSlM8eYRJzyrbkHWbOYcgxrJfB9Fq2wtRWDNAqVllD484mIOBiY9VpcOH+aZq
eNOcO/CCkD9ri3m/B+zBL4V9YBmPn+KfU8QA6+cXlJLq6m9pNfs7LLH+znCjqyV/
Wx/6GtBCJOJjk+PKrP8SXRZya2vMJ9JVeKjw8yivy5G6iEQ+qe+mW509Hj4gBt9G
LAm2G+LzrFzTgEXaSucURpIIAJy2YJ4Huzh6FQ8eJvOjj3A4uwz6HIKPpuSQtEfP
/g5f3ZMjiZrT0TAhBMs+otMuBKPheAHbtFbOuuRXzVxHayhEWVkxIbWbUGbJslVQ
dZwIcW3RkhtUsSPRqBSP2OQAasDPp2gPC+lqdkiOsIIR2WxkEtTHnuLXjtH9pM/4
PMkdbVDHgY/8nkc6/gb2QpImWsNsyWfFFP5+awssa+6VWQDuqEE31MxdQvm8RPGI
AUzYD+WQAFyuP/0FxX5RmHlbh6Uy8rhVZV8+xQCwydDOo0a3uoiHLTsxXNh9yHVt
i3GcS1B+nMxAN5uybera9OWe8NK4cJElFR1d6vXBxDYejTT2HxTJfW2yGigGxrfE
DpPTvshF7lL2LvAYlRkKjSodpgI37ZtTc+RIj37ePXLBuWzKvVc0WReuBzpuadfy
NC1/CviN6l3tgvrvwAN6zstKe0uIJgmYNHhVqHZrWcW/alMU9OY/So3J+ZODlPpf
8sY241rXeTF7XbjxGb0c1V2FcSQtnyZI+8c/8g1bdykYB0G1zLqLu/c7IaALFP7l
GnQ7bezy31JmTp0/L8/O2pD2+tZRMezjinWda5uO4itICxKtpDsEZ2IO7kVMZxID
RTqeYYR4dlJ52gNjcPbb90TEEQYR+Ig4DCZ6HFJky3QcPsPo/cmGNKhr5Os89LAK
wSCYF9pWL0FwREGmLZbwSltlFih415VQM8Ys+V7C3TJy6508DH+Csw1EL0xNgHzH
JUAuCkHrMdRCcu7c2Sluy6uVJWYel5BG2kNOoXLWwLhLdLxUYc97YdAMyrmr7EZg
CtAU/DhytyN1aJeHVS3ydc/bKBg7SAHp4FzlhflvH8t1m0tbhQpNkyaWwFkSwodp
4N9QoArtJZvgPximnUi1G7TO+qgqlQVqrLcz9U/JvSeIeifag0XRbctajAsFgC80
Iz4yEpT51uEf287mkk9SNJEvnJD6JNCCpDH5c0AvoPc1g2+fCBYspBY1tX7Uho54
pdG1/3HYLKo4wRaAIujGUpmeRS/1NlH3E2JFkhq/JDeFaYE/+wRKDMeuMaUlagKc
/aERohU6y0q8d0LwSMcjK1RWoOoSQM2Hvo0YT7WFfm6Uxw+o9YSrH6QadCco8QrI
o869r/EDas3hkIMhDmWY1MC2bL/YERsMoVvTUYLq7bedjuFTyE7Vd1l3BgZRYs7a
qFb2UmcrkWOT1j6IKQuadT/kgdZbNf7Z6h0MRW09CogyE/sTd1aAPN5h4UrBfKN/
KveDhBNYgEfkGCQIIgS5YoO7qejsev9p9Au4fzXRUp5sIKN59h3/6T8xlAhfdnuT
c4VlQjsh2T3AHgtf3h+dCrxLKLqRRhID5mcxcS7tC8h8O4HZAn1J19nvSLwsOMDH
H6IwOo0KQ492WSDL0JIX54BPsGTqKKIYFslIjYv5sPXhsqrrxHSLF4DtQcRuo59c
kNe/Pu8cf/u54r9+yFs2ctmvA9irHZMRnILnF10zELAZkSFMnGzMPyft+pQaD+Y4
Y5Z4cS82CQFhjn0XuFKRsaUTUI2lTutc5dv32luCa+wtU/nQpL5D1fuhF3e0j3rB
qX5cRNKRAYDg5TKyK5wW65cAQWjJTOHi42yKzyuU/fHxwJ/GdSZ0Ux6wLXE3Osx+
v5fmvnNrfzPQ7/OuU5A06Gcp+p/WJwOHfedpw6RtyMVQQyZ8mHBYWTRZkYjOchpG
FtW1GRUZp/DCxBVLw55IQYbcraMgxrpDg2eJyUBccrpGysgVgQCIJk/csIQwQQA8
P+URMq5cRRb/VfwDTyBtTJ04OTI53eC/x7cexefVdqAQCLfTz32VyIZ7UNf6QLrn
jY7TfpSqCBArs8EdRuHTYFJzikwstcu0URdBJbM13rT0hz+XtHee5dFzqo73QxbA
GjtJfMeLb3X1SzYcNdm1C/AkmzWeEd21rGIg7w9JgwBC86Xw3iO5Xqawj8CWwbTc
WnxvRr0D8JoyCm/0zpZm696AigkMCnD/mBd9nx7gcG/kvYQG8/qg0uG7IkU3Jvo6
TTWz46Z+8O6ew7GOWlrlNLm4B3tIPdDfufKlTPj581GxqEwv9cBv4KH7IyA7RlgR
53GpizUUn2FXII4zd9PZNDT8hHLUotch/Wvmg8ESCK4F84WvgTEhPFICm+1BWLRs
Ur0HJYrL1wGu3c2AOpT/NOef43pZoYJeTRnSDQhRfcTFTEnlwCFSuzZe/CDshdnU
wBgLltkeAwW0MZ8WaDFI7Y6xsCoqwo3CVgkfKDInoUfVmMnbf+ZUFZlqr7seEWBL
7mq9rg/DA2hHthdVPWlxqXLQbyiJF4t/ZXpEBmX94HXKaluvggp3HRT/FrBcC22c
DI/jslOqd+9B1SBvPQQtpMOkzmeWQYa3mYUhY+VuAtFVyzqEn9FkFdmOTPE3DHBl
cZ6/aivxwEVrEarMI1fuIBfhCm1+W6untX9rfo7cFuoaaWj7VGJhKSqtpy1pB3Mu
ooAdpOuYP8NAn1VuWxjsabKD3HVMHS8/UfvR2wmPK/1E1Nx+WIeBVAWjaqlGbr9v
eTnXks/tq2Pz9seYuulxShxP+PWoZHk+O1z/y3oh+eWBl0tGRvrSoU7CDbaLGsnn
hO0gaTmGn2e15RHtUkUyjaHxvmc4LQo252+zdhILFFFm/Gp0PnRfJw1DWuFhHiU3
/FIYpNwkOo+oSk+Cv63eivMTxTmlGuUrVzfvxCPCBXIXB5c2LOSNO/6RI7n5l5ta
NsRuewLkgYJesQ/3T9Y83RUww4RtREcSxJdvLVqsnOOoJcpk5OL/TDw9WPbnsZSB
3VBzrZ2jpJSAaIXCS8U/fVXRnkjJnlry3f50rQMokmQ6xYsfsqorxHOo4Uj60JBU
reZE37QC6ktGwbrjVtuCuPPkmhDgFlFLtsVlepYWZAom2Os1hx+akfXBrufHkjTN
cyf+R1BZyt6JCSyNZOTAghkvfzvGvP7lWEknSMqj39YZGswPRUnq82YlR5VRC5zA
QzEy3+BLv8/+GwvMkWlqpISLfMW7UWDIL5zbqi9gNKj2Ndn3gZ4+INnCs8qmagWR
O4DnWZCY0ReCLyxEIijonvX+XLPCuNqA/uYqW8JSZMYTqAksG8dX5pv2bmzu5K9B
iJ3p9orRU0Vc+YPOepboQqPCZ3YtmXNRvJmedtW9mRnuonWEmHdG2M/4uYcUYVj8
wN0JXdXPEJGkb2b1+qq+4DB/mZiUJRdI7Fcar7FM03l6aeh9mxOc9zxcIJwCqoQ+
3CYynTg80RFdvOA2fvtwYCoyGLGyTrT0xxUlOUvNrQ/Vtld62KmsJqT7sQ/hEaux
GzZLEbEjnP7EMe883fqFKey53RySzFHQ7lCbOQms2JoWB4SrOWalKN2VjtDc7wS2
A6KpU/jAJ9SYZZ0+Cxaw/47VhYt40oI4tUHBvQ8qAn8BrX+7zhPMwL4ZpqVAvsDk
/C4lXs92xElsGAx/XuXpVI6WHw4yqJFYrxEOcL8hwVroqSwD0t+YN/IOSHJUVQ1B
pMfhSsu/0mf1BMBMBHbQ389LnhZxn0P1zBiemiRKqj+8dBPu86Z2XXZQtFHev4Zg
xpq3ClOJsrAtFGTPUZ4cMzS2CMwEKE2g92HI9nAITGP89RXOOUXKKIc2BY8ejk8+
OILKPf5HDFKUpyMXizZNN3VOk6xvTzJh07gLR9W+mGz6om1ybPN2iI7XJ01CC7xy
nytsu/9uQLcC+gIB2Wj7PdIGW3RH0Vrsid6pO/rpQAkJTZ6Ej5BoTj42ntMJ4cBN
fGJZcY9Nl8aIXU/p1NdTUA6EPe2aAJqWnUfOmtpAp3VDqjArCIYUQCcS6BOBAqaG
sOunKnsxlm1j6OV76N+sWhGWNol6q937KfDxG0+kImiTWSGTBDdkob7xqnV6MQnQ
AR0uhHg/cfPiBg3KMLbD0CYi6CEENQ7dc74U9DcKHLdr6XKRGKUtSDF+DjG4zZNU
wZvyum3GJNqCbiqy7TGsBIncI31/TtlX6uyD0RbL+ElBj6tC/LmSheQbHr4Qsu8K
bnGqJjaqh9MPan9S5Hcj29GcxGdLL0qQxOsmGeawTfJFatBYyMZZNaPf+iN1ylZO
RJ2Ep57vMOTcj1Mhh7Mjd0CztbleaaDBz+ryvU2XPqKO74rIOw17DpFu+dmitTTD
gpHAJtUDjuaBLXnUCt7TjB7qSVFh/87JihKE7GXyLJPR7qVdPfP+UVALBJmy8ml2
qobDXNwk9WAtXp1qWvMrlXqwFBE/BLQIIk3X5naZBUdleApPOm3qoeMMX4eBCLeU
j/ttpQK0bPp8qzXJL8uyfh2aarE9sMd8PhE1QyLNgjT+Rewl79lrSpDEacWFzTCi
ssD6gWQW0HFRnpBwn73tcAjbEtWPFbote0M7x0CGFa0pWLA1/05FURnZPVIIfW28
fw6e+996YHeTPjbozeoHo+H+Ch+AudVfSEDQfHV3Sps+CEvG7pMIiR6vP+NO2I1l
MIz3dgrCtuoJuc7RtfrRONlRAdXUOBLBr7maShxczMbw47OTq9JK4SgFZVgEb485
A3JNjybqHNK2AxpL9LnGv3UTaOKy4UL9qwbi44fCosdFPuzhqdXWQPrmmPtaVbpj
yczKyF/FqjgWwFfPnYopEmdTjcpITNGIhkI/tvorzk33oLS/3HsC5wynELLNlZXV
wAJ0/YhwFiflgtTakL/VgFLlJSz3YYJgXKj+T1RRDZLarrDIBf2N9KjJARrvUNbn
kp1AbqgJpfDo9s+kusQlHc4Hu34lUTUJHwwo+U2tfovn2hTvhHiwIxyFHF+ANcpu
/aBOJ/qWoVct1sfvRE4cooD4bzywN74JNRLDWimT9KOtTIB3d2yeccOXKaEB81d/
CT2wOj0VUFm0KxWWM/8QYmtI1eCvdgmB+9ejkil2vBqICS+Y7GPzyoQx3s0KY2sH
n+AzgIsWGfhtMSmZ85748qzKbopJAITHkHwmQPb227nUgk7Qg1+VjbiKRiRoS14t
ZtupkqtKw+porW+Of7dckxbT5GXi3joAVogoCD7bR7I9aQvJ47GtvoHst4NC3kly
LyeTN2UCAzJ4/G+veXh8pAk9qUxVEQLizD3LziEzcOHXQsmnoWaO9rb65+mjplI/
HuObqssO+iEodZIZiFxYxGzsnBIG8+fxxeZTjhW7I4xl9zXJ4Onu1S25eWHwFFsL
zxkPXZGnUYFP/WOH7sTmfJICpz6pqwmPCyJbiyJRobGh+X7RV21AFpPelQmlfOvx
0oxdbeP030VlE/u9vYbSWZzdKKCEku0N4ZPm4yS4YWoC0iwJUODFcI/gdistQEj8
c/MR7R86rwRYF+3ImGZqRBHsyw8FCnl8+x/DW+mJhaqR7aM89CIuwETT/2j723BU
oMpKjtZnEgZTeUIwDBSk7EP7NOWq3Gbt/4jpQl8gTaCyjHMPa+6xVk1oIOYfklad
rtCf9VysZb/F2uwtxMNBaLu8uIfXCkVnt226+Eqvq7F0OhbCJe10JbvPc6i9LCF2
eUxhLex4w0P7KZwEusSjWUfvDVDkbdVdb0jX5ZYLUNyJCjT29Xtel6p6boXRMR1R
RmIvM0rzvHkjuDz2Ho5qX/Ly6jxQmxxAe+OSFDclAZv7zlorE07i/XFb8YE8BEIV
gjzaczFkdbJP6XZuNW9dp10JZI0BhL0BhWoWaKu+BzwAxQ3JK2hKW83cNjWJw9+6
K1oBQV52pJ3zK0xdq/+I1U7OdQbezx01jEyUwYtdRpstCEhD4Za5Wv4ipLtWEU/A
6skInqFhnAvnoErJTFHbdYN9b5MwBz+AyU9DGnkR02kiM4Phx3PFriKeuiF1Byk1
8Xr/vLbgdzlWHLTa1oST1wDn4Av+ogVua6jsY/puP3QNIphHM7LZ3q1l4U8p7gU6
UXnEn/0WsYdumZIMf2VxVRBaICKrbUffqvbAteF0VcQXMP0QOciS9X5nLDvlaKg4
jPeDBIEQk3xIZVuQ/Q3xZL7X8mCEGw4BIglk4N923VSEPHx/91kUDyXyhWey6rOu
al1t3R573NLtVxBGsbVS4EYOnLLlrPrRJMx1hEnrmGkCB016RJ9In7rC1o2UiB8/
rpPruO/4/LHn0sK+PaJf6c5Ve/SMbQSFo4WYW91sJVroyO4luyjPqXHSwy34txYC
sTMV/fWOQv7mPfn6GtkMGc0u4/RBbCgMiXVHdm75oLwztmO2Szb5G286RuxOUTu1
6oM4JXs1L4o9ZCIcQCQqFakkpPyo081nPknTyS3n1Mj9Rdsa4Nvv7MSxiwzNNNwm
6NvkYcTD0Rewg+BwAUdLgsc+Rbnd8glSEiI6Jb15G5X+pva6Hytuv/epcrh4o8UE
iQApEbL+M3iCNmbMhf4i2nqs1PyWlfoODhRUmz48+cCsCLbZnCdS1m6i7qDmiM/k
q6TJ6pdvjSG9IsiHau3QLv8dDYzX8/00S6nm8L1jpNbURHK5usDceGreUsBIUHAR
ahpIQvZlHfrsicIjHP4+s1lyxK+sBMcWNSkTZw+OphfCxMhRyFYCSJWqQMxR8imx
rwAkaGpDuRhUEnEo694ovDXJsGCsB7O8j4poBnhMUUcn6jn7SY30oEahyBDmER/z
VEMnyoOXfXarNDN/dbREjuRTZemEXvcIJHGbfb0EE7viskaD82j2OkZ9MPYaBn15
dGmSN3pJV/xIZntsqjwm+F9acH8JEaR6/LzOI9FNBThyPLJ1VaKHOyOwxcigswgc
t05ITzxPMNaq68fKtkeMxt0vALt4+ZC3zF1S7sBSmScDsKQyQoYD9rR1aoadyg7x
AMa0Y2xLOmLYKnM1pFYY1Rv2XS7G3CDqkoS0qZP7dhdmjM+oqmQN6qxERa54k/j7
+0I+m6LsFQvT+9kt5WOIZ2rxglfDxM7j/qdGGoBJ12b9vd1KznhNteACooWQdOjX
h3XywySPq7NRfrRQOzDmj/deMdeuYTYrXrBNwhjd0soJCVtWb7aV2LFE5zfysiZZ
beBrSIL4YDLoHWLYN0yWWwajz3ZpnS4Inrc+7EOTTXYDoLM8qPC0h8p4f05sOfSZ
nB02+yWhij7JwBWoSrnz18PHrcMexbYRWYR+BQEN5I7StcMkS5tW3szum3ALqra7
USqIj8RE02LBsvO1YKEThEVcUpZk1vt/BWOyuDFbbnXeirqCT59ABKgIz0KtSffl
73hlvUl4MKUwvN4P9JRxyJkXWoGRCxdw3M12TKcwdWcJge+xstpSxVw01BsaeeIS
qpmFbZayjpMgqj7uGuJma87BTu6DXMXP8pzzpMcV6zgjyQB/tAX1ReJtqAtyWir2
Tu0HJHqzB+1Cu0XBUMYTlxS7iTPEbYhk8adscLqdk3F1C0CdaOUoWL2M2P2jxk/S
UhX+uZARcnGFc6qQQBbQyL17cFZ9oASOcoFbSfdCyPBHFhSLSvgw/wgKx3IHefL/
wXaWyUNL//JZCZj3HO08bxREn7hXlERyf2Gy87w44jz491EB9VRaJa/tSCZ1ST9Y
EbF+NcZJPXt3YrE7+HCFpalGPo/LLqbOIOngNSu5T6MilSZ20+C/L0Irt4ZN0oxp
n/S2UOYSczr1efbklTHt1qZVGGw3HvQE1F3kpxYBtaEUDooaQSqdpBDRgOS07hqg
MTnf2UsvwttyH1D9egFzUnqxAhWYoTy1DLiqllK8I2Mis38/5CrwNlekgC2SomWZ
UYqhFGXZ02SYX9oaAXMZ/E0+/u7bU9Kabwr05MB4cfS5fqVO33jv50V8lYSEA3SC
X0vFyCWN5fshw4BoXVtrkedWuvErsDTLg9RX8ZiKKO0n8eZtOV+k6C16vgh1vtJu
DqhxzaD0d6NDfBVqgSucx/vZGo3Bl4gUhLHMELYWgPb5ztt6ODe/CGdFC1nAk6KX
XKr4Otqw9pj8GfRrJAUJbVRoYhvS6hoO932IpQhFBUUcm6eKMggOgrtyezn5wfln
LUbw7p/xPA4nwNCyPzgEqaCTvYmBjecLnO3q2L0hLV9BePvbwfhtRgOPcJbGBQff
/A/m1AvrREysSgts21E3nb/uVgmHZ2cgen0YQKf2PsiqwO+OWwBoObqvT/tOMVr9
luvl6KahR/PJSliGVvPrmqRS9QmXQVWoQnYEUcKMNlN7l4ZY5SK4UnQd8XdkKuYE
pjdC+31zlQVRgmDW1dn/Yn2AlnejQzxUrLPxMULUlke5rk7Q5Pd759NAgIc4f9Ue
YBYcksrggvDzcHACwsxlx6cjfqvAc3g7VSrPjeu1UCsvbM9yg9kuFSbfiV7/A5VO
jgxtRH/x6G9VYHEg8EKDeJ/zk7Lw40YP/elJaZS9RX4hyfpuNsPtybKLvj2GOo4i
iducPpoUDDMkyIrau/YgN+Sz7Wr/14ODS81cvjb0r7MylRUYblHF22caD7/g91GW
aUwqgQZBj7DsHxn4esxRXUermJFJ+SwjlJuWAVaT1xfLlPP9ylh70agp+qC9uRjV
k1bIYt8RQj5pvCAwYIJQ8jkCX0Gqb8EnnLGyziKGyPCHS8mDtWGuRvH6cWcH+JpX
xVPG94DPqpPKHKbRRgMNqQ0Jj/U1TWmAa3TcXnd1Oy2kdv1AHJev1zQf33/I1GLQ
G0OIahroOEbW5Cf+XfcEnhF7/rd81H/5qpnOt5lAoh2Z/GoZnTVveGNDrBulyPah
njM3Wma1oj1QNftUpfsPBiMeuuwPVVD6U8iMvhdmlYqamL8uIzFBQzypOpNqB1X1
SqsT5j198a0gdxN7lHWReFpDqHaRJsTHtkxlpsYnyFrWPnRJqoBbMA1IuQ/falzH
l7XIR2saA789OEjNcBxE35XHClYjUqCzS57avy0P974p5ZHkoCmiuYCvC8GsSaNj
1KHztF7Z8a8PmSPA9SE29BZVLuLnmaTqm6rQRY0WoUEUIkcOoM6PRRc0XJuY8sYG
jO5036f+JG+8Mqj7DDU0cXSp6zhSD+ts98TN9s0iR2oXa8N35QUlx32uAh50FtcT
/1V3OlCfCktMqjabLHvtfZ3UqFzlGRiJnTJoRdtv5dkWr1v58GIFcD9aHXdPFPf8
BajFSEOW38Ca03SfQU2LY8ZNDrZXVm1dReRDOakWSZgxqKPtKA1K6YbxBizuV3Y7
0MV0bkceMV+9Lp5JXqGM2QXdOkQw/BbXu/mSNIOcTAJJOI+Rm+BlmYgpKPzLh2Fd
CmIScF8sl6B4Xu/xeZkYmDO1G36TSckKjVFvedByBvOTVemeeAb85jgs7MruMaTX
+zmYptPIThBJMyS4F+21ibHk25TotkM2Anxpyj8wTpjRhJxmswQ/CU9jl7AAh26f
R9t6jeONj8hu61bpXbsrIj/4rilESK5cfgmfjEYSfyAfPx3Cq1aUeVQZNxsLAzKa
NhmJTT5kXvHLUNdIDVBC3lrO0PkQXonAJqYoFe3PIgxPe6O2OO8d9otFfd1JkpXB
Gfpgepn4ZEHvFq5As11lN5bz04TsBYxOmKeYl9SoM9fEIq7X7Y2J6QmbTsqAdruS
Eq7OHzzJ6SmqBCUAbVLisciRBd+FoTtN4GQIUzZRLHs37W3gvbbI75xe1YT3AYIq
Q4GrjFYKS3fTGZmPh26XYOq8ngQiHUKM80Rdqgp1HheLe/a0qY1XLR3BI9kFnMHi
oCWLEbF5h9PXqTb/gRp+nZ1moXhpiKo1xUSsGgtFd499DivJYvUtF7WqmXun8UTW
sCBKOsGzWsSuNFFVsVdRUBeeriqQjhl3NTfhSxMJ1tdHD0L7PE6tEEua9NV5z58w
zxaAChzRbQt5ImE12GRdcOGL224K2gFYN/6sNvYGaLQSX0bqSusIqeC5eaiIFZ33
L1WTB8MPub4lo9Asz1kh0STajSH8JXZCYBhlqVlb9jWc/DnTxe0LyBL9i2oC0xXA
edPBZQxqA8glP/wtdWzWqurnu/Kpg2whBwg/ob92MXf1oMK2FD81s3UM2Yeru2wL
gGKPN3muaMDqgdhPFXPZ5VOVawPB64oLqbZi5niSOCLKENb0NslJd8gxZiWfERMz
vBpFg0MjNgn3LDYMKQ+shwzJw9yJEt+2xQ2pf8IxD8hrdAauwnKbtt3QZYLT+sBl
eqYgsmuxicPtQ+wrDi9wswYH/GjKa/rU/ddVq3PmpIEQbiTxcHCvAxm0zQlK96Dj
obFKjI4QcZp2CaAc0zDMSFdEFsDJzzDZ8KGMqN3fiGqAUV2Ust11Tm1AjJxIWp9+
c93iDOaPlQ49U4/cqjQB8ahqvrYDC5V/Zqr/DHwZC+U579fXfye8ifnDaYUK4Uvl
NnRhYDvBBfz0lZEYd1547ndFoHZ4bcWb/Prme0zMiTDQErkJCWAQ2iRxMhx4YNvm
VvmLsOeQds76t8ztpN27dFslbGFO37nekvMFr9SgS+n6rk1qO0ivEGiilXov53Pt
zjgtvDwCyQMXOEy27cOD5M+/17JD3A/Dzm7dIuy0Qnx8xHgJ+5ucuKwnBV1TorJD
d8LO+CFjJ0KWrRYJ5YIa9fzxfdyAA5V/PvoeI7lLK4v5qkq4p9ykZ5UjHlgEtTeW
2VHWAj9dI+CiR4fdVnZIyw0Ruzh7kXO9q6ZqlMexq4dbLdGrCH0oFCOie2ZyVOY/
yQ/gzOZl4X84xHEnF2jgQOsKDdsw+jMH0EwJ3TPnR4+np9tcL8tt8ndF8DdqCk6L
rq2gmE55XPDxgWcaAsZV0SaH+1eYobz3ZAg6PGPGp5s4Eo2cygllFI/a9rcHs06Z
ox8+F32HsqkW1AqoOo9I8UqvpXa/GJPvHLyNKAWdB8FOjTpltDShcUdF/sVoEhC3
9ulFZGZcE4yUXzxgmaYf+jGhuoJGBdJ3/r1f0128c35pjFBenyPAh7N2u2rMD3uq
Xd2Scns53p0IYwZrhFdxYWru+TGwc5o/uO6vyFs3a9p0LZAkjT0iOsco+GOhHuYO
OVsZdkpRLSKBkRBSSAz939FK3ifJzXRgBDZF4Qt8qzxB/5sqdknLrxt9anSMfe4/
KcDY1fz7Mwsp5Fz1ZQLU5XI6BQPR0uJswtg61Uw9MYDi9D84juOClzNk88FAbA8z
cUwbVme+Jwz3Er/FlfQKQYinv/h/45+eOg2Tq+uxNMqY0P+7ujcNm5B0/HC77dsM
FwFJ5Lrcm8+G35dFALsLMFg0soAvcZI2UNR1BHWQ3PiXcwGPGrm/wHu7SGy0n+ha
7lyFpTG/tSlnrV0SQjICmTF6RTVH+G7Gg09EL3lvDjlA3PScapyrAakKn7lVZYxf
p6nTsuwRskqQa0U68SPZVdSSC/PSw7hlbJj84dxiZzW85yjKT3VG2LM0glDi+6gv
ExsEDUipwGHDrV2dXSl560SiMJzl/aCLDPuMz8JPBMnYgLeDH1/tcPOp/UbBb7t0
kyBbdJb96ebFhRNfMfuKtgtzT/v4uzTfdHMSO6+xPNK0EZaOWsucsTXggS6cG774
2loC1Yg7Peig4zZFvhDxAXK9wHGaI90jUe5L1tqqGSLVwgaSE/GNXe/oau8h8vLy
pyeDpxqWm2R98HO2s21ilR41neEA6V5gXQmPP+xAklkcrBJurfNCB/LkJ/9YhHMh
aEIUNdUfSdA+UHtPIDLVXTTuN+9nXh2t8q9PluvAlNrPLRp3gXKPAgzVgEFWclPF
ds4moexo6ASJ31kTR239Dc6FunKU83PGZg7yfRqqcBqhhIFVb93vnSNzrF7R6o3Q
/veVWNJLw+Wb5Jqh9ZU4IXLXoXaQ21HWOvIsTZLAJ3HOm8hR9cNQYkEuByxNXvML
dIXDDacxGVNoPY/mkwXcawdGCACRU+EGTqfd+971DquBBtiD9czvvWlEoWT6p8Ec
9c7f6Cc/+Gnpuq19BP+8lN8G7vXapz02EoSAFoC3fcz+ksN58L6ZtJhCRg/lxdT8
+f3QUrNrIMXciHyzFFDDtM9W16bOqHqghWD+7tQOia5C1mw2ezQm1uUXfB1tLyjj
LOqp97K1WRn2WPzVHfAJlTZrXKT3cxikVuD70vCdNb2VlkTCJNBfh+mnV/R6SBj5
AttI3jknp8BCnMaQtD58NnnP/7DS0FipAwXOs7BM+u/wrrqflT5ryLEIXePiKT3c
fTBJnGV48mE6396hTDNwJ+G+k7lk1corByhbW98B+KptXlgNX6iAsEIutvRAuIf0
8RTQreluu7oTzDOM5aW6BYS8jCTtyO2er2EgA0MmQK2mtzBgN77sThiNvi2l5BSF
0TGOqXm40diVWsYKkw7CSLlYfDSl2J0gCZ9ohE02n8BVEEv61fGU5QU9Qgc5UFYe
+0Wvs+B4BGXNNievOL0REEx9q+8EdBgWoTbqQz4n26ZfL964JKvlGi5wJWkM3G4+
hV7MPnrED+Rw88be7Pw7krznuqCxlzxRFpyiWIw/UECWG0aSUiKoQs+drpk6qGg3
+zVqNsynUslaDC2LuFJd1DoD1KparX0n4TVMtX2439iwF5IvsO9n+W+ASau4DHXW
yo8eecAKQ5Gw2RFJgNr2DsWYVM2nJr41gg0zMyd4cOaHQFZaoG8+DOjJu41NQ9M5
wyE5G4IrN5he0Hf2bA2A5d0a+9tLiLSc5PaHQZwvVMzeRVAwnGTK+bcCWZbSd7Ob
cR9JYJtJps7pU+WTqB/V8hhavXYRERvqvPp9Ja9X9sVJjai/Z4xEPuMEMVxUIU77
MNxYXwfJFy9pGlVRuMR91zImLyYIwcqc0X4ueBdE4C4BfuENdzc6GGFIzgOd+5HR
koykJvX5YXypGA0gq8/pk4FtqL89lh5j2qZuLDKrSxCo0ABykr1dtHaKr4nzMQGQ
jRnRXj/FqbQC5lUmYRjF7o844hMyPk0/cJVNY5sY8lMTYIS/3hMHrVM/KGoXM6jj
zeqOYMXlH5RcLkJ++mlhK2EAW4YG+Rlndyw3DcvFd5fVebwMdzk6R1N+/Vt9D1Le
CG4oJT5nFbpRLbqYwax+DUmZ2rNG0Zrl1UV6AN4vwogWBeaAmdRNFauLUKYiMxcs
3eXOTJ7aueJ+EDfgew3h4adX86wPc7Qy5Wfm7I89k3TWZdBYp6dl9nPxX5ZJ/oC1
3vCJvemMITvqNfOeMr7GYqrgRxLau56wCMKBRnZQKPYip9SR18G7z/kamQm1lo44
qBfwB6iSudd2cv6W9seZGaisg94Zx+Np/2w+nySNA+fFfAEiZXBw7N7m4TI0LHe0
KTsIOfa5BqVkvl7/RK4KE1tJ9j6U/Ah1eR3SNdqB/TPS2gpeRMNLN4InG1P9YG32
m1sAxY5WpAMa5Xux8fyGTLyj6VDeUe1dqAVEvIpbA6jarcmNOfvFAiIzhvp2ruGP
yQTaTGoOLHzQu0EDZu32t227VFMkKBrOPmaD87tAUv2iNon5jUCp7H5oB5/wCuPP
xQi2WwMy59gD30EtCoVOxYSv6plWw40YjxeXmC0yFn27VnVyK5eJJuCG7nl2RHUs
fZNobmdCpAkcjUJItpvJmUUSkbfyjxK3i6Fs9bEtcEpo5aWVk93LAYLvrMEysFvb
tkMoXlD8FWDFfe9Zlk4hQOnLNI3t4Gojn+quKRyDaIswddhj+IGXyhCJfa40LqRX
Bp75ZVk5OtCdqp0TlhGeYVzizhpJOawk19QwtIW1f3xFgkYU31f3RJ6YVT/JTX6P
zIYx7ugRsHh9/ZqSBVuGHuNrqKJsZpOA5dpVgam2DWXj91i5WS4G3yU+cLfH1KkV
JG4urDyzfYXYhHPf2Tm/QslfDXuep45DYgHjV/ISCfb/AoFzyxEwKvYyd6kMuiYD
flp/GFG73xVca7ZVl0Olk1BYUUbnYx2dh9sUAUQkpUGX44sctno0w8zXqszIZ/Og
XTRrm98+DdurfAgQcKVl6e5jtoQBfX7swRYNez8DpSakbYtyoqjSDqXbAEpT8NW1
nQN/yKUtLQfu7cMfAifgklQnR68TACazNr/2YeXYUCQlo0brCeCrCUX7TP5JokzD
GMytXu23/51iw4qpceKGUW6JDaYibzRZO/iLoJzcbTPOmrQqPKBgkW87ADzF09BU
QVyF8+aeNgUWW6eSPuoQ+W3lsNjR7nrLBOX8qj5C2t+VyZ8DkC/qu0Ux80xmE1Kd
1grZDElNM5RuuBKHhq7mFm3grOlFbhcjvAoeTkSbYew/F4/vRALonmdn9Xgt8Ypm
94t9kZL0QoQL6V0phBY0FKtGUNlZq3b+UAv9BZgiiTCmT/8XZm3wniTYGIOb93+b
ZRrCRX0v9aZLuu6EMB1e4+cLv8M9BHSOqq6TdNF1YST549sn1t4pWej042CutC42
B0gw+gL/JoRSW7zId3IZF312BG37N/tw3yqmnG8TkAQl741EHRxTW+L/LtpCd58S
Gd+2+wnF9DUY5PJ57qW2P20MrOLbOuEgwmEMDDpVautwJzVQFXkEQrp74KsvHeKC
xNDL6Y+KAArdBxEN/pN7cHMfzODaWZi11m+R8HhlSBjfO0Rr6wulmoWz22gazNq8
UmS4dHgQMQtT9qcJI/zhmlKnTe2kLDQDnQc8DS7z2vnsdUaxk7/nzi2FzhZim8Cd
2uoysf/yrJBAlXGo/PCAjiei5ZrmqwLAtCymeqYZ6sP+zAuEKDX8JIRf7Nv82at0
vH8xqTNiNP1d3xJjCEZEAphpHom8Ck6uc4WiVc7NoZy0eQTcda+n2pVr+lBPvq1I
/ud0FaBJHqm1heoePITMCSr5ikWKTAnSRRKfzp7i5Ku5DqFmwB3wydFkPnpMiupm
TQsV3QSOZ31FEAsbENaPZdzuf92QA6AfGzAJsltFW/NuqRHxai7IRzpY1GPKVAw+
WeMBYJ6xfMCSomPE0TLgraGS+Nb69CCbNEYrf8ub9xJ1sslNZKtyReVA6Cn7GfH4
C9hDHAIT88+5ZI7NI0RxZ1c1jXj2wLs2qLrl+TcwPu/cZ5wNnf9364FAiPsnUILo
sNL2gv8nIDttG69+2CEgo9Qog73SxCwmqNoIJt/0e05c/wYNiOnjcUgOcTCBjD1j
d+VAkJDfsFdDxzZ0pQd8npAsSKFvQXYd+RHEDFiXMbEKXaYzlS0QVWasRu6wjgbw
sN161HelhGSaEYJ8m3JfqLn5ZLpmDtvRU0AvyJET/4UZfpQOaEuyjwQNmk0bNwQn
MkpHf+1862sLiy6LoagfQrmXYaAQdskc4xd+QSSe8AoB+pZOEeYIx0nUwCc2pfZu
fr94uP6ZvkEyfjmOrR2PNgHByaXgsBbkWp5bpTcsBXEwsz9DvcCGIw4TIGTB/FTH
xU7fmm1pcpdMr/tN3MNFvLBE4h0td9se5fVU7GNdx+2jISleZqofhUmdW3hZHzP1
KWTWobvulwkOEc3eUoZ6nu62fpvVeLYFcv5+s2dXhe7pRr2Lwlok0i/beBVWMFEw
ZpCoEYsYri9DTnH6HpeKsR1VycbLoKBcTbU432ZajjUx8FCF7eshnxZtIn0hEEZI
LJgcUk4ikZ7iBtK3J+FguR4d7lu+M8tFw5xcYtV+RV4vW/pEnx2R0yUJqZZwZRfF
nS7ygPXKWoeWr70hH4YC49Z5rt9Y8PEBGixUogJ7yzw6QrGWS1Ch7PNKUAROhW3W
dcKI/Ieh6XnzJNEGs4y8JB7vcp2C5mAKa38B86EW/3tnYnUTTypyMFthobS+nxZE
HoeXxJMa0biTN3jEGwCFTU9adJ/4d67/by3oX5waSH87LlAR7x2RR9y0UVMN34S6
hEqOUW93BSU9RbU4qbOJOsDpbzG60jCYKtHxAEeg+u90r7akLyZxTZ+ePKzMORI8
XDw54kuZDAA+qflKlL7B5SSUOdvgmbPhdKnJOqBGWUdll8kdTbhCKYVsC+K3CIU+
c0SmTZwYHAs+Ok7z/LpfPw3mODnELbFmXTrVgfJeQjv91UfzvINKepJExuRbiOhH
XB3vcnRCHfpHlQL7+/5SOJ0lyigaUnwz87OfcvgA8HZNUTRBX/BzgNMQm7FiEFDs
Qcm0eEA/O3iKKk+ZolYYomBaiVzkC+Uf158zYYF1QRgzfJaZYKO5sEso7rDeXDCC
Ch+uSk3ydHLWSmojLng1SMHCAhNYjHVWL7V30+jqgZDj0Grm+ViH1wemfxMle1Xd
wrWb4p4YOPb7eA0yByE5j470j0+KO9K9m+pQmGbgC6rz4njKrcIlH0p8tJLYb+Sj
prZ7zE0WE6WO3uEfaWNPImCSRvl5tNgJtPVmM/yz/s+RI3TRw47h1i86hJOhzV2R
57+OKoAv7LIpuuDRdbCICc5IWyZactbvlVDmAnJn/B/JstF3/w9yIYaScGz71jL5
L2jERnR8R4AKcNivbSIKqoe0Su/DuKDIcdRIEMwYCnoK3TxW7XbFMqnkMBdkbDR9
Ybmr+IPBZHzBfr0Z2FSvSYbsXiJvHGvL3qJgaNzpUfzeUL0wgSZLuLF11kxKMLCT
t4qBwoGO/HeuJ+DcMDhmm4lOBUnC5HuiQuIxGj14wyeTo1MQ6nNPJ0ps16jxEUgF
DcWQBCPOBi1uPVAJZL16+FjuvGCk6swMLHVqxwaeS26fVQrilWAumg1pC+A3KCiB
OZ4+tO9Us3jkwPgsPXTwUNyv2xFRxNJ5+GRNY5yq2MxXI0g6otWIzn6GM9QX/bpr
lVIONR+z3Fsi/P2Lu69r2W5iVli0A41Y3ogM2WOuFqROnO62AMHJmMnUUF1NrSvS
EivR5ivn3EoRrQRa+psuTh5PEn/5Z55KF+IPioTkICoDzTo5J8YFrHwOTuSX07E8
qL1GSEo+2bDex5wm7HQaC+AUXie0FxnYAljuoZSZlAlxWsO9IJK4n7OYbHxc6ft/
ZRXdxL+gJgPatoQ7OBYrPSRjHXgANUR24ozz08WQYNBfcCXay8bsvNZqkCxUrny0
xceDJ3qpMugLtL+sly8iqEfRblK3uVnUAuNVRXIMlF18f2Ie7RKY0lPcMdXEO2Vz
odn8ISvl0kkSdEf9S62A01PENWT008kwDoIxoySx5bus/hpztSECGKZnRr8SMN5y
NTMtn7WKPW0f8Lg8SaT/PKTu+uzbI7TlmnJZ11BgEQt4L+jnNV3Wi+4ZGR/hNNrT
MSeVxEoIN8CGP09J/KF4oLAZ01fT7B/gdHs7Wylp5YOGYC3AowUFdHJPi/LISvls
SfI5nesR0N2HLdEk7gKu6Cjx8w5ejrDdB4rGGDTuwpamBxYIwRygRa/dprIJmBEP
i6sS+FtBmhrqHH/17XCYXfOmqFjIVAgtu5AA60UNxNNyeDLPHXsg/VXBCP40norh
JQ7LZR5yDMKAoF4xWb9l+GEKmxZkM88LHdpCibpZdXhES5FSgzCdpyAnZZb2fAiE
neKy34h1vzbssiu2tXbh2rxedrT4i14QjlFLZ5jJhvsKfITmaISl8ayM+HMrKKqI
XM7y3lPnBbmNfvSslV7MgYPbW4pJXA8+32rSjxVHdRWAgmZAmkDXxCQwt/iG75/6
kqOdt1tj6TLdL0JBRBnOrbPQLlMfSjxKFMQ7gNeoiTzXpqXuSZLJxoOwCQnb6IX3
0lQDG7zXm79mYcGEy6gkiKTcujhFqiYZoK7/bAlHBVCC3A2yfMbl1KRembG2kPzb
zcOooQd4K+i/9C/rUMwJMHyJfpincbZn4mFUjFYGirICoDrV2SLeBNMQruvkQf0k
VfX9ygr6Mji5/soPwiWMYgqyj8L5OA0Zb4S353zETw3ew0IzwQ9iWXsOrwAd9Qrj
v4prmztvAnEzMzwUn29lPdLTaH20B1OB+NalOASp1/zX+DGZMcjsNV020D6C6z0P
fDiGDpcDYWQySrdFnJIzdspC1Rv07iBtiYQUxyUf113McJxr+gjtxsoQVpAzK6+t
C/O3YrzfFzRYaVS8XpWIzLIWr79vrEo6EQjkFlvykS9hSAOq5U8KNbNZzjrlKqPv
ftG+0vy5Y7GaNWzPaPWRw1QYLLzmwejAHhHDrApZ+i1tE3Dk4FcpFF4lCR8ZSiwU
PHHEq+NzgrDciZ0FN1Ce3mr70O+2ZOw6lH6MppkpH3Wcx6VUgwR3T91dRanIKLDE
ajoYBFKZ7hhyxFD3ZVbyzaVBRvKKVfbXabRqe8xcRmcEp74JvhfjGhVrGXMLN1AL
J35wGfyIeNBPIerc9ThVGuoXUcTWt7rXU5Ejbgr92dw7rQIQNnhzMdYRCA/KEZbD
kvQS+18vEZDxo7TbzsDSbQ6PwVZONrillp7PNd1JUeTA90B4c6xCsh3d8H2NBxFM
aBJYdq5m/g4Vztav/p/ojjf+aTRwh4zLvhstqRHKAiVg0WCKCSZbqC2odTgKMEjG
sfqBtk2u8N1kUKro3+WEue39EG2k3s/+Q5ojVH3grTYufIievLYcGLnmzDo5iZ9C
wbDZFcHyo7lUvWmdNDtMC6Ous/IorKiLOjx/TWVxsr9YtCP3TobfcZLjrZ4XVpGv
R+x1teYDg8TbNnyJ0GTq1VZJF10P/wDyv5vMWRj+VY+Bv04HZ3Te5mm/jcioPFIs
flTAC2PPs+ZcJLvLcVySSKES8F6GtTn1Ezig/sPinKynBBURA+NN8KMPN2xsdl8d
LEve1WCC+nn/b+bT+deOx2jmfxbCFTuuQwjEwtEa/EzGLrsJB/fRYkZw99A4HaE6
CmpVtMiYhtDj0RPW2RgN6ptJQq8gOd1p6z/FMyX1jT4BYrdI36u/wKeIe+Ap0pdh
RLNV/WQ4mtmJc5mMj5/iStRInwhtE8cw68fH8AVPSXQHKtFxDOTnNctheDIzjz87
zOcah73VreRGYaLYL3BqfVwp7J9ANWGW3gnCE6BOoQ8BiQ5+mkqIkFQiveLzKwLH
I6P0cLdlpuDceOg6W1qxzZCm10Ldmgwzahp1bHtZucIaq+ZX/dG0RSinrryCtwgf
AoZJm4MAXBRdxWC/Hf3RJ1JKsb+4C/Zi84UtlfrVGi8Xy/9eg8SO2QsLrzW3YM4i
UHIu/gttpiW8pAiYTOneHqhiahUSImsYw6k+ZUZ5M0RXHfnBO6SqzBf/8Uz7PehS
XAKkT8xXeru3lYXBwmH+Q0fkdjETjnPa4RgE889dSow16IYouvpUvhOBp5CF3+Al
V51HdPJba5aV/WUjdb/O3yehlbgpK1VSs//f0j5PD1zTzzD3suo/cf3jPzKlrTpe
ehbXRZW5r0n6Cc60FCJ2eSDDqe9mY2IDjwTIdRJ8NmgbgRp1tVY+NoDhzAaVgw4d
s/1ZTgzJAprAmLrAZ8SHm7+dIVidOG+tx+IehgJB5jOYKHJG3fWz7+/D4XQ8fX6+
uV/gd3XZah9d/uBed4NH1Mh+NyVNQ+9tuFb+I+Gie9LjdQf8NSxxyZdv+4n6l+hL
UN/+YJRJyIPRBhTMhAtC8Rwb49Pvz9iz8hPhM3AVvrSBm9sC5PaOhgkpX9S48B/u
iIpF5/yDnzsb8lKoaW3mZMrCLv4R/b0rBJbit+xvgOWP+EH6oDVtDXJRRdHB86QF
AaIwFKdWS7FmksiJOCDr8Hp5LDMeRs+vzG+B6WC5POIWYkSNYqtCl0o+cN4mmOQ8
gYr7D6rvtdgXhwmaFkhcQTSJmg9TuOGlqfErt63HBORxir1leVmaOyV3ZTZXG4gq
91gHfQ7r9VxmlnrrtXfJKI+CJY4n8PEmRJbpmBgKyRTvhRVFHdLVZVBnLIfdfnuk
9NbyjOFlGgj1lxby/pQNemsa7Cmm22ZIVQpxT+wlYUBOn3faN3+tWVS/DHZKKPvP
//0N0HyJ/wv0Y5i9HC8UdEFVNzZYq10HcOtjuZDy+J8wK1cDRNbXiTreZD1+UvW0
4nmEidoLO4irF2AXf8GkLHg3Jd0+dfpXH/YBxQNPoWvxJWey1Jt7w6mShS4r6Hw9
vYultEve01lKlBzRBAfwd+sUV833Tjh3o+eX8dC8xRrx/V5KcaZyLtK0SYLKucwt
4tFAb6HzH+8qelO7pOzRahvk+EU47Gwegt8iocNo86TvwWEaEnHdEQy//uJf/zWB
tfYkqlH9BBhCLCLva/FR2NxrkmXY045rN7WPtNcj/KWYg1HavBPqabQMZwHqjC3N
3/FugbQcGapn2kK4a76bGWjYzr7GaKNt6IkLNAJo054G5H/LvTrUi+hndfCy36GR
kxf2ZqHdfZBnk6I8w7b3Pkr9C3og5meTwWZqf4G6u28xjNcJQ1A4FE84eB3138l1
W+SrNublq7GUGxFo4/qZwAE+JI9FPfZuBPXv/7M67NF3BUIreUgFVSCvpiYRiGXD
9wTb6fP626FuLk6r5ePjanJTBk/fuh8vhV/iD/G+hAOOOe7qMQc2GwxfjA8AyoRM
uAH0/gZ2aNSX+1OvrFN5L0LAHRATb1hduNR4IPdysxtydJ7zxiHFg3n5icZae398
9SAIXqYivDmCwJG4SM6bfEBHrdnNlLVQJXuIavPW1WqNBw9EypYiPsiKd6Q/wTr6
qyjLyPsN8XsA4Fb0uQK0y4EevV51XRNxL/CplM6AMxFYPOeIXTWtqYnv4XPHxJtS
i7QNWZx327r9eQ6JMtq5thNF+e2Fbol6cgLnqS9NRMXxOnoUYiPz42qDI8Y+TPIt
8AxXrOARAHyRDVCEM32JCj3BVnAezNkG5+UMnqSXVwhJodJRW8TSsafiwWKmN3rA
QlXEbBl5fWjIUr8hkj2cUnmDvg/iaouAyUw/A3UUKfa4GtPTkrmK7Y7M3J2qDLyA
3cQHFnDwAXgmlkthw7EWI2291aiZoH0QPeWg7gtFkg2UTvJn0MvceOmBJG9BdTij
y1uAIElv7imcPnq7Fc6UzTjpIW05AUlKXVIdrrQ+Bvzt6rwvu4fRE7Iiv3ajUyj6
yEXUAv2kFOli2fQ2RaPc9pVguEQE0quGpLVdAni1PrAfNDDuatI65HQY6HP3BbWi
4TcaNYfOpqUDHKeAmXUUOVw1gqDeVG8I0V0Rn68YgsHCQqNna4GVirfRpvnHo8XQ
1pSAprvuidfnbXFCRluIV90OW/PJogWURPC9xwb85JfP4WDgUaS35LRiVhXcBUwP
vDeWlAuwTQGy1HWb21X/KwOPRjIluBUG8h2BoIhQNXNKabtIq2hfVQO8AmNf5wpf
9zIN5V90+8IMny8/cplt7w6pbMdAmz20+9Lyr42vHzs1hBDa59kZ10q1mQpJTUpk
a3g7kZUSeqrusfdCb1PXn9nh0q40vocuQ9YaIGPjH+U5VD3l2JZxEbwxVAAStbmo
mo6oAiknGJEYO6ZDfqQmfzhd2yvoDiAMZHKvH46uRErJRpW0dQReuKyQO86chcxN
OgqlTBQAN0Tc9Opf56gHOTFpKZbRYeavqxL0YvlBTzpdoT+jYE+OxuPS3P+KxUtE
IArn3drjVfZvgAxJtNHfe7/owtL+vDruHQvhqxwYWEEBG3iTfuGOPIiNJoe+wg9A
0S3pvm8t3Gn5SP+aTQzjjttj5VQwBGYWakF3S6XpmUIZc63t/5y8TzD5bq+A7M85
tAVIv4jR86lAjsRuPkt4qA5Qkia52i0azp7yJ3G54WpQjuA/LOzoY6seyQ+yEsI0
sz2u0yXJWvbWw/c6QoqZra4SQjsXTWB5soMAsrpzm+WMRURF7++O/ZczhawaKMN0
4v8U/Pw9xlIRWDpgfChni+R8T+PuFHmANy6iBbyFOymyCrAySs2LRoeXGbtBQW3n
y6PyriTED+JHiZ3q+/hlayg5cL1YQLdnydPNGtZA1jZFmKSL71eibO/RoOE9B1oG
YYiSuv43iIQ16MfcQ4WCt6lfS/E6PIYizslocgoBPmVqyq2wPP7EAUgScmiRF/YS
eVxoXlAvSsY4AClhMltl6gulAC0V+lDSqdKM10h5opquY9O7zzrlwx0AApMKJHrk
0XZF8av+KDereVHS2GEsRRgJxKyANxNWvX00J07WqmXooeV3+7CxUNZ5OTKqNY2p
9iy1gVYgnnLu9h5iSY7/ManEHsRDzNZ3Ux32PN0calB6Bz4OkSPfiw70t+tgI/O/
Nnr8NdM5Kdc4fjfvuvLavhoKbTHTNKGVnxxd4/sc8n0NeRLcG9DNQ0ukwT90THv/
1ebfJmm3im2gMpKPEk73g8V9z/lxzyP4NXznXhHCmDhJo+fb0kbNVgMtY7XQ3eef
0za6kOrEzl2GQvJ970qEcsRukRmuzJedlm67x1tvzdN72THMzSz2PTh5fAhY7TAO
TepI4H9ktgFq7Zx/DpsH5T6lTtuS2vrezjcVWh6QFSDMxEK0fhJGg6jyZ9Fds559
37VjH15tZx5PPNXy44ruRDtV4qlHz7ZUQ3NZlSIEbsnHSfszaRv90u7NqBawtF+y
zeyqjIyiHmV0pUOEgEokJOKjL+xYvPZlSPX91oOunt57Pq3kX1/+w9jRmAOSinFZ
whIezOlI1uShk+TqhEJcuTnIll1X7jqMcU+8AM7DcDMJcL32sQ6qtcdXD5u6yq4Q
c/67mxwg8rDH297OfKx56y4QC2PlGXYeFWFhuzQNkx3trkcBwurWhWJv7nnr2EYL
m48PMTuHt8CILdGuqVuyp2RIa6uvq+0is5qBq1VbiRHCKdCLbGOhsi38tpng+rcB
0LDdg/zqdHK7FACAPBRylIn5z//+IoMJeV1Dh5dnNARu8ZPvdefWoacu0MHNUf1B
Z5fHlIW7SUhL1g7DxtHRPH3uFjg1fUQlNUqZ9CR4qCF6ffuw+jmsa/P5OQLRn3/P
Nzh7Yw8pq9EUTapQq7OIJwPhPYoGtmfSGvP2m8X4AcCWm7TIYaIyV1XhU8wE3WkH
27EN8qW+oSQ4zxkrLqOgnFt3154JCRIzQAemaDQXUdNO3I3C3T+GKbnqQwJ7za3D
Q8RWJGTBdHwm4LU9NXxq7rPxPhVrnqb75S8PhWqEt6NKqFZFqSMdv/KIVANlOrzZ
DIQ2Y2ZSX9bdZ0KXy5NcpscadILpi9cX5Bp+eQde8C0MUMYTtPpFtMgLvJYqQyss
6T83vebrWxa4BRrykQO8l3Gn4QJKw66oAqybyHAj07ABC66+CdbfY1D75kRDZYlO
JsGZfjWe5Z8H+iQmVbyJznwhN0qFTavM4N1z7QsE0T36uKMiY4XezmAFIeaDFyCW
dffRo1rO/hnrr9VGbMYypToWv10OIy7D/QPgHA/w7HHtha1rvK4R3ywo4k2PFEPW
rASEe3Q+iT1U2p3eXr5Rld2we/GTAW7Di2PVSKO3fSzSmqMwpYSvNK45YM4qxZaU
1ZLs4nB5jtWRhG8MNRfRp0EMcOZUzAp2MqOmMELPkafDOFpxXf0srdoQiNd1WTzN
oah6nqsfyqHZMnIEupc62tUH11zB+J57os6+ct3xSDwSuTbHndiGdYURRViL1b2/
MZ2ImZj/VCqogeTN7kZXRdnjfo/ZNFfosg/ZlQJ3nJoKlBwI6yB75WU8HS1eVVTO
eUC6o1oO6PlQqXfrPL3YSFrP6I/CNVluLReKwzYk0iTvR/o4VBL2FIesxBa70miv
eMr9yzBxpUSF3o5Z8Ju++5de/Wf6yYrDw5g4MhKXDAHP/a16/1Nsjh9BbIplybo8
gfTcZvKc0I9pUN2rFXs85oNNnqMuRArDHuJ9QDAcYOLegc5zrfT4DeDWjwbjRDXA
4FJKWPIQVIFDjFZpz6VBH24hwM1OM3u4ptni219IPTBJd+G2ezZUrb8D4SRZgscH
mM3XNs0XLxSauS1Kbhz7AZc+lWG4HAGh2XKYN/Ls1OsprSHnwDjHJ8bkIWv1mFxo
UwzxLDQU+9Pv4zjtaXwSt1dC9R6nT5cSEb8x9w7LTjz7qBhMgHjG3ne7nhMTNFkn
lav5JtgnRCfkdnuvMXu/X/ToCDWv/pBRDXlgsLj3nX0SwZ0uPnlsRkTem/sp+HGv
EX45PsNKSBWoGO3YLh5d5zH8zQqXla+lkJusLcW2Xl6vKvvNWz0Xp556bHeFJ5i+
+Eq4TABSxcucS6wAfitxzsNklquOfNxCCZIH7Sm57TOXEMmaey0gvs5Asqm7ZeNR
Lch7mKvZALQAJLaq93tTud55xWpeB25ho7guUJZxwdTukGxuohqQ7AINtvFPNjIu
kCbQD4huxIByXCZAoc3829gmoKhWj7Dk7xoGhgDCkcdrNRjupcJPqu0tw/jyuGP9
eopZAvoc7pyyFI/t69PrGks8I+H2//jo+ONZy2r/ifzkbf3AE1z+UthrzozAyRL9
FW1uGRyZ6hxYuxdN7QAL98gopCEgFV1x0msL3yoP/DF4g0/vFS9Gu/dKpcAs7hrM
v1Mr/uq5PM18wwgA5tcycerDQJQsL6BHunIlYD4PuDvV7G+NxKDvr9yY367WRHeA
OkRBSsNVggZ7PODvPXMGen0zbdatvTJYSBi/gcPaOLAupJrkbJFAPeC4pJXtuQm5
U2X7MM30HTXN0Wv64JVFG4AsdkT05tkJgNg6+D2Tq/vbXvAzzTRQ93G0Io9HJh9W
e+PZegO/g10KGaS6QZ/1PKnQzRuGgkSpWFYVvHADE5AQ12uH7b1hzWbplRruLAl9
mqPkn/cOM+rqQ76BYtHwcSfh7L7LDh9XsMDCDgMENpLgrxuA4+u2vdc4SKvEne91
TqTKt014AJ092ueejNjgwrCe27+VrXm24MzLxae94TRTyh7RgSKkcd3iAv8MkFNV
LP5hO3MypcShTaMy2egc+p3a7XQ7OhYSZ0oxJzy9xfFaBlDTkdQKtX3rVVebfJEN
i4cyHqcqoKr4bKQ0jHy4vEhNu/O2b2DCS2EwLDuNl9Mxyi8ajH6W0ncETMyfAjlX
gRg30C/pr4lU1zRuqQUfTB/CGN5/RpTSKr7Od11FLnvftIzmEX42tZW7GOfkvxVF
Jnt6mFhdMW84cjoBHH72ZWMkVsXX/RjumXyJtgUyXwXvWHQQVHFKpOdr5RsogFkl
mUzWa1gnLs3wbSTcYt8OigcbKO87m1DtPMNu1QoDD3D7MSQNEICQFX9CTT4CVH3Q
W2TEUdvO9Ti7A4xVaTyJylg9IRTdujkon9kA82hk7Wj8HZ0pP15tpcLPpegYtcYw
z0Gp4lbcnBtoYrOaJJUD7rsoJAOSJG3LHREC7/S5KDdXhyMXXex9PwBiLt9yytgS
6cqvO8BOblkLyl3VYDONTlCByu83k/XZLZdZEdcLyWkfnI1AYMeq+VCOenVaQ+p0
x8AGE4Te8QNZ2bFIOD0iKVgU15bTa2w2ueTQSoiLXnx8g+Qg6XDSv0rCrHB14I2a
dvIAFOyT9j6+VIK2YWDYJ0Tcth4ekvFzD6M58yjcF0wGEBzZxLax3GSpR1V0JIjX
ar3LLhzPvCWY+B9VI/e7/cPuq+jTLW3SkPR0HjwtHpIilSnaT8WYmF6Xle6ccvAx
1qDxnDvJ4zn3TCqoVRGKppDg5De7RNLPG6dDCf6enlxFTUuxTnJLOtSIY+KGwE5B
h/oP8RFY0ozT/YfBgxsNJ90xzqoaNWvpm3rbQDymDZzARf6StWPMyAzcu7x9BC1o
uMbsaDU3crzhfx/ke2TVi7oMMvg28cG7kERHq5H9yrIG3WzKQIQ8/qHEZP4wPV9A
Y8rH3FfyLaH5RQGWbOT2OHQkFRx5sXgEIA6MNbH9yfKDnpxFqc4rPQp+hiPkjT13
HEblYRZZLkWIFmDkjn5eagc6Z/KVUr4hpDFPoiAX4JRZ8msO5mrdd5CJOSfuypDj
mjNkUi2Oa0f6oL8gb8+WygoUImAqWLOMfkRVWcbLVV4B3FzQjM+XMMD8n04z1PT8
Y0N9KAST3HZpC/aYmh4bsWjCs43ruX/LETkdiy8gRxHfL+FsKKBQxiKg7PYmWQuU
woCsfu27clzX6RWl4fgNF3GOyG9zmIV/nexHKvjeu6ylmYiSq6qUjrO03PWvUPWq
gTYxPs/wmIyqZBD9dc0d0dUrIsG2pwCIX6I/Yl/tiqc1/ZwuOIsm8sGZFJfut2Oc
PdJB0Ypx+VIsgC2xaC3fvlxo/eClO9cxhJRVR9rlttWotfLu6YzBfxooS9Jfp0Ik
LTHv6yzC0ijldo4ba1/MUfCuJIba6MHpT230oXg72H8MVAx6tv0HBTBNeGAbn1Xk
N2h/7k+eRa9wrIFPVJ6olXCkoj+fnkVZGykpZlKRGWImpUlzVG+uk4f97OauuCsX
P4nMmNTm01vwQS5omWNmWVSwPi8I3QB0Rc0Uxdqo0/wNzq0U+V+B9Xaiavrj5cQN
6N3M4CLeYR7rO5PH16+/MUmeo4r0Y7tGD8tU1BRpUA2UzDxcYQZJS+iFWgzCZ2gr
GUoOSss+tzxkK2CBCBKbidhJzDDtgexQYZM78qAlEDJr8r0vmFJGIyjzTVcCuaFh
EnOcvzOltO1qsb7yjkmbhCha2hm+i9jaY3wgFWLJJ2/daSy0t9+jejYAShqVDYzV
EEkLAvJkSNFYkuL8NOA9+SEWJa/VzhykDOgJqsOwhvpKcemFU22U+ChFDp4NA4Ez
95mKqyspVVcPdSD6kkbMS6+95Mnh53EiK8WoGKoivT4qgpZRDQDVOhWURYJxMnKU
EWzakodhzuRvIS+znKf2uswcNmSnQN3KsyM3kxWqwgNV6DfviI9k1Z+Cq+5XGh2E
fr+N5+lCkMozE+zSU+vWpyctHS5siVNCiybvNP/EwTPqNXH/tlmoTpvJRkOWqxw2
cMByoAeul+4ASAUB2jiuQS8Om2CaCV+ZFYK+lUysqog1dQ+rxViqV0ofQW4ix8PY
XSOlqDpMIMBP5bm+d/+DbMFYKmJkFz65tvqsEvsvNgecpxq/W9DqT3zOdjWTYPdl
9lb44+yhqSzXHamLzfpcKeKUSl1HUsKuvRwhSRNqOV+MpZUqls1oMMtOHVD5QeQf
dMFgC1IOSe9BE7GOmivqAoTSh5S+42kINhXIHiwSiSw73LCHfUWnxwULBUxVMULO
ksSXE+8yjUzA208vOMo5+V0IDIgqFsrhKX0RSCZnf8i1RbRv0817E9o3Ke3Axfw/
GZUy3K31yrkTyrQd2LcXPlvWmICIBczkzuSkwIQ9WS7eOltS6jD+rr1ekd5kBy7E
GXGhIbgAE6Iec7hiHS8/d/YqDDNscDVtvE0+tDNaKKcDCng6syxdTQXKHyE8bGeS
ETdjkxdriSH8AbRkADhVKZv9xnDi7Ahf3iv0NTSOBUVXVyEjbiDAa+67BBWPrjqx
MEw8jlAtaWJRARW5GUcBqiy1CeXum7gghANgbyGsAm0fp4R7j3ilcRYl+rQbKWD+
W6DBZYB/KBkq+LXECHoJTfzL6Ijze6T9u7IxiiMLmM4ouLe6uiSU8kKUTsgIYBj+
GvGZg8NC+HXvPb3XKODY5y2cs8XLCyCYa7XrPUoRGZAOfvCKZOYgVadLjfIZKL81
sVf5/ByNEV0TTR/rowOJjPxhGcDJUILf7G9pqi99fVEjFVcXQEg4aa1ahmwdb3F6
zOkRnjlYjRVf6shA2ErjkVFn4ZIa+YmWjyjkZvvvHUAh5MJWfjWZTMcaef1RV1IY
muA6tW7p8GMq+IOvrYqz/FywNMhcPhZDmaPklRsRymdlnvgUIBBZWObhH8BGHUnt
Ua6HGVqns/kJASj1ev3hoW5NxuOPPkltEy10w0zQ3K5M3yUS0pqqXL9mw+KhCcqg
a/9unX84vUUhYFCMoyyf1h1D1+afRAh3A9+/l7dcI3KetZA+8wktemYZ1tUgUNsk
HeHL6m/ZkY+oX0QUgGzPwCEO+JNVqGp8XgPCI6Iff+zRT9wRP/VZiKw8xYPFaMff
LAcXKFxH3qDoleQu3SMOOCeYMWSFtJO0TlbKq8Rtx8/jIDC447oZV/Ctbwo1cVaW
lbTV545Gqp32328JZrKVqt9rY3W3gHqtZagMwvxj4LWtRmTz7JGWqTo0wwyhgrtx
J+hqNRaZc6RNQmnnHIEBDiZNBDQuLRhmHuTL/RCrDc+YBzHNpK3Yddg0NOnamxn9
EE418qhm5H/iMsYPWcGxWyDLQ4iEHfwWHeEK5zTMmCvqieFYiGjuBnTH+Mk/mwWm
FokGD25p6zyEAg06foeXymoBOWkxHgbxgslLGGLJyTYY4wkCiDSulLY0/IF2P2qb
12q4MkKsgnsWTXTs19q2juvUZrjneAyZx/2juUsCg9d9EdfMP4YU2Ly7W9gZCKXz
z4zrwn9JCA3Eqy83egUENP+seohdzXa9Btk5yo+WWO+ieQ8ImmuHmzOnf5MrXd7G
Emx+QsaA2zQvmyi/AIfjgPagmu4C8EZFzBsZAzVWQnLCm+jEb+bHGg5Mv0nHbPwW
r37mrV5Q9qc8tMgIApneJNev5uk8H0eBPQQPr4tfnyDKVtZUtuNuSmb/S1da29FQ
mwVwCOVSmHdJscDFb8uLsiC6aISNdSvnuwzRfavoePGPDr0GL8vi4rQ0K/N97Uuh
gNLiPqmDJwJWhrGhnqI2VaW67qFE10BAxybbYSd3dyGEeVczxo1vn4jLkBiaR9gc
iR0xGBJ5czmIAWataJwI8GMC3TYPKNgGGm+1Rd/EowiMF+ulaWO6qxZT6RaioaaM
qHaMDZyw1olLD1Xjrcug9P6EjETbaTUOmTZ4tEzukbQNZPhrc5ENk8EZsGA3LEQm
YgKG9LlKDsR9gB9ncnwxT2Y5k4+0hg7unJc6jLF5Q88znY+KRnNL3J+kD+aMOp3X
rLGlIirhfjosvkmFJTXUb4E6m4SejqbpKOoZzxDClMlDWuRbb+2JHhZoqG+vOtF1
LfV7kvcNrt82f39jdg+Uc7z8OenNIgbD/DYmZ5cC/GdwCAV3I8dUckXFmJWqt4eU
Qe9VZ2cAtxUr42Z8roN097aqMTBt3e1Zw6dovYevWgSrxMmCL4STUz5HHzBngJb0
R9JeMLBKXMzuE8hQJOutYBdb1d64QUAGRWNjpD/kAgvjCs5OAIM0gRwX+aYj9T39
vOys06QY+po0sJOs5p5xloFENw6BUUQC4LF6W22YlmUs03zJsKPNkihPrw4hy18i
AZ5gjUUjecI4iVqI/07+VNRODgCwepASOSJJyNn/HbKffK2VPBGrC7Qf7KqFJv+R
rVfXoYIcBK0b6UvqtCnEOW0GJmW5Tq7U2t88WJLkOwRgik9EWLN1JEWq3bqWZ67W
BMHFB/AskuqkLlbcnhd6NUGHMhBy50+aMZ3ObWE6lHsJCjpVHNVCpSYvZ8Lo61v6
DHXdUliDjsZAg0wrHftgaOMnPHv8JZsg5m8JGaTiCW8+JOBM0AV47/k8RL0PPZ5o
kJTrpU0uSIC03EOIV5xFqAVKY2zprXCSB4PPeNXGWfErLhQtFIM3OakoBBzGG8OQ
xHEg7hNZTBMSms4Fhz8L6oaQigTSwFF+g6bYJZm1GEhiFcXxUeWsg/11KJZAoD6l
LE87AO93UjG1mQJWuQo6hfQ7Vzn/sxUpeIIBSe1sN8IoGDQj9UmB+v42ljIiayk6
IeaGsP2eEETuUF/h6v0M1//8vsOTZgfupNxdKED2CbwOA7UYoeLp73WZd0JsK9Oe
Ci9Jih2B8czLt3fNGvBqCMvnxzAFGEU/Ny5jnrOLFE1o2FYxP/eHNinEWHS0mcAG
e5YagCRdNwpXq3qUT9HML6tuEGfsuYhIN+do+MGA/TmM+lSV6LSa7eD2KJ8CSCVD
WVnSgl+Wy0OVHpyOIgfYEolGJCI8RFyCR5mqC25NVyzYMcY58ihtxy2sJoxdBH16
l1Vd/B1vEuKOSNimCRXyqQ6Cca8ajc9yFL1duVn4Y39c78mTsIi6Pu+tLwBVLtnN
B7AhZq30L5hS7bgSEBm0FIAh3lqFMQI+BmLYA8ugvwr6FjxEWZlse56UzS8YfS9i
vccVFWPTJlFRqv80ERaFxQchn3vLyFC/Kw5futoq3bgVtF/gPho4HcCoCvk64ey1
5L5bDsQrH/FJsUKA4nlNe7opSyImXHu7DwnkZLjE5aYZ/YR/s+RW7fkUus9jJ2zb
MyoEia18Gm368aBClkdratzUZyVglBZL1voJn2do/NzayUJmiucZvKSHxrYkAx2U
RKpk/MdnAfAzk1723w07Ta4lc0cl/lOUc3V8krOfweUDaky9HmHCpBvVtvvFUNvz
WmQ1W4dqEquWcXlXthVwh8jio4+Gq0zw4PvuQkECAb5UoRdZ+obT5upBSFn3nhvI
TL9EUzUXiANYkbxGM3RoWDqhe3LPlyde73rNXPQB7vc9aCB6oKpVMqHU7bPH5nhY
l+flnjBhpQ2cljsHLUHgXBBaJFGhxkwPmFJ+jRByDobYZFgHIbTLZ21Y6K5Vfb6S
/gCfkXdU/DaL0mGFeg3hbYY4Vyc5qq+0v2vqPoQK01kDwmTOgtlj+jGSR1xhLiEC
cxqcYa65WkGdKbDLFxP7sEsd0AlaFGTAsuxTGjpDTT1HavjuDik7tv5i1/Ih+pnD
YKVNxAvxGxmr3oErqGs+IoIeKDSLSSxSiyGCllsuiixDyxlKJ25FVLqcKzYtEGs3
xhIWddNuAhWl4o275geebG0AMNQp8EM8uF2xTuOhmIz3T7TS6yafRCN1K/F9hLxN
7Zc9LVlTo0yfO7wAy04C3fjdVhxoQk5doZ4a3QLe4EBux44x/bSaFi34Ub0UyTM0
NxrxaedL4zEkVfUVZEUoEH9Vn3dEeduDVhuDQ8TQNYXTMJBQGFtCWVB51BKOMuU8
/t93MT/EXeTa7O8/Udp+rtFpENtIRNKR/m3Zjvt2Rx0Cr7NScaRZcnuEOObI6T64
VlSB1wf8OhTgHefnK/LJ3KGFqRhLGlMMksD4Yw+CMvnfboy71DL7wCaKxc9HXuvD
Vn+MgQDsQNPZNLFO1xgyrHIpYLipEWK7HfLyQihvRLHJi5D4DdG+MDYTMeMUj6s8
c/NJfa5HhqvQp+hdSpSXFhbl0upk18APDb3KSj2/r99i3OazCNtOYxngS+q7nkfG
txKyswgbUQOGq8K11La7C8x7dxu99PezLPy5VbzAeGBZh6lYVOv/N7RmEmmKepfy
xBgXDSkp6S8QohKhu8ePM8C2lIz1wBKx9nSFK/c27UT1oVWEu8tZeXL+P6IakbUS
VjtHxfjAXS/zECxBjiV20BaIJfnlm0S1tOJnIP2z3614sLLgDXEebP7tttu5pShu
anZPqLlLSHY8o5CTHY1ItNtSPWOOZnB5ZEP1LSqvn+rh1+bK4+tJMvMXzEXM3ZvH
ekYzSBh0VjHwlFFb48MkTbABxUPZQG6TNvustKoNgdt0SFGt+cF2Qb3x6CVWQD5N
D2tblvzikJL5pCHeJIZMYr5B/gr/DSpph274MuNU5Wa6yUBWzBOwclOmRsXQ8DbE
sFS7eDNKi5JqPywuAN99PRqR27krlRTyf7VTyXcs+A6gNEZqIvrcebQFVKKgjYKk
VZYn4QHKeOrnzlGeYB5XsiMZPPVRs/cAnQ4Zy1biiLBkYKpTD7WW2k54IKUaWXCR
ysd+3iB1MQUBiwjF+Wilu8XaDEmO/aC+hycTIYKrSvPjfUR5q6smu/YmkjsbSMi9
aBsqSDyYhPm1Hsm9oFi4iMospAyNs8Uskd87cLg6S7m0qHHoV/rvy1xyIo5PbBC3
bKIea2GYUVCg3KIrgkbm1GRtah6BFRptS4Sywr0T/sPwOIO6Abu66gA81zlPgQXU
wOdigDDwghtN61Ss2jMeQCNK5FBe2IoWc/SomNp1wstvEptzi8ekkfQ6G2Ksl1cq
xlre2q+d1+sZoYYgL3F39srhQKmkZ84qUSMAFhP5I0Z5FH/TqyGnTQK45032/UQ0
kCYUc18C8o7Z9Y0ScYPhxV+VtprrKPlDR6nxyRK71pD4V8wGqPbpRZ7gtvVLHBhO
FOhq8D4m0VRhOklQ1c2oI3evtnVmnNrIjgxD48rXuowRnJ0blILCl6dJPRs0SVru
mT+PrBIVGeIIcOHiIS4qHNT1aG4mabGZWqW0grQgH2sfC2DX9edCIE/EQnKLbrCT
VyVggcCSJ3IRjHpTizlDg3MCZCXknhBoD7QSO1N4aSvgxgkU+CnS4VRMmrD5yzm3
eBR8lXS4ELEGBQkYCySpc6xrDVZzzcQcld6NAJNeQ6syq1HsyWN7kq5iiaCvxmrk
qAWGx/NoXlc41TaCNBjpCWxLbMLmOTrZRxLqIshXRxK1x0bT18aBXXhw1ygshehV
6720tgtNi9JoRVd9XXnGBXN2tikEyGInFa48OcdUWwOPKJwwLJSvQzXEz/uqZlds
pwx6O0aRvKQVmZ83vw89OgLa0xzmLMYbHm2+dv7Zc7jkqGlDF2VgGlp99pz4gD0g
x3ZQb+SV2+fpKSOfG3gSsRVDkrT4nIB2EkJ1D6i6YFknVlKqKP/4BrPXuilOdDSm
uoI0a7KBWkBbmkseKSKDgJ3A8jyhja4f0NxxE/dmK0T3vMgdH4kGg0An8ygFsa3I
0Z/RtnhaeD8Z65cPu43S85p/fzaFR4wlw5WjakPh49PJjp2yGDQQrvXLmIZEfuC/
7dwYAzRJsNtKRByKqqT2iu2aNYBXsb+M9n1zhsivAfMnAqPsmyrtx3zVX30T7yMi
zOwybTz7QUblItM8LJtLXNgkRFblgcufH7R+zf02YJ+e1nQGl7uFZGlAi6jsJ0ob
NIO8ynL9PtRUgk9feAyHKkK5TSt/fIHp5uhPJtdKs7/B0ydOzXIDsDG47TqVAhg6
K0ycktdNEIjeAt1dxPD+OOu4/sXDN4dVTB1FZiaNcbtK3fWn0mXWEwPSfSI6gC+U
jn/D56vURcq7Gv3kKZgPuMzMAa03gA2DwVSA7J/L/bFqIF1XqqD6eKHdrpv6irqr
IwLBPYwuR8q1olJ4bwrdjutwE8KO9lIHE68cE9K22kr0mEGq9Jlu1A34AXxEYftR
9EHV5oZhMb9XpbkB+S8NrT0k912J47mD+/iRbsX1mJF/UTrOZKNYTQLcchvAl7xK
QsIIwoMNt8O3bQvwDGzoLXC9Nz/U3Jzgg9Kj8xFRA6Zk8JAU2wQh3uesAZoKYhIp
Kl41jP1MRlhi9cOBHmU/tXRGkCrFeU2iHk9HYDRQaUJkA9uCujULaz6dv6iz2ECZ
oLXreEFJFGg4DZrFZec9LZ5azQcJLvXpX1N1CslTcDLZB00wdRmo340N5AU3QZK9
SNdtVlf3wgurFMfwFPUnvVfReAbdFd94kIJTqtFpJWI5eGlFPeHUZCFFmjaoWLMh
ks8XJCT2KuLedS5yaz1Bw9l566nFrw4j5Va7DwcQYeZbuwEEvycX+McFR8azu7E4
yL7mHLNBww96uDp+5/j16WzGRhtbB98UzqzffdJv31HvWitatgsANyEjtGyAObwJ
pi/L9YiF4+6U34f6aHvlV2D7AoUn5O1CPMsj17M1LnQnkSaGWljPf+hQWFPjpgNn
WVBNfUeD4nyphzyYFW0ZoxZS0E+EBUZ/wdINaAI4aE0VFax2yDEgedPyjKGdUDgm
ppflJq5tsYVzs5ga6VXHHQIBhuwBMM6rls9HtjCEG7zkfsHAV7N5pxZVt8IkT3eN
FPdTuqfHSbGJITeKBuLwrKm5Z8udS1OzM/C4bSW5KxhcJHD6bEkir5l2VWvjgmg0
D+KcQSTzZlPOTkVzTHKIgklP9AkG3eh/m/hhkZ/Ry0v4dw7RyhmWCqiBNgYnBjUf
d13J9RQoX70SlBRUb+m0Ht25kzuWQENXjBKoCn3tM30s6h75TRAK3LNvoXjG6XIe
/HMEpuAOluysH960zVJFr8U3UYN2pmihiYyQ48zfP3sYeBpWMVmYChRQgUSbH4JY
Svx8XSFgeN5/bMx83k0hlDKrACnmSEPPy2TnzOOcvwol11d2bsR+MpaAYpYZaXiy
b9dnd38kmXkd6XyIoH5oVnjrdbwCK0AVhxGjZvFe+b55EuYqPEALOfpwvKDi7ot0
RWmqQa1bHvpz6rKqkb1kbC0um3bnWIEOuhcMzc7+V9rCOvGnJkuFdxlX0U8SD13o
EwFTgi5N1WqqrPLL7tKxe/UNfDXAByW7wpE5aNstKzu9PRkG7hdxI4ByKEtJ40v9
72Av15GCZnn68J9ASo3kU+cCXi/hganJpxJ1+9KGTxCSa+OSQEGLmQxHFGRY1/xc
u82ZHqOeK6SlUrvhq2v59Te722JQcBppU2w/cLPF60xgbgO8tPWOt7eFkjMPtWdo
unRpXLdI4d539BtExUnCRJaTVaKyJ1hSeluuar7Src4Yk/wT6vkbUUsiUOqlzYhz
K7iZKQFnO1mbpEyFBY6ypBzvkfZfDQ30axugbnIMa1+3RaRZxnCgJCskhg4UHaZB
YKz7gRH0elkTOCZBoWC0eiXnkRQFLiSra0atNfEZ6LM0Xh3OGkhXuH5zKu2YNYUm
tiSQanHCfP/sWS9oZiTmMB+qkeC90FezVnsn4WM0I8H4nUXydTsvLcI596aX4YnM
dvk3Opv41mpSp1rjjqsZazeDyI1eSnsAkxox9cmbr1CrW2ymbV0RigBk2//tzmfH
yKE5P7Bja65UUOv94B0+FTPaEhdc4T144zW6A5v1Kxe0tKvYCmBQh/fJt7F80fy8
yX1ZpqQwgZy4Yn7VEpxuxpz/muCDa+h4xZ8ccAoVwN6p/vC/7cb4gIIuD9un2DNY
fSYuc2ip5Ps/b6SjrO3TBzk5N/ipsgMbQEHcgzm3K3fWR/5j/9i8wehtuSicrQdx
MDn15aO9m4IvTNtLetEKB8IzNm+Y6zcD3Q7Se7wnzLQHQ4dn7v/uJRXqrbLZeYgu
EhSvvKl/PKbl+Cnyv7xEwMZsVBx+OYgVRgrAA30imcSvGFgcgy5UiMWNdvkr9bLw
+ssejXHAb9KApCl+wRi88zV/SwnH9u3SGc2aPiHBYAzS2qdd/2hSqlKoEmNTbFSY
53MqYET7D8hyJZbvYLNDu0LjQLkndn3ceIeVHEv4gnqbmgrzHmEygM9DH3tqm9Bp
Gfh/ZtHd0/xkjLjxlKjmyFFqxpaxo9t4siItKzd2x2plJ9K+ywqqaBu0wkMj4frJ
yayJf/sv1LVB0ZqrUUYz0thuSbjA505ssO9EVJi47BQ8yGVb7oYAq1HRw+dWHBVo
zUWReFU9IiVtwsPN+95HoRafqAwMePPJ7/EsFir/4u0v3EtGbh9MV6Mvup35hh/u
KKncFS7LD8JZn2ahNISO5Y57a+6D7tRdkH8HwV3xN2Ou8R/GnB8ntrcn+8oL5dqM
sMCCkIdjBVnHd/BKs8XNJEeZ/1o9n7oaFhjKKQwfL0Ef6lj7CTiIlbkQYPiG5Aau
/66F+a2Kn/70N4luhCEMGNnju2x8ndIYVXvdvZvGwNY756a/AohddJ63JMmb+xl8
3r0C4CyozqWBc81N5IcQEKrNuZvCDgFODeaB+XcLjT4W6+KiBf6wum45IsY2nLU5
HjVQ7UP0rQztD/y/f13Zfh/8iROAOJWA6syDQjKa54hM5zp3ugxDobWOlSOizP3Q
OlEtVd6UTALg/LVcCkJ1aKpaFvDPhs1hpAFxDnSVgrXxpwazTtW1hmxSqRnQ87ts
rcTpr9OfRHZYtlImMjncC9oueeLqv2hUkbnwMQKG12KIcaz/UCSbyjmLTACHbX0h
SXFJ7Y5gTjK1AMkTZTuaDS9aXbNgc8DiWmL8IMOJTeSvAb35NBLQKMIOfW1HXKGv
hV2FuTxS2zsDhshyyejtdytgIRmMteGa7CKA9UFbpXtVOPtdKLSA5XBPOuGiqoAX
MLy/8BRpemw2qmwfcN41JrPozJVD1VQbO4jMvdYIiipkcuycMzbmt8kn2UdNNN28
6yVJInIDqhwZQDOZSv9ttGtEzmszTK0gcoqWEEdwOQb9ArSzCkDy7wtaXMfTgubM
nB30hBGL5dojFde/LgxnZPMKcnbqAiVuhL9XgAAEfqHNkd/FOUSrHtzlHFGh//EZ
UMAp9gYdjw8CwutR2dYL4PIZ7cP+cT0R8Yeu6RzQ1v3N5nJduIXLWvxGS2ZbHOHA
RVIRmxcWxZamsc3A/9efEiNir52AgAUbo8znzYiaPjNewJ7kO9kv7Xs7ZqapVuHC
pTldf30BEnQa9xwdr4VUfo4O1qqIhbxkDXNWri5KfPmNCsO1SbWOVQWo9qHzRLYg
i6j6ak5MJqEma6Xh1OJdAsYAOACn7VZ6z7cBJjACysEquYyErLdNE9lpCVvFzDoz
FfMP9Mkl2UZkqIkaB+HXxh/eGGt5p6S6EwCqym0TH0Grc7JKoXKmgqqca8cP7vSq
uBBjbEmcjV5UrqU7VG8oifSmZmFBhV6mJ8c3QfIHB8E+Qq/4b6+tAFgYWg+uCzG3
Lv205jRIp3A7pjw5ebSjEUFSTp3cr9peI6TtBQHkBB3CXyZ5xv/UgXvdolXHKERp
4cj8e1UW8Y3Wp5ALe7GVJtk7FTck9GqIL93CdVgL3LWCfZClMSqlORD29qoHKzoD
XjHyt0GALtOKVmRTBxaWSZFyhpBu1Bhf59Ip2ryk1pBC4YzoL871Rvzr21VLsR6y
BB2JF+7k1jZeRrtsj1w0yTGbaY8LkFUdMFtUmv6NSMTlGl4Xo0d3hX3T6PjIT/qv
2jKSCSB3F4HtO2k/Dz1pu/UgkJIFpiRp0hE/rTFkLhW+W0yAJBBFaAKPHpiwW/HJ
covsHh4vuRhg4y9znHVRHYLPV82x41CPPLlfOp7YdCRQJ52T0mzlE6LJBGeXLPCk
AjURq6WWC3TmR9ri+WqHPYmA8AalFCf7Zr/Gp0RBkXE0zYdvTdzD5sUKLFRW4kSy
BO1cN+2JcY9cjLKwIsmdUQiZyeyQdd/sWB3psdQOdLZyghpFKr4ZJlxptSIbG/+s
YuyWajEyj1ak9323SM9cgB1MpstiQWIKmesP375cj8N0C01H3u5KlZXU9nobzdeT
jL7YZNulg3Py5/9UHtsSURB1QECIhyrt120dC/PtdrS2D6D7f5N1L6QCUEHX1oTc
8LaR12xmZOjKQ7P3LpJEfDw9UJd36bXQHwG5E3SQKfRX6SfMpE2XfGxDvAhaK4rN
5XsrqC+naNcNOhUrFt8AzYlu3HQ0UQPXIv30emoIwHz9wX+5T2pnOPv/7Xj9Y0WV
j9r+kNS1P8wDSUhwl2atBsr41wE4ZUYFzekMwgtrkdSny5387TLHU78OIxqdtOvM
1qOdle3ui3u995K3/ve/hNhgIcd0ekLTb2tPsGTpp8r+q0R9JI9RmFBof3otQAVs
9+SnVlDMaJjrfRG8COc8QXnWQKyTrEunDMAwrVgirVeEZhVFMFam7PoDKTKEum9v
r6reHb+zZN87Ntb+AQ4LQ3xwBWrZSMpzKYPWX7Jjgt0qTW984NSDWgBr3uFbanUK
f5hdXyOvD+QgWJ2g1GbBA8YKKzaZZWptVVpFUnNnVE+N/M3zpUk6Jr5tYLcZrUO3
uGCOhtx/yS2txG073Elmn9Nu1HCAi/NCvgzn1DlynRW5i6icJlLjiKdIa86fuHBP
14JJSnRlwGnLO6Z17+qaIpW5kjdWEa5Ry7ghr/fIO8uVgCmL5W1Ki+iXXH0g8ZH0
eBBPhXE1nR8EFAHwUa5t8wNF36ndUmNEu0bU4nd23ReDf0PQrPet99/2SmojhITo
n7/e2Ajunw6Dx7DUu5EkC7Du9cT5QsKHF/kqm/51ra2aO2/e7NBtbbMgKR0bIMcW
p358bo4zARiMSMM4ewxVZQFD0B3Hk8onD1bexpChyo64alIfWOOvpfBhAJ+ngOpr
1QN8d3RMOtfH0QbNtQhQ5RRGOTO1CaNhMqKiivW2t2qBaxl1BbszlKNHn1RqKEsx
tZfEl1CaeXmCmgKWGGYP7Ow/EBICibUvUL5r6uU678O0wKtES5QDgN4JFco9KojW
uxSgM/doKm4L9biETYmU0S9A/EhAUVZLsA6e0ouqPdNXQ3BuWipC0LLQOy7NaFTJ
e7r9jW2bRLhOZr0+XTcKGA8tCm6JkLLSYu6LaFJXqnVlr2YV8J7YfitfhLcO+htT
do58gD5gDL2F8fbn8pXGQSbGDX28MZXhDTUQJhbQQRBaDTaB0HUNAWh5o9DbjF5G
5XsD8wcu84RQCvej0axP/Z69vu3JtvzWEFO1Xzn2ROcBlC10yBlwX+HjXiGVBUS/
grWxon6G7pSvswxJYjDa5/Sz5SanQ1msytxZSteU2kRxt5oi4Rx34vKtyME9gd3g
1JPuiPjPr1oT+ZA0yqv8jkYKoGnL5G7uv9KT7qTwUjgx/LWyowf8qGzjIkROdlS8
An0e+Z70TjKc0YpgAxcvA00kaDtu/dOTY8tdVR1vt0jEHd30YdII1SG9xuzZObhT
eIconUK4gWTeWLqbo0WCEul4fpey0LTH0OY5kldqMXtbyGoaY6ugzEjaAdkoYCaj
eBkuqMXCuQgzpppDrNHs26L3vrEk2aLBtk9Fosadeq4PNDAwfg8TbCwffRTUakmO
DAYOYgFcpgAtdfRR/eKSlag1lYvuI+bTeiOSz6rySbY9CINvf6GEgTcySKCBfHzu
GASgAwSRg8nXwvPbxHKfPs9TyAv3uz3yDYwgB3oFK/s0jemqJ7cxCExDZXL9wxkF
SZGp+RkDzYoVGCKE9SjIprh/KTTofhOSLKzhVTKb5EG5NJRX3/Y1aODK78kb8DrN
7lZ5AK3Dnb7gy/piPmuUgvRDSunbaUiLEHhVEsmnes4xAWWoS5yfGex7Vttxj3iZ
KiUljqo6I6uyVYHeXl+dlhYxQQXseWNge4wgtiS2uIU6DSlA1vwCeU7GDDbiaSeP
8ceE4CF7pWslU/HezHMYTgqp3oHE2MIJKghhne4m7dhX/vJCWhEtmx6+LOPr3HEf
SAAxzAAZN9eis4CA8qWCw0mzB/b7VI/JO3nduXJjM0E2l2mpeKHKv4NI0eT593MQ
pYkdiv6F8eTPuiyVSC2ug4NEZqpPC6jA3zY8sTsOPl8T8nTytbXyGsilJK90YCeG
jZqQ1RA5ykSOqScGoOsIrnLhmKiNlgL7/Dw/Klw/KFM8qrqGsOoDICFBxT3FkvqJ
b9IqRCikZmNt0kOJxm7YZTVRx2TuaxzV8ldaOaSr7q81SkYe39CUQO4LTaOL4yCn
zKf9qvlzttk5o+bhgPjaVa3JWbV5JwZcqzy8pbMyumIzrgyMd0vAIL6rxmPlN7bG
aQaHaI9Z3qtcN3J7KnCyhVmMtqWuKVUBLxygGCDPd2GXHGNvQVypyOA2bmO8HUH6
Xcp8yZibHcS7hk7tbmsHexYyiQ75BTYOxDFioAjbfDgS17s0waxWcanqWDknZzGt
OVg22kWxKzDBB/+WLFs5MkkRFYmhmupPCWuCeHsbJP9T9dtq2EtutHpLF0PwtY9O
fU6u1kWRcFQ0auivnFcaZWjKSDVo6uV65607IPbpbwzf5QNSQi8coQBA7EaLcJJa
MhbO0DrkgVGtG6PfGYvZSW0ixKMJDK8y+0m6fxmvq+7L1pK2v/MYeU13HsUdTflX
IqDGaTmYla2bRc1S1WM9yrn5Hi5LQjc7I29pRgdXA65M4XBHL8Bij3RB7XQ5Vjm4
WQa1/0zfp7GqG1Te9yNb/GbYdj7laqA9ftlCyZl8gGAC0g4uxEOzDuggJj1ni5Wf
RFynm+Eqe9Mrb4rJ2IUuR8xcfr1WQcUD91ptChwyd3OmDc9dVkRSbJ5Atf/h3p9Z
sVxU9/5nV46PhEDmlcNelidI1zT6jhTFcGkMX2MzPbIDazvmEZASyXN099O8QooC
U7/aF5Tp3Au59V7Xx133112lA4WXa+d+yzleqwNZBAEh9an6ZoSMC5QALLzqOTlP
+bEyfSjCY1unpuVoFsnLkhle6AUt20/jaNBBrpBCfONWD382JYHmbiUUMdknLHVM
xEVAuVRpSDy3qsvICBK1PTQTmLBbHfAanHfrcJTzW2x2+/uxusXfzHMVdiUOw4c+
fBJX+mZ4GiSYvXYaBggArfdykcl9Tr/ijzPNL81NiHGPwXzhpcVPLpgt59QEfm4O
mY7H0sfbimjdo2oEVAWZZkKWIDpZ7+CTfzpXMa47SSLvPPFBLopQCCQBgi+CbbRD
jgVMDUvk786sXAHLZJCq/87m4Q1pZ6AURsBwheXdutK+4aGUE/zG1Nvh0TZht57U
u9f0gEitY6lCtKzOoDb2SxTG/haSkjjCIr0l3pmwsLvwdab5rmu4Fr9NctBx2ole
j4tMGuLERNQg/3EHRz8yCHFaLlN8w6+HBTEOO8co/csHmLUATnPPwv45bfhMdZVm
SWYsnCYZqgPHQKl/A5lr3lnkcAwhFbqtQfBG44rzf5C8XnYvdlqrd6AtuqJgQY32
Vkmd+HXx6xMUtAg6nbZacnbuE3n6NQ3y2AZGaivcyCPxb6yv7QWLhCqwUGHXzlEs
awyzOAoIzOXOcmnXVvY8OW9sd2Y7y5FexO/G9AXifdjqxVcYkcXIxb3zqDX9fWSY
t0lMQYqd2pcxBSR4lOG90QCzZmd19PFk1000tzHfV4G1wig6Ek0/WQdzb2k1pOa5
686cprgznNwXdlxwleoTwc1b2m+tFzo7hKIQuSrlda3q210/xJ+g/Q4uCMec9AEv
Y4ydIhRCKk1BBwFO8eUN9a3/2jSLbrqylvJ6OucKpXt4qbJTExG0Jwp834lp01wL
TMQmy9wgl79kbc8i9GPKS7GVLvlPaT5YxX7pFs0vOn+SFelO2ijgauHxxm+HIZi0
Qk1d5xPCLNTiooHTXqIWbwj7X8WdIqPHt39GJy+xK5/UjpUDtz4U+k6iO6Yuryxm
+GUOxct4gUNiBJgHFoE2BfwHVDYtGBvvKy9zhip3z3a/X2HUUvbnpxr0OXIv+Zbi
RH25a04AhnP9ZWmLOLs71wAAHgDjJvf5CGgw3Tqfkx5tXOcIbWOiXUhvE7DVXiTM
zsZnoLMvstzZJTInqZC4eChXP0ZUb14NQWxew8e0ABGpeITspgt8wsot8ELOcvzQ
pUrNimpgpZFO7155ad70Y4zwR5W5eBorg422okNNO5ZLB77g8Bx/SMP7JJPyJeyT
qaz4I3EkerjYlvQHIrhf809NNWm9WbycQhi+Rv5wsdN3Tod0eBLJyFWWtK2/W1hb
VVipR+7qk0/7hkxEWkUQwsUXPXD3dbRl2srBNuDJFomJ1NteloBiX99btLuKjKSE
nJIqOCEYncBtV96PWxHirS8Y37CKaSTpaH7PGp8sSFjq6lTVsGNZI4JgISUHsnie
dS9L4ujXnE//NuKIEywPcSDgKaDyIOKPHiDrgZ9aEkLzN1/R6ByLITj+MrEe2Fmt
R/uzidB5lLe1st8GQf2q/59XY+xBKz7FyWrAQmXQnHs4miH5sZy19h3wKWR9y/LR
ndoG9hLy9oCrkG9tG8KWS60PO1geCNWF3UM9wPtx3mlhoUwkJffaf+4uO3mEUfmX
WAQM52ckcVoV1jwwo/jWjag93wAwKXPavXaLzA3pvWFlHWd2GTLMsm+CPyBt6G2v
JPKp2CYAq8B2RYosBSL2T6W8CWo9L1gmgk8Kkv94JJU8exRV1obysoGfdBF/2IXL
n1559zGAahrZeo53LfEAvdjdsMtwAHv5dDJ/mwCEhaMAdrWHhBtFQPacjxp0tUO5
iNxH1khtrDs5eMeWfxqANnJll/su5+B0ZvYZvUpGuXsefmdv82hF8WXzYzhzMzgG
Ryk67NzdOwSKqu/mwPW0haEm425B7WKqZGcEnk08ga6zxpqx8b3w9ZD2nJexgjA2
4KFgg60TNsQOpglFmqPvqlhlBZkj7g4vI9/0riJnUxHHvvXe9yaWFw32Ch9WIND+
RUNSNOa3UoYHW5Wr+WTYOQo1rJ/dmJhkVmbN2LhknNo48WDiW14J2sjQZB9kzZhS
j4qkjsc93tec0tlgB+pZDFdaI5hDKMXgVrw0RuuxWpCI25IWm4ziOxssFUhEAPWU
J9oW82xe+fF2USQ2o13SKH1Djwd61riOe+e3mMZl56HiiB/oFjqJivXdiMtNYgmG
Qe2N5WDLkoTqX/PM7CaZfw6ubhRYmirdpGOrSuOtdDO80o8v2TDmE8LebD/AG5mL
f3o1XgymrLoI9DvNXkKPq54DrbxU2hg8jFguoAkO1+F5PzC1qffht/vCz6ovDsqp
R4bxK1t0dXVMBVKMcTSsAv6ISwQe0AvSHGZ8xo7hogXrI3YzChPIw70jJLQ9TeYC
WTaWHzihjcEhzKEyTi4GJQ9MUUPlJc/7d9evTYLf7avKI6Vtb8i0U7ob+Lyc6Cw3
1plT6RxYVtpMn6A4lj7E3Hfhm3yMDFH2FSYdifAuN11hU7k27fzYLATjxgeN4Cnl
/WcG6VBduPHtaWQiIWbk/HDbx2Rp1pyAnXeOnOmYRj2iokR/yB8WvQHc0K/CP7Gm
D2k9B+CTJEpOZSIl9KSvxs2UWj/S/cPUN607KHOgTvYtiao/vAKhgLaBNb7N+FG5
50FsVRNTGx4Sy7ObP1sKZo71AC0txNpBuhun0ZKzQaNqyC3JMP1SWzQeaOCgZgwp
TPklXutx2Y0NPcOMbtKbefihaWtsG8O6gKEw6Ly9xvA4hckT+tEx6Tl0d5dp2Fa/
P0C9vdNlRdvb/igP66LJcQIyTFs9bnhAVg6iXONFMUukDk74aXQMuU3gHkuiqyew
I1w1JaTzXvsIOraO71HAFUB9mMk35rjyjdepwcn+P3kNGn+4VkQKfknM30ujTGeu
Mp8+41R8wkDSpCjMKOAZ/RdPdtBtgxOCgVPpRc1fFBQrHmSmG35sJJzegn3eu55p
75Mdl4t8E4wc8NjvO8bym3KM1osK8aKc6VLZ40Z3VGQ5TAuMnVdyzxYN7Ji+gI6R
e1Np79xl6y+DjN2cDHDqT0evKDZFDyMNePQ5Hswj+DifJ7JRMVRLiSTw+t/Tw7qO
UPxtcFFOe/exmLaydZj9LGGREFbqjRqDykvQZQ9Gk0o6kr1HRg0ylBaaEshT5Gyf
WcwOSa+mXI1e2EL6l9ggCF+r7vvpG7l0gkwnSMCpLmvbyJsDsDNlwxLTBWsDBDYR
tlxTYjCV+cYvK/dSTZwJWmoqck3ckL/GD561EvcudPXwCGHhrC3AsxOEyDJ+0PE6
ja+mY1yRiUBqQygcPSczNcaLfxeLXrFwnO77U3SdMwrAxpgv0H1JALA2dNI3dYYk
LpOUZudNXdv39L9GybYPEEuYe2csTcPDUxwuTv6MyaIqOup7ScbvqR1k6kb1dSnS
IPgWh5fYqq9t7zZpgxoFKZiyeRscEbZWooDKOjhVlF+yF5uRB5AEap/AfmaE0Eub
txVN1t+CpgWYHoLJq+OHQjD6RuGuzpa+xHbEHVkDA5MrdqeDXA2KRHCY0T8JHjRD
vD/gi+Mv++BD7ZR6c12bdS6yPRmGZapkHl/jJTGrKJYwnT6Y3iZOghsCsdi0Khls
6c9GfNQEfqGF5v4C5VK13cTni8FusRRMXFqCq8OGKKP9KbmhrSNftpPcwn5McP28
SxqdH7e79NgIndV0XsQZaCYZ+l5hduXv0/UnRef0CiWC9c/5cjT+B8p/U5oLdWy0
dRVlnWvVpYHHPasFJ9SbQfVR6KNonO1VhPxTpsXn+Vy9+0zGTJGbeaB/d+uPNBMW
AHPcI+oyXWt0vKFndo9RhKrBQfIzMdhTUDp0/4Z80Id9syrsfWCHfnZq2iU4tpdr
TL71xGSOlgoejPJUIvi7C7S9JMo3GLvK3tfsGwJMu+na/WVq4yGoOuTyfwA1O/Qn
oMlbXoj/AKKe82foU7to+Fl4cSqCgC2OsE60SikSzFbdpPoq4+ZkMrcTNyY+mbL+
wF0YcdgKt8anALMj7OPNrZmp11ltk757NOo/dna8hBZveF5py3wc2I6ueFzEzTL8
u3I6X1Glx7J6MMWXMEqOJ6Zggm8AzGlq7VTp28xpxarz4rKzN2eLZAzaBeTMtJ/y
eJWrGM5iQLXdDYXjzievIXBxF6LKOoXrnwHkyIrX1oQV9XclFrgvz5h6Rr8eSewA
EIy83n2c5RLHJhK9ovItthz5oXOKn3H7XlesiaZ/TYVL/9kEeUWCWQeW9NjK6TrU
4ZpkUe1wyeIsYCDNPJ4FJN+1Vism3GbdZTaiDopKvA1QderVjS57UVzvHcmryU2Z
PsQwskahRCOYLP3tsra1bXhrAroVirzWpsLpig8EV+j5kJNvFzJiEBZRv1cu6bRX
gta8l8TYZaSXJeUyZZAK7OgEmXEn1FW5JsKUGcec66vWZzAYSv3/8hxvzee5B9nf
dKmYg3nuV+n42YO/UJvWYRH2PjHro6iDS3OFYYQSBHA45ljy0hvoPaurmmnXZo69
NOCDzAD5LZ12597tSpP+jzcmD/Sc0w6/SxMn/na/faJdS9b+68lFkgbbs9LWi5du
9sOXVKXZHH7fqLdfAYWeDvt1uQwxQTdtPpP+0XEpwQhkL39K/MbK91rRrHOSGsi1
tqKtphk/EEQQVRGhcwTvyupXIjHkh47RbQgPvygMd3btoI14/o8NSvgZCqgaJLZp
Q5TDFPILwIRIdaIsAOqFdi6LKJcx1za4yNlT1uuTEOI+9dqm/YfdoDbR9ErFRoqN
d9YhdV+gbfMScV4T7WdBUfrwMBAOOdBzQc3cA+U92ZVQbuEEd740N6PCRznTj8qz
mJIqoGKmvKrppvfOdvh7uR27GIx0lhZVc2HKt6D/5d4A/NOEPsLVJ/pBOdZrd0bb
JnR2fCsgALt4nc5bFc2bMQdw08/R2DkVDKa31EWY/eeLSmReNbYMEAS5ax6/X37/
sRZ2sF3tWOx6c1DJ8YmiIznHby9UjK6xQOy48a4I9zs7cY6kXl3DJZls6+5k4IOw
ps1HNrmKjS29UxWrbES3HFSpbSCeAKFKA/J+DwcC30wMPmSwzrcwlC+gGXS9E/Gq
NXe5KUwppj0VAX6qeVqc0Qxd8NhtLQ29RQyYdqhzkMwlSqGeeTqIrnrY7Qn9DW+X
y+Hm25KOI97fdpXY3EhbWJO6MWuM+DpX5apYF/IkPIeBIqxt6bt/obeCU8PdpkNQ
CX6NUWvPgel+HjiTLVFR/XXXJww2R+p3c3Ivs+xIgFuEpjBREg3PaCARs3OcBmO6
clB13YZ2lW7fLFfHrKiCIWjzQ2K2DFDJTsXNkY6IKsOLDYZ5yF8dVthpa5TVKwad
p7VrVYgrDzozRNgy2CXwQBaVvweeaQx4kLaRKjGECOgGM59jUyUb3mEzSC+hW6Ji
MTRyz8oAuWh6Lq2aa+hEPHOz9rIwsj1qyWPT9ka+lriQ98bQsTtk4G9cAg87yx6x
i1YXxd0SMhgknYL/gQWnE4gk//vhYuuXseYYWS/DnU92MYkisapAIe2yd/K+f85r
pfxog00r9OpZK2Q8hlH6yQGRASQYuDsVEV2CUtGwdhhVx9XmEld6edqswzSiU3w3
h49o0kulk8fh5rs/eqjzQopYMpT7eGzPeuVP3NNPaHxfgJhGKHrvPIZHbFlxmW4A
8ouYBoN+1OwPYqKjTNkE2wygX0CAy0QeJxOujOFKBMPdcyMqlitNE2tql57xc5Pf
HoTH14lAHaJUJf4FuWSRDFlY1SgxUPf4HnizYFe+4B9Daj51sWkZNysJpjORd/jk
FdbdCV0CJ/AR67RRYRS7lFDEMfKRPdFcTlNxvGc1mEzNsQ2FGU3jdqmN5Kz//6h8
z9b3y857J3vsRatV5UN3UUaOOclpE9cSink/JZ7/SCiIOedgrgcBBDqfpxXFRntn
2oDtTitbRPlorqbooR1rVw908W2AadbDtt+n1kYTE46EBcZ2liV0iovNEM6rKXse
V6KPmklCMqAgszT0VwfghXr5spjR1fCcm4go57Bx1cmBmM09ZyrK2XbA0aAF43Mi
Zq5hPI8g9Lf8Rzy1N+1tGrFAsGwZAPQ8nWkIa9m1a57o9/RQDZ3cjYAGS6IzDcbs
2SNYf9c1oPEWgooIGBhUv0UaABLAAGTZmW9GN7sCtUfQtUVoDURG4QB+dT4M4VM+
PQ2TILrpFdtfTD9ZavFK9VfuIcfg5fe3/yBWWPQottcW43BWTjAddCFzKPuubDxG
0FK+/8IsDm98NXQN8lvTd+LN2CBHGP3U91c/2mrCOmG8g8XTbRMFbo17AwXFNqvX
LhVvAuKhxue6bplkJRjmTqp+FsqZM3RYNC9YI88nceuEv86R4W7zZ1rRGJiPfMAw
G3OfRxLc5DR3waRpJzDkrVnVo8CQi/JQoU8uAYUDE47cIb8vj1UB5Tde/hS9tSTi
CCCTscQunKokHhYk+SRcWQ/QfrRtyfGT1wdHD1FyyxmSuURI1/gfet4ZXNzMcN72
RgO+9mKU7E4H8cGX+83mhXN5o/WyPQpyWst6ycrDMdNKXocjexRUNz5kdWHxVyhe
5JgW9fYmz25JGt5efNuKo3ugNmsL3zFqb6KCb46OffeHstvZ35K05Owg5zzz8gMy
6YvG0wKHS6+xJoMeVeXBwlHPfUl3iy447aXZiMKQ7dd2S6LLCotuCZSl6bVEmF+7
2gfdqZzAyX34bXUaV2NDoWOSV63I2bS9m9PihlebCScJAymAVANQJHot7SqIVLs0
cP0dw4lMrZsyYuehLTdmJeVjGQZqIi7Pe+GuI0+lBORvyFQ1Z3TKU+vxjl9faXtu
gPwC42EIi4Gz0JNnqkOz/MZ+ISEP3xEnipQDg8LeAOuy3W/a3RHm2zFyK3nTjgui
zkj9+kr/kMHPE+KwLWLjD9juK1m4KWKqTdSQTRmq7Z21uCxHevXtxZDjVQQxKMEw
XhLoHBW0x/RL24k78tKpEN2G0nVy74eRhEtSzTZW6ZAnFU8qhrYkbAe4Ru+K56z8
9jZvfh8kcNOkJtw2vtLHPD2ATiICkl+Rtorhdu1aBCwHipaDV2NNWQjqjkIomDFh
U/y1gcEiaFmBlcdu12dPQuzcrffIiGZsOf7jjlEZ1XMl70vRiWW5jf2tyRNx0flv
aDOwXhiY0ZhNJ7b02V3n/7CYm6325BV0Bd9zt/wJrSEKoN96kwqCWHq2QjgCK5Td
puPY8a2+LNdmIXubibtEUhNG91zZJK/PoRg73XuyxIUHyNyWhdHQ/ywgukRyhJJ3
G0xT5zTMEQlYJRcWZyD5PCVcmf6OpDuzal6uMtOs13QVILB18S0QfATLuTWM3Yf/
qlFFtameTRGV8qlus3AFSKnqaAlNITuD3d4NnRRtaH0hxmI6i1fda1n1L4zQTPsb
mi5bzCteeOqm5b6VEEEe0ID3j/sFindWwCMlFJMPaUMxLNIfTY1eX0YFKmLS3XRN
NF5XxY1fNlFkOkR0F0xT5F7VOW6hbKAMgtP6EzzyP9pKvstvIxbxVsoKLkxfLPe5
K3gqxREf1UEA336kvXmirkJY801SAP36BiTrPhEvdm9JPg8ovVDv0UKMzvYiihIo
QRbVOWBUA+Uvy4kx5vAhWnsEdbQ7MULMqJJwz5CdCwbDVZFgvv8dioVYrhYUlHzS
wv3hqc9dCxOdOZbPdm7tiCNLCH52zWMjSCeOwD/vq45GbZt4q60HcHRDdQVyKvTx
WR9h1iLw2YvgeUcq6mG+GM6YUYdEkgpwO1admalGnXN87lqRDMomZ+8MR23xgBY6
aSi+yPQ18ewAbFAhmLYUPQsx7KHPw72r9vaRYMalZUNVwpbxCxNAn+0CmmuAiW4P
wC1fhJxGiEUyIsxrYg1Rwp0b+2ceCIJZ2QtsHlZ97dSI/PL+96nWriVwxcWgVwnX
y2zv5SUz5Tx2k5CteRf1AIqkTDL8TAtHG47Jz372hPj+zRmIY9hCqGDK3E1GERyp
mQEzeBkKtYpHzsTe6qhQzAETKWfIp8WV+XIGdd7AvfuUxdsAYHtgEH6h9Tw0KSYB
p2ddcz+3gEFTZdgKTI8X0J88cE+c+Funa+DQl9JSUYpmfAsmARdUY5z6eB0e76Gm
v3pwrlxjRdd6j12H08qWXiRpVSrLjGzzysl6zYBy5b7sPOVcsrsE8kd10wZrmRnv
FprsEcAYA6624SGX4Kqt5R2chRMzHzxN663iFYvpeDXt3kexitsYUaXczqoO/iXg
7iYE3YCvIF/H8JdCQSalwwN7baf7z9wDYR8aOFMkR8sO3eH8cnbfDYPLXNr5om0V
MBK0jDh9QRBJrf1p48I3fF8iX09PhvN3uYobVIbXgI4u61iXolZaObSjJb5Nz6Vq
mC3k+rj3d88QLGJJkh/1o6w4RUt1ur/KwY2QmjziCz0Mdm8qu8+4lYERBxi6o4jt
jlhohUCPDy+w0bH80xIT6wmJIGoa+wcSunx4Fei6mUbO/qPkVVJADI3gtzcfTvYr
StvBOLTJTQVHyMRCK42I3GnYkEl5qnSKGsTmq3D5jwnGoZxE6GNuqgf4rhWdzbkd
PWg3AOz7EgV6jeWCOd5m9rRAuWjJ+SPkuc8aAV7WMOaZTY7SIDZN1d2Qvq3AptVa
CJs5kwTyCUur6H2OjrHuNKEKBUKdoThlrBSXl1fMu7iRV3J45qyDOiOnq3BnHz2O
hgPq4L+GpsWOWH40dQ0ZE6Yz1EJ8GMP+paHgTq4V3RatVYJs+FgWoR1BQhW7O+ys
wfElp3PEANcUiifstIKqGMuADKJazLch7EqdOz2EGBOrVnumSgEmCr4CZs9kpNJK
uodkcNOj7peT807dCVwN4eb8czC2oXrk/W6V/z4hlXlA47iXM8RTVUuRzv/S0Htq
QVs6DHZYOhhUB8QQsK+ajgJ2cu3xdmEqjUD5FrEsLk/E8yEMX7a7awSYhda/eBPN
mPFX476Diq/LM7Qg1V1NX0bXFSgE1kPCCcR7vSN3pPuAWAC4g84fN73UiIS5WaOB
qEc3QbKg8WWHyd7aW6j299YKvz+/07hYzdVGUUq2XcFkICus0WX82r8lv9pqHz83
LueAbUn16zfZUFxTtUmpoclCM3mCjFAdRIN7Fdhf+3YV4ZFwpqGTp0ghm/i5zZqN
UAu7hVnVnhhHVzaz9bHgNg9FPmpNgKscxNt34nXMfZucypmtftctm3F/UxljCOWR
H1lGWDiwKpYDEms02XeZDz96CaVWGwIzg9VWQrCAf2qgq1UimUzbJ2t014qoNaTb
3bCPN1N4LbZUdRO+cwvEi+B8YRgA7tcmP+vF3ByZiTTdrh9BiKAudCg2gyqK3qPr
Qo2tDPSjzvIWs757AFQW4OoNZ7phYBtrq75tvAOP6oVxqO536rBZ6COvpzT7ijYd
Y4+nvzcdgEOdeEXsZKdKt8IiiVBmos1BovdYN+xrUeUfRpRrVFWFTaiyuVyj6Jez
8UHVSpROCOcfNvA0Mfw1WC233A5ifyskXxFAxNJnY0PR8owKL4pMhKhTHDsdzar8
vH25IyR0P0MO/KDKXkc0r4b4cu3j8+TabncXYjdI5uYjGKTNZCZmz8YlUZEPEUmC
KnCb9+t3/WLZkXngWgHXVzcCHh49eMFTVwH4xnQigFe9kUdnKekFCVdMVZD0Yikz
AdTPZ1hKyoGEzqM3fDGh+ZHmwfzAEKNydQcAUaxlp6v4y6ldQpiXwovJ3RXd51gp
4FVzvtXY+q0W0MKabKVZ35eiQI3fBadwpxDk0sDCp3xMMqqpHeW7HMEStrJ5Dti8
N37Ovg3uAOm5JlWmzW6P2varcPi/TI/DYa9VIRxYGClA5DXxYQLu7W+EjHuF843/
NHWZtV/u0Fg1+FCigFyeahGvkK8Y11xX5umicl7GJe65htfshj5aArdsjShlPB4/
veH66htbLf7ROGLHx3pxQJbj5QuCByIM8MuyfwDK3RKQWUzPDMpCtiBYCSQiszVa
wpOSKl1nE7IvqH84halLuW7pZDv3Q/p4+kujpUgMZ2FSwTYG3vVFfuhumjfb70OS
S5yJlTNO7iHIZpIace0r0XeeTp8pDLRxQ94sgmjiL9pamvphQbZGdWIV8690/PmL
47l9h3V5tVuvMpVA8GrxkX75w5M3Km6h4m+P3BH6KXxPPRgprha2BZ/OdV18gTo/
XyaKWDoZ1dAtkno03IeG7xYDLLCFamS1148jZaCjZYGUv0/hBVD1jTMig8uBPOcD
w/r+xq1fBMj3z0CyO+nGO99MoOZ0xAkOavR+ThQPbA8LXVIBT94xR1FFKO8VIsIs
dlJvMAefwJEX6luFJatA8x7fy2FpIqbNqREySOqbjbFidPkDSUQDqJ2xG9lMLBVc
TkLt55X77Pn+VTmCgOF34pWAUL7aW8Kl2btfwitRyIntTs0GE115pswtVH7760Ta
VSYZZzWirS1Q0Zc9zVpsXHujMypZXdr/9NGPWeFic/ugtzRSjVDfrMOAoz24cGM4
DYKyMxOtB9WguWR+fX6hcStqJWmhk3MdHL6V6q7hjBnhPZXSSHyZVA9OcmaMrvnE
4Q88FmfCbgxBEX+bLfNhGg9VM6HezSben+0cSRy1cQc0V3wfurHxrzj9glkPqlJ7
e9WX0Y4DkuhrP3Y0rFxG1ZblY91PLuM7moCD/1pCw8apDKr86851hyju7iqGu7J2
OwUzvWqAz4PoaZWSXxls7Qp+09ibJPOXo0wbogW6WoRWa9GIEIWjA0m7aj6hvaub
kVrDHWcQzVX39w4ZbjG4eKW3ulLVv5Xk9hXJQ/SaPwPBEdlmIIvoF+wmRNco6Ids
XAqwjbndcT7wu7SihCtdP/k3+jNCvT9wiG8FSFjLR3D7jjrN2Lfl7t/X6m74vdsI
RCor9wlX5QF/6e65WeNWlEXHih9eDFohNxmda3Hcjbq9rFg9bVNqPYOVvP1Ei9W3
gvHqwQxLlOVyhFjws52S9vjfwsWzbXnCpV3+X9DcmVdwXRA0uaL56AypJH35ZT0K
7SEvOktTQSAVqMYQfLeOgkPcwY/JnbJ6vVRc4fhbnFKj3ADzWCnQad0jhD0fkWlh
+fDtRr3QSaDRQdigGFq+fXLw+VAmihP1rXRL68mLjVMnOTXFlXX+L52n62N4ev2G
ELfQol3+vnFB1xcEsKahYGenZKlQW/hvh938O0VJLL0oaCRuC9TIeUQI8gQrk9P5
vyq9ZLrVhac7CF/cT9cclwqYZn8cV4XJ6DgqBb2nPbWtRSylY0Ka+k3IyIQxUUDN
zuG/ExVKfYPrt4pdvsvLU2ZNaILaHgeyN95UnkTprOISMDmenMhFrngsxzfVxz5C
G/gFEJrFSJQ2RKRrbNETW3aNso17grfp2RoFshZIzGljcJDpYnQyUn0gFY9R4xoo
umk2yh6jx+K3GKZPkiHesFL6/iZjRQEOJBlZTW1u4E87zRZcAz9DqFaA2mVJmYQI
p9nIQLvKRzuMGVcGvJg5MuobTz2m9ZCnZdShp08lfhyW/roRSdotcNAECEpwSVqV
XLHQLHPmtp95Q5T9LdRvmFZNcRwnNUosOIYzRbokzglA2KFiAKhzHxAlddogFr0e
ta7QqicGh0FCJS/x9b+5fgsKDy3KSUY/d7IaRTWXg1B47NQW2wV6vsES4hO9O2po
u9qFcPQY0Wh9L/fTZSI35fZ52s1EZcrDvSKR2UqGVvKYA+tX9BP9qjRPZ4cZfcTC
oMZbCXsQOJxcFQTsbo53MvvslwtGzI7TLL/SDLZFbwwE4kPjncMMNRZAiXPB2WN5
Naxid5/r2NNqaEkI+She1T7QfarCPRuHG5RPQSOatbogg/97uaaxvJGKYOYc8emO
zLSVZuerL6Gbe1fi89dkudPBq9N2uL+T9CTNjoTcxP9vtYbKhA7wLL1uKTNO66gj
mJJHvst2+QMui79x17JURyDuWWZbhpIqHZENatbQ4wBiR/5uHWRZwa5JphejDtNY
m/lZ4XDlYMFIVAPJOIUBpsJVwB13Dl/d1BsBtsKtyhp36yqPU26ekCQWvDUCyY/R
n+S+7/kzmq3/KXfAiCeTMO4YSAYNbLXNrS5AsppI5g/dEhkKRkv6rIhIcOU7dGNQ
+1zbGPNCU5C4YUpI/unGUFw5wIOAWQTcsi1wlGvt9O3x5Yqlli9gO6jgMFnECU0o
KhJSEbsuRmRXl+AFQe2eE32Jtx60s8uH2eduhblZbjezHLRuZJAqv322h6JxcJoy
QKWYkzUJaPylF8p173IOW3ZLQ4Ef5uzKkTDJVGymOjN2K4V3tP9pfPLMQfJue8td
lV5R+JBmSVozva6dJ+cQr04VrYDVM9KXAhMes2a/CIibYcqxSH0AUWeN/KbJz9D+
AXKVWitglRD+ARHv7JR1RoQI0/v4cYeJxGbEnYfbRiS348XkFZbRtNKNWgNn8lAa
Cwp1CIVa1Ui6LBEA2nwZPOfCcLUFLIsM/GS7hS1fZjEsp3YWuqS5ZwKNKE7112Dl
7+SCrvjydRbNJNVp4i65NuxFUtrekHGcve+gwCb1Gv0WOnySGyI7BrzJdtsoTd3P
cZ+zXBAN6TKByv7Dk6jEo6KfHUDr+ol44SrxBCSiGxeXezE2HWMrfLUi8GJyxywv
Uq8Ni+LblQifYYjIuuc9LHobtN+PXUnAieXK53P+tQfwUlhpC77zcYv/FS94JZUV
HvbV8TcGvzHKkOfuvdb7oICYgkjRjH4EMN5SVGzVgPjd1N1puiSB/N/PEM9kw1iF
DkEQmA/SqMoVI8cOmrFKUiYCk+ttG0yYvx9kI9bNx6B+vhu7DiAIO07vJb6gTuRZ
5cjgB89o9NqRhsOxeIfyK53vXYKc/5OmMzBFb4QrloDXo6umkPonLWuIx7kpNKHS
EBS1/OjKa+RjXPxS8ftSmxD9sZLAjb+BCN0q+yXXdpPD8xhbsEs/n/VSSic73fs3
+xOeZEcnqdhqjZA6dOeMIbexVLYR81ykgb3qqTPhQEInHgrqdjXslwfD0v+6ZaBE
sAQ6xZTF3Kx9kiaZO/kChgyU8D1MME2CGH0LQakke5EtCUta5XHBPe1B+moIeec2
0GynUeRtYPlEJ2Fs4i35yuXSGpyyTB8w2rFdTAn5Nv9PEU+o+UE+3Jnl5/GTwF9/
MDXouDvkzOkzips7Dp6iUB6UnEljiEcSmfDK4LJY5q2khpNulBe2IZk4oD1UwhXD
vU0F2f6CZ7SdmnW0yabwdYJwcFCOmu8ppisPh350P8Ax3ejwCGv4S3x+i20IF01t
SQrdTmMUTd4ABZ5MJ/hXDFTPiFtxzmgvEyp6AzdzwXc4deb+NrbqDrLPkmyVk92C
4joe1OPQBWycwWC8ikcJvExzl8/AWqeoQS68RHsznG+b+1OcCdT2KyZxDx2il33a
8lbVSV2D02Yo10v/6fDuvsC+PLTKBA5YbbolVbKhE4G4ALqjjhqXW54sLIVaxDMS
DZbDMubWhG5WSPR0uaGQHa8kwPEYXz9N2LMEBmrn9Z1xf3VIBSKzNWeRcWZP4hGC
VebQxC4MRXO+r6YpGg8tBZ25AVsXINtdb5PJs2oWtribXGFP+HDOIqEZi2soaZRD
wmP4dCJMM7FScoF25TAv4MevV1uWrp40RP1jFxcUgXYNtgpw6TkoEvy1As2bG0fg
mjTBpHc2SW8M1P5BSrolzmbmA6y6TeNH9iwS8+BdCLW+V6dNTIy4mfAM4xS8PDYt
/tIWacDDnKMSjJeymYcPuEeMXhslwRdwoUZvxf1Vv6abcLZkbiQ/xI2kYvjOLj+T
t+RZ9hZGL/6zveY9rI53hJVCtZpD0asCxFfMDIeYoEBMQGqjlVBxXoB0Mm/tT1gF
lC6ayuLH55LOnaLegw/n4CVPL1r9mj8TnakyQNa5tyJPmyaEQKWGlrP3Ts0kHJeh
UiaNq0MqUr24CC+fJv13r/iVDq1Ic+80mCBScMxWGZ2UwJJZihd1LSk+AIe0m/eD
yNznTWVZZUSubX488HUw6Tj88zsk8xEIo5IlO0hIbAK6QioHn2sJeswOs1YRrWL3
go7YRkos0D0aJMBLd0JXTEIyOrrzBc+SUldq/7TV+s/aXPZ90gn/zUo81klXAvUj
hmF1SLBJmvgxbBmOgpouzqDPN2kM9IqMJLuEjNkB4TJihEOpi9/+MOOtIXz9nL7Y
gQIDNAZli8gQA2QItBxe55uojXXl4HcgKcDl6q6O/zUn+UCjcADK84FKTq10EIO3
7lbki2JKjAPVcdyTFAHfDj8jkYjY4Utxbzc/Sav7plt/RQWIdAC+cOMv6wKt03Kc
1GhmEO7zgSI2fZTcs1JN1QUO4QXiZR911Infy1nYjCIbIdBu1ZMq5xO3bYUwJzSn
46V5yXg1YwKh1GIU3AbShrJQa5qOfPM1eWoQNszUUFyg3LtSPzQHhYa8cjq5mmNC
I7VkLeOh+lu1tmXak/jwXwWXmbFp0jpDJXlFszlP2uigSz+KNhiny29cFGMBxzUW
nr0kbv+GLUjG/NHsXQYH3HcSLFVMNjMpJ3GlmJ2r5U/XxFE+H4DrGzTeRZG2Vyp9
o8QoveKdcSUSWgPWv4glMSfRd5gtCRRYRwMfdKDIhJyPT2SzegrKX2CLUnCmEa6M
X7J9wMlwprc67//X+pE7fmvNwKOOqhrDsRU6cOiAHFeRp+Jc+VE1JHrVguuPIepG
zNdy1AOhMuIH2eBeOLzp29ag5keI4brTwMY/bBCm7+eaml2FBZPFW42BYlHKS7eX
Ufz3bM/aNrCiIKBKQEMr0R4GqCtu237IxaqSr1w1BydUUbx25Gz8qYxE26Odj+ns
fC3+qb2fVIWZkbiltbSiaj5ApPCQwT6KlLHcf+31FWPO0QZGu5/hkcatA3euxxEZ
p1DXiu0HcCfAJH5e/AWqaRkXtzRmPWQ+sLu1rWOhvMCH2dpJc1Cs26Hsmm5UKz/n
DP2jOx5X8E65Gjtxmbb0PzevNk3xDx1b61KvJ2vlv84x7LCaybDrsc3D+YUinOK9
Shyubn3XeuBZJh90OOalv9xmKh4sMPx9EwRolwBEcjhE29Hj+wVv0LJlxBkkjnXR
hLvv5AfRNJavm6Qy/KMsYMzvR/DAW0X49x0cQNPdf3g5ik5u/ThwA7NqKsXv2IeA
hHTTy9EDBcs3kTRAS22fDUye1u1f+Ad7dRNmSaNIS+UePLf8e3f9gNXkJ/x7i7CL
CRNYHdIph3tO/Or3BbGi/rIEgwzdEfaFfyKyFs8h/HnIXHz2aLYVF0TjBMUfeoFG
DWvVctSnElfPIMv+Eqrz2iGTH4i0lbv7+zm86JzP7VnfOk+koyRxKrBpW17nUctq
uhpEA9NG/o/F3nbbyYQKYfWtxG+EirCavlbC43UbbVUYYBJwoXmxcahE+ncHa1vo
s7FXMSQqPNXD7dJ7phy1h5G7D46/A/EtooxIOLrk6TTwP7cGD2HCWQoU+AjHAYc9
kwTsUta4y++XmONlev1Y+ThV0wPpVUmUH6KSB2bGpNwh7PFpouz776U9f+SxMQXx
FobvCW+AYacJUzLojl0rCTDacqLL3nxPOCGv3H8FEOV2D42EFBQPHE4eb2iw4lyq
NypOZtuvtQkrF33ewmbwiFA1YtzIn0eIU86EkP/u49ROKncuYf8+3QP2XogN8mWJ
9IMoWcXivD2ozucI4lTnfZiEqOY8sYF8+mPZ3EmAvT+3l0Z6rVM6uMcODGIjvjrj
7sCg2N957VOj758IsMsOqdIUOiEt1l2TDEkkgjxFFfjBLi1sNpCaiqHYhlHixu2g
oVjUARsFu1bpiHz6ic9brP1WUTf1j3eWhiL7RnJwHhDq95xH8SaPhal0bBOWsujx
s1VGKycdFneGXxDBs4CDmRGYBuaK804iZHAMgT/GO3nsN3eklJBPsHFVx6800WXw
4MyXZtvq2Tb9MGz3Gjt01nhPUvHcTVWyvj8V7tOyA2AyYdH/xG2WMgScBWsf6gw1
A1gZS6DvU+Q7MjjjV6e92nSAOl6otEph73xBalQ1vZ6WRNzZDIdow+D+Dr3uLsjF
590/vA2yqg8TU1AHLotP6yeYxI6yAoortgGKXC+zJ0wCAYp5VBp8HPry4sm2HI9p
Klw9s25mT6ojSB0rZCIwAKrfKSwC7H8nXY+bno4/S9gG1u2M4aJaH+z2tXZmTYTE
uNdXEYeYQhCAZj6SqqhqyAz+qoEnc9Ps+tqVIrBPYS6u9fQAjSjwe45ZiAKh0gZU
nuwgTbkn3BqzunG4rm4n6uzJDzmugflRVB2i2LYrNR9mf6wYuy+mUJGQFP/2USIQ
ayRJpxATuQ8iEE4mXSI8lIqpOMwMltSkCiWTh/jZUyWvy5YIKV2Y/Qh+kZ1AvmWp
sSilhKsrg+YYKJLro/t4ZlY7N+svXJMzLYuDB7ZPrwZQBGqTQjGwWKxmBKGdIrJ7
77WjJ6Y0gEnBnVELw/TvDkO9EfYba7C6CpBP5iJjNO/S1EX2xgtkhVeETrtIUA9j
oAeRBIwIjplL+btOBizTcECrILNTQbSS2pJLtg+ckhPkUAXoURd4BK+ohfdXkkw/
1SqyrVSg6qhHOB19V+O7JlwN1mBzn4PtpH18E6Zm+4AXu55pBuBd2wqsD10PU/cr
qtz5CqpKdeG6EJXQa5BXDNKKswCYet9iqK/Wq3+KjKjGcsgkdNORdntNXmYD4pq5
2W93Y2/OZrEMR5undRTQoqVah2nPlD+IAXUw3QkIzi7Q3Kj54jiS6k1Iy5GMqsaK
3hboE1z8vL494JTOGvXgd5gkmRfPqUon2PDpwzWHwYypbEKUFTRFgAe+9bCF/8zl
jOJWR44OqZ8WJpaTv9V0gHBTyXoPlxJGHqAIjkHgPLvv2nTrmrTKJrxgiuPEIYt5
ToH6S4HCN1HZlWHdSy9LOMJYMOlISnyrj/3W8jAU5mO5MYcqv5Tf3GQB/9FRejR0
k1I1I+73jEFtR5NU45qorasObBz/qyHb2UJavtJuPY9yJrQttYWll0XCoe9Q6f7E
5KwrXaV34BgA3g7D2gq5jaul8WLpKwQ3wbLjooYfqu7qOo5nnbzSOtwmWXTX6w/F
zLFh5irVZqVUwNfkwpk/JGdgDEkuMK6psHmES6FYkRgdRrQzYacOKO6VGG9R7Wsn
6FinYME+6AL+sDYmnSurH5cjjqB1tGDp2ze82akQ9LL7lGR1YuVKxJ7kK4BFGQvE
4jidQpnvDCxN2qsaIn2at2i3nlX8w8+YztRy6QGjjFI/cj5RR+svrtnagfa9Oidw
HrijWwow6g4dwGtUsi5DXMCpdl3cuM3WDW0nJWAuMfBL5kUTmas8PocQT2KiL0O7
ZshLLQYeSuaUo3+9YcKGe9kYyBAfbjxuFlgKLPph+GtgG4sXJe8AiAGnwxJ7UZ+6
jdigYVpL/U+/l2eNwi7B/rV+DeYM5z+teSI/aKVdmdfnPP91MbTx/AKBM9BJhkuc
CBOPTtAZYwAPsLlGycvkE+vdygh/xqkXJLd9X4JTyjfIwAtRjURMBHmxADEHjYOo
zgsNDc6wJXCSpmX6S3SwIT5ghIjBf91AIaCeZcQsjLE4Gw5buNPtf2WQJdtekY6H
ZjnRUTkBN+dCmoQCiIBM8hFBrkG/CKALsH1l9lNw7lFdSJ8haswQAyh7xlpb7TRR
Id/bTmRPdrUlwIK8A9vHVOeBYXy5vO1eHFTeX/4Z4bVwiX9bfl5F1gvKHBohKH1a
W211YypkA2SHAiH4FHggUwCRNiCRZ0Ud5a3IRci2MDuWMA/RzMjjuWtb94k75NYR
EdPDWUxTMpY/OZGrDX34cSGfTgOLo4Wa+E0Bk10xhuqFdzACWxdRQn3u467BRjfd
yDkM4Wrrfj1cPMFro3woiZxgMvMeJOuNmpfOvw8fo/noscj8f5BIq9Al2KZWRC8K
aK6zodJG+aij9ojXxSb2cBvk0eXyMNVhrPhnCcOV/uo0Hx+x6lfClpKol+01Eopm
3qEJ5TPTEnDlql1I88zSBcC/utsgdfP6Ax0F8m3HE3tJCOqx7tWVyROjqD+n8bZd
j1vcCksb7jmlFvnuigeTRZRv9qUBsX1U84YD7J+MD028L5ay/FrqMAKwy3gb/uF1
6YN7W/mdMfh+UWLV3hljUUm79mnouPTB7gdGSqZFmaaceTaMfJGyqnv+F0gA8CSw
riK86hY1Ukv6+1r31vfDhCzUxyIYYALmKn/XGdX86zg5uugqzSFziRqf4nkXTJeM
FqKl5hrs5ZlCbX21Ksi7+kEFhfhMopDaTeZVfJigQ9w5wz7AacqbYhKvIKQdZ911
lSe5gqLTNSkDbvwBJWZ9bqI36uMzEHp2qpXImGsTfYwaRWskBceeV1e34P3uHxbn
WYTEzPk1jXa3IVyYr13TzpOPc3QUMgZPYUCvNjfru8OXMS8Z2vwlQ46tYmguHkMH
Jh5Q5Q8/49wiVEcqPoUreqEAV9JYMZBc4b8TPG5ZMMGXA+62W1FiLgczP374tMEN
Mm2Jvf861Nrtr/gfij8lSw2T1ODRFuU7vppgquXlLqK+BfBvgSvje7HHNJc4kcGp
/gwFbf1ai7oHE6PjDuvJLjn+d6iLIeqRhoCIj8vNeBFVItf6zcQsf/OWZoTK3jNY
/O2K5R4d6b4hKuqrkzD7EY59rgDedizfKFxYeyNINUBR8a+Mn7ygpd4HkW1h7tRQ
zXW683oT8Si9TwWFH3wKZ2smcUk0mMNitNl8jZ/7YHVoKkGkg8c1hFrc5i2S+l8U
wjNEb2V5O0fPsMDAOq6MLGqmE4Zmnr366gUogLCwuqTuuPPkB/ptvxbKIntWTEC3
uA8DFD5ZAQTurlvC6uc41rfW4f+2kiNkJh4zGQfOH4y2I3eSMor5RRSFFoGj9FVm
zN80yx3HvEXbKJ0gOcPlS8x2bQqF4fO8uDqmwiYE7vkyGGzN4MxHVlLFkOkaNO05
nz8cIwj/mDnFohMzyJ8oVflHBaZyK1Rh5pf5jPDaSZAabZ7AyjRjSt7og/NvatwI
maez/PtLDqczatDOX0uIE1ezmaf3PylhhiLWPL3PrYQLk/4Js0OR0E6nQZGuUis7
aHsajzh4yqFu2gtjOf7NahFMi/Ob47j4be7v/k0nR9y7LR4YocTzNrNz7T7eWldZ
OprWJfR1ItL+aF+MHu0PBeJ+yJbE22zj07Y7G5kqPEx6AkLM59cC5ARcnUCKiKld
0cTswebuwl0CYL7A6EB1ZTwNnrWZxjU8dumQWWETy+NlWCtnZpTS3sz1y3loIkC7
Cl1qchYWLyLUW6aourPz0AQKWh8xh2jPN9Ju2bru2ZLYUmyPdjV27+PicK9WN+NZ
mXfRs3kkU/gn4oAErDbFl2u8x+J2rDp4XX+G17FqkKYHL/aZ4zsS0SrS2XfHkqlK
kHTN+8BFRW9vZmX9S/Pg+SgLWkYSZ0lrRU3ckqxuObhybWAsqqO23I5ZxpQWlUcW
gHIcg6Uooo7anR8fFMjaM/iwDrDUB0UnwrV6Y20ldzL94zz6BbmoqGuz3fLfITqh
PLp3FWdygVfweVladh/zRcdbiJhnlPcfHm+hgUWYUGR+9HbrAg+1STOPSAnvBtIl
Lw9wBPtX41S+9M3f2mWelikb+yJRhttx24UDjrod8JTTT11Th19OWPTtMGfGEPAv
ukLO98rEhE6ylbApOTyxuSnroqFzYl8mP5cBjyhdM/dna8cOtqroLnDf/ZoQlEe2
0+c5uhBaE24CeVQ7kG8r0W2FuEMGxuS+O8zQM2tAsInaxnnOA476Qk0QhrcCphRZ
2q5O52jGctCvcsN0frrbL6+bHQQp1Ynf+8gFWAFOMie+KsEIXwavOPW+zCn5314x
zs/8zrsfiKDUpgozRckEDA7FiJt2ZQr896ssFiNIUccEYagt+qSp+vkcUSK+2wAs
N8z7krKB9o+uvwV7jxsXkuMizttG/pAJvNzII9/ZhAIxRo5dKSj7AkNgHfZqj4X8
jyOPBihpugnK29hOqfBfA1d1DRYauGQYOBbRe9slTDXPky9ddS6FpmzQZNPjeji2
yOGEgm9RB5P7d8eu2KgBKasncoRajfkXqLjTAUs0gAavYTO8cIkjKR/wBDhwyA8W
H71VoNqda8EBKBBUUjgmIYHyKE2u9KGL+hpPF/3AxDpgPbOMcPRV/HzL2EbZwaCK
HHWzsU++/gWwHnnAEjKMbfXawuq1qYJs4yQp10iTzJ14E+8TAJysAes07fg73wjP
LoBRzr9A0uAfm8qMSTekeUiKQlDuYQ58RwMT0ZLnQc+djBfpt+RAnt0rOvTFAJw2
GE7poB0MVYxiUNZjdqj0AsVqJmdUhx9xAlof77YlVEZjxkRAx7pO+U5fGAgDBeqr
2Xhck4eR8Hx+sRqMAhB8gGqyNWLJQoa9JUSZf8xqBFmVH+c1EIyS+dpv7/37KhEW
IBhAedWa8Z7br6/jGKY5+A94aU++7qRi2tR/v68a6yT8/fmAixJK8/+pajwoNHDz
x4unXrE9x5y+UzypYQC3tBYnqczjQxvcn3lEy1ofBdViXpOLwJJ1X2StTa6ll9Uw
Gx8GNoqW0t8NdwM5I0Ys7Y40hqw6i+DPKMN3IniJ1kbJqDKApt7J19GQmnOmMsI9
661Hv/WyVcvz8SuZcZp8/gh0KP8pvoyzp/VkFgUhzBRd7z7k/VghIiBH8pgo3SNt
iBxW+2F0Dgd/XN0dr5iwpo/AB/E2pQRMIGn1aaHAWIMKdA98izmHHQMMPauqtI/J
2CbbqMc2T+UjRmV54/iDlQBxsq2lXwWhMqySkN2/Qsrxl8nTpQeKc415toqA25r3
sJ3/ETZrI+appF8Ygt2dqwpyMjpehhI7kaQ9IXxwJanZHw/jsVq0HTSxNrZI7KF3
/Dg35EJSKC+LTKTlKKjdiZkrBGnETHv/cx9Jgw++/1i7B3GwHA+0Ze//NWMHjDyV
PN+OSp2LVltc5MrpOFi1iKtgmFXfjfN+SJknVdROxttENM06n2nuQCEWG76CbkV7
ZJTJ6Rmuj6FdvsutSB2Ty0pq1NVXM3ZW0HqekXYr/gbPgdW5ZKjfZVeoW/x8RCor
4U+rDsZL6VxHYD/A2KJSm7/kSE+6levIh1b+KJvi6vR3jWCObevwgOZrZHd/Pezy
Xi7vWjvnzJoKxw1TplVtje+QiGEQGitOFW7y8HqLyS7JXfN61kb1vTgIYM43+i/C
kfoWdz/ZL37xhvlRFqtAiZJ8JEnbTutj/HDpVEy4WMWb7TrfnOnF3hFWVcWu0iy+
yMiHebkNdLhPOwrNCXXFs1+So63oO/HB4fhe0XtDZjaF3v93GGPhF9Pe6/I4ZYKs
kjwD8ULzL+rOHYQ1BBogaQXAXbM+m4i9VzNmGYCaAdo/+uYJ3t1xrVZir8FY552z
0eUvu9CFJJ8zewu2kpshlPWTAtsojlv4v0KjZw4PYHM1vMILTfAMtl8ri/ZxF+yX
jRCL9Z3sUBSOjFpZUPhoWZRyrwuUWwli4EGd6uV4JVRPd/jnN4JNDawegmkbhCGb
3+I6S3ilZ4w8RbqC5Bu/f+fRVf/dqpzFi5PqSJSl1ScJjdFwyXOKAG33pCYyFiO+
scv3AHs3hMeAODtuPy6v6dHRgr2o69byrFiMl17YbkMVAuIxNa8JtFdbNawprbAD
I35FxLOwZrUHlW16wFp1ykKZ4ZEn3kL0burwVsCSLxI5aKRJ4v8rHwjVYiXD3saF
bf09FlsA+6L1JcmzhqsVSOlwPOwUAm4VtwkCC8W6La4W0yC5mWHsczon8pW3IblR
uJO18kH3utuyFqNcop2yneIteLVDKMUj5B6upkaz7iZssx2E3MNXJi389mDiV+2e
z94tqBzt9aiyrEq2UulDt7bBkoJhklXLA7PQOGpx4VCk5wHQhFTICnyE8K86F0ki
nSQ0I8ktjAJzlmHYiOFo272OlSVn/mYfYrgyz9fFFAG4fNCXMCpHME2Rz1I+0llx
3ib/p+3rTbP5RcsNUhJLB7rDg9h7CnAcLahgVDPCZ3dQ+KfmNE8i/d8OAKa3BstT
EpEJbft7jHBPbZI6g8KXL2mwRCF2FEp9a08ZGcbD9KxacKpKGtQWY6BSv+ERgNR2
lb7G/yqubNDWwYehvehqBtpZt/fuHVRYsS653gmqQF5TDTmeNHV1oadalNvEKnGC
eVzKTiQK07lWuIFlaO3yYfa4oF/RiNL0P2V4s5n4o1u2JQ2s6Tt9jlb35ryYBxv7
kFiYA/Qpt+x2SbP9A4HOLM93ZFppnMoJCwZgluFn03v/RTTbdVGYYcC/zumELnRF
rcWHcZ5mb1fnjgT4twtUBg2b56oL+1N4yyRWZpFMGoQEKp/FcGfgaOwAmWM649/C
lapEHVIK228t+7LzEScip/dhfYaP2iDtGAJ5fgiGN3bwye1bxsK7dszruwo5uQiT
0XGuqnSEdDa0ADHjrWYObWOkYaPBGn7QLtBhQECOOlPZIWR1cNgMtpXkGyeayIcU
JwyTbXmoXfcIFzxOrICBRj22ZEkOCwr+LmsOK9XGuWHt6ACcD1mmQkEkkxoH75I3
x4Mw9F82hH1WForGgdwY7tnz4LWdhnPS7rlyLtcvZN2YUY82Qkf9fbbWioO79PU5
dPZCWSL5H1DRk5CO5Rrpc+hcIMKDajzD/bXxmoBDo21ZTDDb3wFJlc2JELWzqqLk
VceztnjiuQ/ZCUIw2AhaELNrZe3P/ivz+rlYfnuOIMht60fB+JHzNpTqCiYTDpXp
IogUA8dAcI+7vGzjKpN8Su9T6eppX3rt5SS0KiLBYNqdNlZKwuZrhn/p5nMRQj4S
GBal8+Z3FkAHwDDZVc2Dq1xWVBEpt2eCRMTHPyj02X1928mvr1QfBkQV2ksz0Brd
APcKL+h7r5bz/Ws0orWSdBdEheiP0xwQ1h3HS6VVmF66zFSzymMq8F+dIJD8kaE9
nhRBREgKsjPnxTuqGBtDaVv+mTYDi+ZCIIvqG9noSsxQsNXZpk1Rm7SHVdEYasyl
JjwPfopxubF7JnDbBFXE6KuaIy2yQPgWmEk/4kiARo3MA8qn1NLXuMOgBFym+rtV
fcfVs7TzAGjTICCMTEgjs29omblyc/OD9eE/R+qLnWg04KY2F4QxH5isXmL1bSGy
VAVU6J5z93JNeAaj2AaD4occ2O587jUZvNLLI2ZjSG3bJe5OP8almKx7uyXmUUhJ
599QxUKIcIz1jPz42rF+2ueA7aqeo3AfeGG6O+NaoDSxI8ES21ijA/O9aERGZdkF
iCEU0washcqhZQRaGWubPRYzJhwiTgG/s9o8hOeVRT996dQ7tjoEWT/n6Mdm6iMe
xHt0ZP3PhT5zaNj4v/+PwxqD1t+4O+SlLlfFagNjVFSIJ+NRGIGecUkiHVcxKu5Z
9pODfErf1DKD6VIna1GM2k+wj+cPOZI7mmRRsyAfo69ezHk+Gi6hOBldT+FtTMRf
3EeJjrFHTtgdGAkGus+KlNlDxY9ncLt9YT72nPOf7vCg8Ax02m3kk/F8Vs0aKteM
zqruQQmqBjTke2ac3AXxKQRcFL3oN3nA3/fG2ZBZjlaJbTNgkNgPI2A23XlGeUwb
gx/2r1hCjWxS1Q1JT0U4vQ5qSMbIc1WGd+wOFJ+j0n2cSFCUta9t+PZomGGvwM56
nH0zRN5zldzt+5mgnCVJZqsktgnAUQBzEw+k+tIIo5z/SDuNnAeI+bIMZs4EB8Lx
De/2YGoUUVMfn139Ar4mpMLapLCI5yNKc88h3msr8XKU6s2N8ZkoHhczyGm/j74R
riXY5obFmsoFx2wMp+cFax2nra14L7m7FH5CBaDSz2+kYGTGpN0sDikI/Gt1GT7K
6asgfx6PPlIPxwr9DA4/a4UwGZj+jfR9PqwpHwe7EtM9IRHIpPbP5xoPH11SgmaO
T7ZYX49Vh+NIttPNGMTlBit3Upgli3Pw3uJIHALsDvGvyBRjBhnxEzPzOSfLrgJL
AgelukC15S8A8HGoAtBC3y7cCKFZEDhusNFg8vgGj+ff6gi4VQFB0BU256LNK/Hn
jQTqjzLkdvescMUtzghbt5859zPco7Qu1T2Wrq2LfuxKuVKjY3Cnjqsn4RAwkbxp
0d1pEgi3QmwtE/2X/XedF6p2o/rBLk1SqcSAyUI2lGCbtNT7wAui00vhmdWb0j4K
Zx2s/5qOaTMHFWEOVmf5XF3vcLvvIJsQnSOTzP6p1kdHI5gNUKTA7G3mYM61o1Xu
Hj9oRbq1sPuagv2YOWtQ5PHL5I/LKSHlTa51U+tTvRC1Vdh+uXVNgAX/RdWYN3MM
9dWI+JZOFBTnN9QYYiBbCOD+W4nueTR3WhR8vFlM765X0N7vq4Zgfk2k7+YAROVm
a4nPeoajTiFwnjUUCzdidxd9MufKVMTq4Db7BVxYZEbiPMPUzTAIbhKmseEVccBK
L7qRLdHmD1vvNn/06Xtvp7ZV7Ah8epHt+74a24dpJOtL5jCL0Tx/kREuZNwr8JoS
Bxfz6M4n05gpy6JzoWlx7TonBlaxZGirAZ73rji+cucigt2+mOPqnX7bZWpB0nuY
1HuzDig+1R9KY42wGpeCRr3XGLMCwN5PvBkZ8sBfAs7ZYvZt6ydy9/iuF7bID2Zc
YRZSXU66NI2gLPjFo13GlQ8Wu37QcjC9EHugDsi63JUEgmspy5e5WNUWzDwUWqQo
fLTJ7HYc1MTTTvO1vXrf6r6tp4RSsm4Hkz8+Q9ieamdFuv1WkLd+DfVVP5zFAXEW
AQ2W4M6eNbJhbXbtjVjA+YybmeyhNFg2e/fPd063FW1HMjq/8KEVf1mLZwGNXVEB
Nz+hOpdzHpfyKNrpE/WLhN7Hsv40xRK2nBZleSgpXiSYZVNkKxUroHsuQmGS54H6
jyS4LW0saE/PSSxME5OkSpNKp2fMQh4/WE82oskzLot2T7LMVBP1+1jzu57nFMHQ
7Eu3WDo2RVXyR0BIdUl+LsmJczu53DBPGzg68Oe7T0uLMOizhTBq9n2D1svM9d86
qbJtfbB9UW70CxG33wejeRiiU7RCdknPiJCtKnooBlEcGfvpxcIrdZXw02s+8Yd0
oBNVXDl/kjNj5eQsie2cF2VMgUFzzq1QAh3m4CO6232Md0x2NaRDzjwSBHqgB7bT
FenUcNxiZp0PrHvjs7i+YMzcat94mk4Rndc6nCd6fkQPo6giZuG7adfcQUDYX8w4
uSof4avjUT4rAExSNURqT0e3Fdfnr6FqbSx2pl10Q9k43wvhYEfnkVtBkwLqiFzI
mDnT6ImqN4qyqBZ/RxryQ1jGSIUZCIdxuCtlB+R2/kiiPqT6ymw4sb9fYKbqvHXb
5D0YQ7amJ7XqXEy1dva0lboneUgbv80CSs5VYHkn/zidclDKB5fGqaPgGxVviygX
4uCWrh+jFYQVIpoO0ssRBA91bIR5ckz3OaElSYayf1p8v4Ba4t5TPO8rcxyM2XwR
I6EQcGtf8WiDPg/4SiRMZs3NwrXEkLCWsdnh7grpGxsgdkmvH9rZowGXjPQQpU65
kc5AjmXoMqlcEqy4uQTn7LsZJQsZTP8e4C9/iZYi6XnwepqNdOru4nuljRZmKXWF
Po0lW9NmtA/4kX7Ei2hZ6LSbbaSKFxkqc9NjfxCQk3cghI1jYmloOqAUZr+i/KSB
3JRQlF2TG+YL2lxk1UpoumkRwhmo1+yF6IL8TPS2n2IBx6K5DidhMaVSRXVPnPa6
gaokEhKpdbx5bn34Uq31wpguoM9J3Va8HOZwP/1uNRl/bcx2aaYWtX7M3zxRwq2u
mOuyvyBDMSgOhxsexWbLZHzkowdT6Oy5NxaD05zrTDQjeTCfl/DUc7isTYEH86+v
EZhXnCac8Mxvv/5OGvjt9ItHPDUZanOCL6VzRETRXQANqk5TQnYkl8rBfIMx/Mv9
OJKdU/1DQhexrie0eN/twKFNeG88QxWGuweFwPSgpqTBYiI90J1CeSxd8uj7lXRd
Ety5nlep0PeCmXM5buP3QJFitZHDtvl+MQdx/l0BXvLMIXtXd/pWCbUtsswZcjZ7
ChaE+3IQ7IEEjfUhvK81Dembj5vuBGOhYd9iPnen2UoberGTbxH0e96eqFcalA+J
V4lhfGg8ri040Mpf0XlXhmkBTnSAoSMbbw1XMXYd0EMH8INgUztJSZbreBOraeH2
8IhwA6aMt3hJtaUX7mYyyjugvW4ddHNkZ0qzFG4+Ii17Nrjf1i9zsPmCUUDyexSi
A7C7Iymn35UHkrlWCXsOCi1YmvKZAf2xgDeIPiVRu/pnRIXlVnKGYsXJTbTwRgnm
s7QTs2cy3FSi/W/KYy5GBAZ42KUCAUJB6CosYMdjiORr5xxwe3F61ONydbwgZ1kF
1gL4D2yaeGmlg2oetkUKxRq6eEG+xoXaiGh1tcoBhXJTh5PrMmEoqr8J2iK2LwYz
KgTMfrWu/q1lmxy7K1eY7wjqi3MmzHQlcMwMBxAuM66pqoQq2hqAlzSSQMRXkbsW
DFCsLZ1fVXPVoyrpMHdVZHpbK8xVNIpYZQOSerXVd1DeA5J4JMjicwUUJ+speCTv
5v+fGOvo3zeNE0bx6XkjgTI4AoTznoin2ikdhogPSV5a2SkMrGg/Dbk8n9PebPpq
JTSKBCGlX9KfL93gQKuCPma6xFBpuhTLf6+KEhFUOqaLu34ORYvw6/Yfk0p7G0b1
QkOmY9O/mlGdaS8fMeSoXs8SeMKQxW1ztlpF89AjJafTFVapSsBlgHkWQ2ZIcKG7
Xts4L/VvNn6R8YdhEvehofSTZfhsfZr6Yy9gpuz/6h69IdwtE6iJR5vrgoBt+SM2
0Gtwwy/P4aJTp7yUy/gcqnbDM40eHY2Q4vFqLcV68wZszBsGOw1ClYkqdpdUnQOo
f7A676GbPU166PeFY3zidcSeD097lo3ANjxG8VEYetN7pyZT8ynqJZD4g0EoxAux
8kuzxEKIeuM+CJfTJc7q+ht4fYav2o6AFr4OfDZt16pVckYmzPkYeePIIds95aF4
XHU4p2g7p9kv5aYfWiDg4eX5WXIEqvsGWVWrYP93Q1tNYC9Z6nKCO+Ppe6Fd5qXW
oYMiE7knpQ9Jeq/sLZhORp695h5fmadJvwldmvRiO+UJ5ZZqO6XqFBDJFsp47UxW
q2o5feePjTgj+KS8Cimhpc+o0VP5gB/PeRGjTS2G8rMAOXqEH4GSi8phtr8jaoRZ
8XkmD5tGtdfalxgYTXq1ugGdy1ak0jfurcjH97XNvVVYpWRsxSbfV6dqWydpra4h
dxukUHtRDIICOWwmqD93M0CvrEI4Kz7HJYt1UsPd9Uz2Yhy8t+RKo+gnRN2Sa5kK
h5DCZZLCX3jfhhYn3bn/nxrObi6cOtA/guk6ahS2RnKVFNEZhyY7JC3itDAl2n/a
C7V7gtb2a3G7qqIDa7XvCcb7ZtwWEujHlPpYnEyTEz92LYaNlcUt30MLOWpIYwSj
yhsXgUC+10fgpa0JY5STo0m4amB9L16na90DGwN4PufWmjsqQVH4Hyl6tQl3Kwb8
CLtlXKK1kWiD88ezerodqbTEw4+Vgu0IHg3izC5ODuMNNyjtI5glQufgbimYqg3j
H7gnUIDJPQWG+DfhDBEBSSN1sClynJgTKRjafDI4JoBdNWC6qjuW+A+2jPoFCfvl
2j0BYZdl8CBpZU633DFCxZrJz1EQ7YetEIEYRfcnsnAuE+Q9ShTTV+bhmVpoB7wY
ge4sRXXMitW5pFc0MZzZ5TAUjDZP10qiyETAsWvVDdEj3pTIAHLrBg99zU2NuBiA
L0nmR2zF9kPHEqaG0A7zz1av8FwfhkXeFdRzPhfELdOHsQ8W8IKsgwf696M4KGLo
tGVBusscjhzYJPTQq6nNgYTuMoS1MA5i3FV8cer6N0otBdTYIfQSCPkAcyqvcWHH
898YflENHZvosWJfDfPQ8p3UaLEi4jGfMSY9PcAXNtv+CFMZVM30yAfwnzGyhU16
1OXpZW5HAEccK/wdGfDbAdBEXfE9toQmekab3JVK/mk+i4W0lFzALw1ZwxtGPBdp
7s7cFrSxfQ1bsuuGf97XR+wQlK7axt49bQoe9CpLQZLWY7RP7QKz3ieDTOCDsmcH
y0DgCwo1YJ9s8v+WnIEb4Uw9TM6oCypyf2rG+tHUz6RliK43FQYWeTTgrVQ1BP++
oh2CUVHvS28wgQIkeNSynA1D2d0iJd+i9bblLn2fYLoG3+YZ2mgbL3aRlfra89AD
0N/nnmlWeFOYd/88ToiDeHs3ZvK9lfiuLIO3TX0cFcDqWQGBl/l/aY2eGjDYTMI5
9pIXoHbp3t8nHKRDyzE2eL86nT69Ipr2fgkG6K/WCM03Ktich1FSCQTp01DRH/ce
RsrtStbVRHiIo3EVz+wwzwHBgCT+ovdnQrjqOwIRDNl2kyzBpv+3Lq18rL+d9lfe
0+k8sIdj6eO53Xwj17d2vRLVoiKorECjx/GH++syMzdOs/wjQUKm8GYFZ6PDIlQc
3YjqKcwVq6XwbRpvn47kNfLifdawE2XHsb3OIMINpTkEDBHha4LPAOX09g4ygXpU
q7AzrM/cvVg/HQgXz+8yHS1PxWQnbtVBf2J2kYX9wzq8HepPeGT87kfPt8z865Cc
gzWld34BHWe12fcCdk0zRi7Sw9sOd/PH42NHFikUfKmQp8ZwuMz2xvNcOBqmXzTJ
AkaZqhpLUECbg6upuaYlz1Vfk16MEFbBf9Qyejb1fEvLh80d+uGgNyJHY2RU3Juw
l6jmTGm3PYjJoCmMDKpWqpLG8DzVZAlgbSK0d4atzDHsPzO0/gD1ZjCoRHgLvOSp
6T1LBU/RL43d+ef+mpWMZjCuBSZ7kSTCClwDAZM/MM2NB/5klcEHvkj16DcCcz0D
yZQASnaCA2JKKNQGk9UCXWRwYHCSuCFJ4gRvgVTObcrFJMhhLuWgkrghD+rNbLc+
VaqhBba575fhYyOarBc/jaCUdnY+5bW5qv060nbXogIS3Nk71h+GvfxB7nxW3k+C
Rll6aYQnYZLU+tkX9a1FRWvO7h87rXPKNmvlifc3gnHHmRethuOCAIlvJh3ZRXrq
hqxw3eLMFfHylZ9Oqwed1atfcsuM1oJ2es9vfDmCciN6oEvaxRkrOj0/TX0TKdKD
60psRCPZO/CrgrhbThr1JV5IenSH3W/K8mGdDnNdTVaq7BlsSaWS33ytOt4QT4qw
dmXAx0cQExYF0A3J9BBg7qrAdpMW5AZ8sulpm57Gvulcv+X4z0CpPUeZJJlEWLld
50YNIrfznfYshoC+olsPTs31D0jzl+R0aFN+O+/EFYWLsAAfd3lcz+xcqJG2/2pV
ZE//yDd6vnsFhtVdn2Jl5mV+K1zwed6Qud3h1Z5kN9wzUoW3oybugk5ykxkMf3Jf
TvWS8+NsPezcwgLzPBiiuMzCoRJkNVi5znojQ1WZqZ/mRJljogRQkcxGT/QRYBQO
pndJOsBFrB7vsj0WJzGqDsy5WZSUEvdDMVW/RWO2ngIu/hM54PmHoCVBL528lh6i
zNE6NE33/N52Ib+s/KQxjVkets9t+1rgyKCOZ0RtK9tz44HLS3xnIaBsgSnch1qC
j/yK156FgraYakMc+xph06DrqHmRcYMzgFaW4r5U9STb/AH5pa8m86cuXIpuEoUq
zaxVbd+R1QuRau4qW7lke4o2GDIAAdFyQFEn0txeCVO9Tuj+Txoh0QXMYo1OXOR4
phOG7ICATrRY/J9rNiz5AE4HxGqxNF6u49c4+1zfhGde56YKzhKfw3dl7mAIjIRj
c2X1yBrwT4FpYlMd0yvW5OGlqXSog47fldYmafKk0ixhScxe3YmBj85250Zq8ZjM
lv3Q1nY0iAjN5QnP82Aa2ipmXBY232UqIPyDaFUa0/WEt+Vj0ihoFpmPnlrm+L7w
8uwt2Qxr6atDjI8O1POKQXUbtfc39KiY6Bm261uXqzaLWBzD5Ea18rwAyBQjaeBn
YAk/vHN4ANVExMKDuY8gFTDU5JpNSytNXZCHnjU0zcFeWUfZ3GXLJriqPaVU+2KC
xYmfEKTuctMty9N6g9rv5aC+a13/xdq5pp9e9nlOQAcRG9jAqMUVE66FGyPYecnP
R5UQQQoI0fsEktqizDjaIc1la/FpsCkIH33E7d0XzwaOkzYRgm3+sorY7SWsCmPv
U6tuZxLuHPtgw1J1WFdqX9OcKXzPEHHDHb1n8ZmXbHjrKrqu/kuwOKObC07SSOJM
EdgKZFUCUvyCkltJij/r9cJGffk5wOE/6spIyOYu3vqkkuZdGV5AlXZfEss49Yt0
kriAmamUVCAqZI4BNkQf1QSM/Yv8qPRVE9HDwm+TCLNomIWJxBeaZaPbwN5+YA8H
dc//V9K0HV7EepHlAZiZaHLinYGdDqreJDJ5aTQe5+FqAvqeUfFI5jTHlRYWCfiI
j9fYlaZlUe1n+0m9EwK+g6dbNcdj8BugGYVTueY+61BdtQTYhKfurnzLOLfRmNUc
aUgTF371YZjLq9uY8aoGSnV+sBamzNgsSWEVvpxAEhG7vPHrOklMiqkqkX8+y1t2
K9nVR//HIKMgY5CFNj8q4q3nJcxOAFOFtR5zPzB0W1Itjhc5riuxlUy9XtL7OUk3
RmfUCs2aYUjxBRNBgv90xEbuxqB7RHfVtLnsnyEcRT3IDG8AlP+PPOZ/ea7HNr77
wZaFv+KHgoBzPvUv4p/17lcbhpjn3/4n8axP4jj22Brk67cQKFI5+dqdqKFVIZOK
ZfzYRTpzuPQCh3jcAZhxl8fkNWj05RyutA55cAFr5u6kWM66gZj7bIt7190aEz6e
9Y7UPA+8p69ghq3uFrFze3LYAD28Lc73ZAnnxqMXA8KuboG4GbuLNZSvSeAyXvMe
YFXvEcOtd/hMJ1tfLRM3mSSqarf5uL8JLYxsY9vV+fVyPoIqT4KvQ/GXSEg/rgka
KDKuixYockx6hKRjx+m79j1nVEBvkT6HItueNG+dh9wILQCxG7dZLUw4hoQm2tXx
qttqRc39lKZqW4IHcMT+hZe5L4Bb82GpBlNksE1/jvdoLO9eF63kvVhOmp2wAkOK
ijqsBtz8m0ZHCcyMM3owrVWIJI911UfTD5QH+jpwP1QcKlcsD53rvRnsciKI76SZ
1xNv/9evhhKnNib6dlioMZwztZe2GM6T9eLRIf4afwdR85XICQJhcR0oBejYNpdx
QJFqOEuXFxP637Ei8pi3xpyqwXWpb6pde4XFp/NI8HnRZbeW5A0aedTUQ5EOEbem
10kxfA6iPVRN7vGHn+pV2CYKoDBVpzVL1hSKqZqpvvb34LfZMP0mJIbsQxNELTjf
qMR9jGgpJXVQ/eLY4RVnKKuXDq9N/FTMapyt2Zmp0TPftJOPjFtgXSfIscHpmZyk
FMqQrMbS+jMMQROgZ+n10NT+skCY2q6G+xu9u2aF9dGMvIYpj+0aO5ZsjXUZ+3dj
OFdUL5llqnrdfeqXQn0YtPbqTj6BXK3msgaLeSzeON4AoUSeUBUEBcY7dzjA+foK
IjX68AWhBUvyQ19Zbcu2b613z2qzGwPphpy2kUQ5D9fvjSLMRB26bMJCUYgkkjtH
3F/8KpX5Yd+CYlxUlHLSa2ikd8o5E8lbTKTTw/3bYDfyhbUDW3ToRMFH+0srWzRu
+MkcXb8WSBvLjrYgS8cN5QejBorriRqadjQK9vXPCA5rQEM3m0LIxIWYCCc8idrj
yxnSznhTlgdqqoHN4gKHL6nE8bP+t76lsdfxDt0QFtcSHEOWXIhqO4jRMvXJoOSx
6w+VA42a4IGUxRfb4HLexKJJcI9Gp+Cg11Y7pJiVA50DZB00JXeih4+uPNa+rAtj
rS4OmLT8QEB06RPUBxI2njrUAN4duI2aeWxsH2CO01XLNryZCY68sfvTg4AhaChF
4XYtjiTrvoFsq85Pcjzcjt17wdNrcNj+5AtjywZO+UeTNEAYjAYf4AcuE1SHznEq
oT7m1EuuQ0yTnqtUCLOVqpos7OCBgqVaA93N9CcTDOmSG2gq/RcgiOEUIgvU4v3O
YX5cqNke8OK3/toBdWfHHdYrPHxmUpCQyRzmrL7PYN96H3+E3GgKpAmEXVTJQqnm
Vgl9RWsF/BLQbhHbqb1zxu/vSvbsiYET2BsUkve1dpb3S9d56YwEv0k+tt9gsZQR
AGyeZAUrGvfJsh1BkBJjqCVrVa/Ojcw9iV64ramf7+QBOfEM27j4IHvG4eYCLJnh
1jTef3bewmL1XfL2XeGBvfRq1oVaitUiKTbxe9+Kvalz7emTbEnlnZwP7V2JnmeS
AEt8hJW4Gsa+o9uCvuiHI7cysQIDFriDI2i+xZCOEokBfzG8146KOCBdleKM2+gX
h1WES/PDemXOMOQyExgkOjVbGKDIfBScOgJL02N8nYtwUDaS1ON7Q688jYpJZS0S
wBlPZQtC+oMyQANtZ+tele9USi0VNBzDIgvAh1FbH6a7kIJWfAX6JwzDUkpdUfMt
oA94GrxYhJkHr9ZGeVAT94nIJFnHdQHummtR4PMZ7ZuCNCnyMUS0gtJFh7YJpSQL
RDebYotgQlv+ZV8tGrSIqxqAu9onO5xF0Q8SvDpOG6QMNxx8FwB3q0Iq4/bqT+iO
BXqjGjLFMZHl9cIh6HuLhXhgsvEWBmVDPiB7+l1ODotyzdE7lknzVOx8hqM8JfpH
gzIJN5YVwGADJ9LKmrUR84ZTofJWzErT31t0pn1gF52EuMWPwKkOgzH1O0JwENjk
HjtKFSg+4FF/ou93zrusWFWaM7SGUavyxA2ZTm1lTxlKewBhAi5TQvBfxUz8iWeD
EG+f/u/n3+r/PNtiQeygZBht9We224V3TB64X4Ws2lGJaxvAzh0y51cei5qj8Aoe
jXh4dvC20i+LUIdsageEgtkV2sgT5vAHYoimqLlGRy6bI9FlU3aiZAfciVew/yGc
N3yubG7WPtTE0Hfg/4rriieU2Vh0MNVttA46hpKTkQqCcpo7gzIPJh4OSpfYAEIx
3BjB1WxV85QEA8DiK5IRKGeY1hiZ3exB9dO5kPnRUmYR3ZOh41eHCbPcY7/7581i
4E0g1j/pO/3RsLVKePdXqCmnx78YBpOZVJbGTSjxg/eYAaN2GQxu47U3gGCV14hZ
FIOtTD8sA2J2xKQ18E3DwRBdtqg/dmisKNQGgwo4tWBrY28+FIbw3FAbpArhWYBO
p/5Q1pY3baNmmRpEUHoS6XXMnWY0deSXJys9Z1k94mG3J4OaidRxExGHBVoF1XA5
BIoVm2CdXic0nJlYhTpHvs0zLPr1GERUEvMK6bdLssJU/b9wW/Y2VxBILOD1UZI3
jN1G+1VI7ucgDCI/izphiWWjnV9fvFXHqSkgIeqGwkY+OAaqnUW9onRJXzV+6nSJ
bkcEfWgGKIpj3+FMdd6g62JXknK5MDApxTaGwIiD1QfdpFd4Mwk+AibXesdJuaMP
FAj9KI41RKQg2m4/r8yABy8uEtLYlWeYTG2KHNeEW4Pg/5pYgSfoXadrHxkAiEtE
Vk5wwvD+Q5v3fnPCHhyWcYNZWynsFoa9EAysUFYSGBNTX3TgCPIIt9mM5Dfy/27G
geQRt2xNdBYue2CXsA5CLc9cr3GdK5uzZ+zywYZrnI7tjCwRQq5zoH+TIqtEIYW0
gwi52gVYM98UMH1s2fCd1oVXCnCexKUOe4br8uAo1e7BDxuazjM25V9ZHB/yY7qT
a6Pdj/HLT4yiPuesMWzyelJSbYMbMsFAjgmP/skzQaA/gXBC5MKMotH6dH9bx+FM
/6qGUkgnFBom9cPRjFSFqNnik6eIRv2rJJbOq3BJhfNpiUEra7nbc4RULfA6XkK6
/to8SnpBayjGA20//T1wqcJEPeJB8+MtYeey8m5r1F5jBFkmZH7Sk5QBDKgxO3Gl
4XBFXECxRjj4dH+Bg4Q84c1JQlr7zedhrmNg652YzzmkMQYPwmfbwA5NhnHpDfp3
5ZUKuUmgONBJ4mb9/astUAN7DfT++ePKote9kP6KJWNPyLfh8cx3LyOhgh5rM6wK
2V9MAOyvgrzolqOqPe2SNA5qihZlebP5fSUA/h22TIjyS/ByHAEJwpqwdHxFFhqE
hElQ2L/Kp2YmmKpfgeZB1VYX250XEZBEK3Vk2r2D2SWOGF22LaJiHymOtDPby1oa
Q160RSDQdWfYqlG5ljzvcw1vX0moAU1mh99pMar0THlVKk2YM1YW72yEtEtnKeAD
KivN0/0huYvoltaCyHFkmF7g7cjcdxO9q1htKDHGlI1A5HpLRUPOe/GhrS5SlIun
h1VCW4hviBV2IZ7p+EQNnKv1TbKc3V0dATH1g/2sLHJSESpyfA11hkgwrbV+kkuF
jn+OBOdY/DLYowqc3YXYDomjvv+eO72MpB59XQr7VWmiLTJExlvRAvkt7uq1i98/
4H7RbldimfCRTvwp0IXaR/Xk4Vs40ah7qp/I8NxmA9uDL0uONfluSOLJO4QKze6/
SiOw0bwIAiVkAABH2YvJUvT+KpajSTeVQO3VcxY7XAw=
`protect END_PROTECTED
