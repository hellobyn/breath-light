`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeIrux9pV+g4aAPWiQRg9LMbHfGDX7vXCBKyQvqYozI9HURseIecGvntyuJStk4s
+H1rPBuSeVVvPr9iKhOZZJPFKgVan3p6kG0FjT+mViTYd8QTE10leZLmVrUOAmH8
q3v/ueFptdck2lYaBw8p12TNQVP3SAHPExp9gX4DIcZsCgl2FP+28jlzVtLOq9dJ
HwMRSbnkUXwmvu6lxySSmEaVjXxyJuowTMwG+dSenMvRiPrKZel2rtCwj49jhyQT
VcnoTe78bNI6WL2u3/lv/Y3EBa+wus6lSjLaDemGCM2QADiwWyeaDfXhaMOc4ZeE
Yw5Bifat+nIfO7CBWDjVtceV5LLR8oabFOy0y8F5yvvBoJLqP9jwt9KmyGproEao
dCM2gPeRw2g7Yz3kvoX9nTOFIwlwWxmJ33oExYxUMguOqWnBqkI38Z3eBRLiB6JT
2QScud7TA+8njnGZTIdGrTO0sTz6mz+oltqrdtElfxKEhOj+5pnYRnJuFjCkIado
ifpEJtLsnMSRO0pHmy/d7bbGOHseOr4GCzEwqbYAEwyyJTfChz77nR7p0hRyVqVI
awT+iWjpkb2lDPI1+jT+naczQ64nCum6zJBvH8vWEbLg6lo9GRuuXJhuSQVSVrJw
ZTiBey7DKwxM/egbQYG+ESQ9i7NQb+w/PphucYVlYuWsRWcY9NjkueRaCZcctBix
n4Np4cDe8xdgqnd8A4qUhb3ohITw+BQ0ecmQMa9wm/HSTsdPTI4FahUNTIzpTOTd
0Aat4Lf1ErOM55ZEp1eYA3cyxk8O7hN96cHZNx5DGfuOhjlLdrgNHd7hZOBERwUr
rhayqh36uNC5HIAN2OPkTEaQZ78cTMXEDc5gzUk0+4ZppBK1hsEfereJ98dxgiyu
XpQ/MTaC5PhBTQjd2ASJQU5I2UZ8JLI6aMSPND+SXh7nDnysVCvO/cYrA9feIgkh
dfayYoFoDj3M57FdJbxI0EKucqOw3RFsKjQFfCf4tqjhBxGeoWTj6OLVH04kRmW+
S8IprlWDqlmLEj6cmjmqoDlorsH9kyUB6Tm6zdjugAOhp0uUjXegaQIEIBnSCzcV
hygT9p2N+P2f2Czx6dOezpa6p+Nj7R2FU0WrbZNuyUUrJlWsMj6Myo+NKDBdtDNS
vE1T1mA9WCj71eq9RnwE5Q8tuXxvDERWhZWy5EMfu2XqBafDDseZxmVHzH2a7oag
NniuTLXTnjYb3pHDSCeLUxFMqWSUdgO5KB2+Mywnf4Ndlsl3wlrgsTE7LE+iicGL
IyxSWMARyhL6FjuPxx1+FtdsVrBih1wNwoDjPQ2edOtNWPHdvMJvLHKsGTfX/6ro
sr0H18loj8GjvpPcSCsJ1wEPjfC9u7fRQ6ryy7VbFF/Iwodn9qFJsA6r8/n6ePe1
s3rnu6IkXj9Zqhp2YUhtRACFyRkrJEyVAddkxolexYFjQXkbxf+KizIajMVVIGW+
goqWxVU0Rz7F1ovY50HxzrPt5D5w4DRZnToKPV6VynFrTXBkpQ/pJ3NVUHVI69bO
NZpH6cqtyC6rPfXVvIfozK04s4VlIsfWlCMWgexClS5rTPxkAyAyaNRD7+XsCAA7
pATuvZV1zLYLmLoEuoNUmdnsWF/InaPaF37JYMnr6kxWTh13oRozBsU21RUdfw3Z
PAyIvouq8vk47f29uf0SX2cfi4HZhwGGaPLLD4aPoI64leTfCUlCX9q+irqiSreg
OQhp6QPTBYu8XCxHSPCs0vmDbu+RsBLQPPMgExaJbmauG/bEE9JF9ewHd9f3bIAh
gh1PJiggUiTtmj0tcoyZb0J2u1AzSmMUegnmWkOJHLwmh6wygyVb89oDRmaYldBW
wIDt4qZE9gmlfNHjLrqBLO7L1M6jyv/tum6b5J9VZwLXaax1hhw6Ds33L9EV+7Kl
CWle2ZsEfONlUGo60RbwWXVkZ0Lw/cNinV/NrRfNRstZBFYpJRa9c+pUZonFjJdi
yu4TV6/g0kDKcTfT29X+cv3cjVLhWNWB+gQCXR7J5Fy6i/h3Nw9bLCRTPosxrGTM
oSZ/lovSKCUO9hPC0NmNIc2xczpY6OzzZ88+646YfvqiBoLZ8cKaI71HsmyTrAow
nrR7CmaFYi2MeulvhHhBFFjVK3L/zHyN2Oe4OoCzxMnqEmvUsui7GtH3zQzDj4PT
rmtXhfY9HSpccHgguYm4iMD45w3wEjlEsybUAZPr1Le1cIMnGgauhbx58XVb0x9D
pq1s0jt8dAqw6XCiVWpY7pn7x7Hg/78aDYfmFsfwVDSE+Pky3wgnaiwNzVwpI7XA
9FRXMn682Tkjks+f/RhtUlkPXjQcNlW1rIRiVN0PmglRIaItyV802HdB8xd3JhXn
Cu1Z32CGaQxOd7LLbTHzWb8KVuGyHbkJjXN3RTSZ9jUlVA6Pv9FqkrXINk191sZh
nK7nuhkT1Aak02CwR8C3HB0oYyUOpFE0Ju/Wpb7JtH15VqCuEh4LN1FDCZ5yStYl
HOFkE0zEo5xr1A7gwj6ZJMxvdEmH5AlnBzXEoM/B85pCv3hqP+SrAGEMgZZbF3kM
znE8SfSMOqrDVs3Z5/8MfojF6uMhxVKaB6BlVupi0RQshIkW80Nm56gv+3FTUJ7D
Yft+vRLdqBH+Zue4wgAZ5ZyOuPtIwGzbpE41qrqi/okVjsW6o2n/kutAfkLCqxxU
aujtJi8FaA4ytDLr2LVqt7U20cbfcDKUU5WDK1M6XUwzcjGRIzsi33pKAIzSR3Jv
O7wBW5E7ijzMruxQeMud9QZ++ujYZZ1LL/lyp1NTRF5/NKGWZTz6HKG+ctAtudiP
emjRKnXpvGeg09sdjBBKYZpCayWL9RuBovNhx+4pQNTTrKRr1jcgeEthHL2kBjdd
lCAQkCOtpnihvBT1cuQpiOLXaDtUi59zIhAcilkbXUHSoNjuwfYA5k0NvBcvOvOD
Zd0XYyV0ajT1iOO2vHfp8zfJgaXiWULFbdUdxQhmHJQ1Qs8n04sd0vrBCzLzoQBu
KJJq4a7pOXGiTrcV+JyTe30MCsJiI9o3uKKTSxddkdAAFwrqr+nMxKxUSqXV/58p
itvt2NrkcFaNAlFzxsXNSmyobDFO1EtoYr5rr3ToR5K/HlMdcydgHgjgobvggHmO
Zc/vr2B6XdSl0ASb6q/E6dEFzLCOc17Wh5vcvLk05qg6D3ovoCY41r/2XHA7Huh7
aIWpkrwa804Pg8OBXlKmK4cWAff9JiIETEDoCEyBhsOvIxgNuV/tgJCzihCqK3PV
kF/3YYUE+YCFXaLZUH0c6PWU1AYZh5GS3Hfq7n1sLYoBr0sQNQGHE+hqWt3Wky3V
R4IXJGPQDn8XB8kB30BjjZyE77PTm+lOm0yGkWAjO6Kdrt5b0fpWF+1y+kdtanU1
KA67EGW50QDsOxUaFhl+oKvf2Nxedu+H0zkq1p9knbpXdwKxbaOIRifFhN18EZKj
LJaGT4S7qA94ytui3dn8acrEbj0UHEyrtQ5h5wyeUBiaGMT30eSGv+Jcuf094WN3
FqGX7niJO338qdnHOT8FJgV0d2TAZltOU+Csw881PcTHqWXl47f7/A4uLJqLeid8
LGdQMFwOfKrVkETO6eDVTgVv2mEIazv+NDT2PISjFS4Du/buNVlFL5FdeSfvDyr+
WxLnHkABszprImypB8R4diRUyTukM/eJw9Iimd3xbIXto0Dr9ljuojIAzdIi0uOh
iDJbR8WVuUn2RuSe0jC49O4Jp1e7w81VrohAYU09BWKIc8SUTl1txe0zOidy4dj6
cJElufZQ8D4SZ42QD/9RdAkeIHHYphGHHReEGXjQ9SONG8QE+j6igYpLQrzyEPfx
xn23iMVfKF1T1DndK825pCjyU2lwgUaLPM89uVYdBIFDto7/EHe/LD+HvqkcX8PK
+7GwBBHWTRtBIpJd5huDylw8SRqPRcD2T/SJJCd1/SYreUrz89XUOouTKrc8Q6k0
VD/Oh/Y7+60B4nqkrlq24je5jtpnmbt0jxBh/47lgoBThfmn6a0mxE2DYb2wHlNL
/fWoHc8BHbbLr64w8K2J+To9csIfRzooaowSme6+oJVji90eObDLQmAJfJ3RHgrs
Zsc4UqliPEwFRNO5gBxGQ2CwPrW2c2l1vpwuIk+HxUQ6oJvD/8uR+snenqxyHiRR
Kge4//KBiNEpQ/R9n45bdrAUh5riWdlXIJqVjwlF6GMaRuyf0StJs1Urx/pit5Rb
w2K0SF1g2H5XmoJrQTubXqYWuopH8RMOl8i0yJ4H2f5ZrJwqB8C3fTqesFNhlR5Z
BNqqnqlCKP7+Xox/n1YBbIWG4edLWr9eInfP4VrFaadcj7NcTyI49yPH7bRgIxQe
e5Tqn8wMojC0bAcE+JAUWhvAhboXEC7Z6dhZKm38OTlRvBQF6NVwsRmTbFZE7a+M
C29SMysNw5Se4sqO5NNSv8YRD5qIGmvGfJG41pXT8HJcMPVTgWurg45ID8BjPNEJ
BVkMZuS7z7FTt6u0X27J49kfFdBHI6IX3tCgu2IVpHolVBH5etVJV844S98Lo2Zz
iXfTqviUwUSgSNpthunoBWwKRBISiMsXqlefU6QJBZYjEyGGYPX2PDIoSJ5omvGL
CJVPO3x5NCOevFpySWX2tLFROrKTCWg3yc9F8xwGHtuDoFq2AsuaLXu9rcZNSUuW
WROOIuug8//VHKhI7kNzHdMgMEX4vO0B4GT4ZDoUjMG2ZSHNaGDQtTqAsOJHO7pL
hVhKmucL9I1hscJPXTWGimUugbQbbvMXRsBssw5QZUKD4anKOLTU52p4Sf4emH6F
UtEQk2bbHU+pL1G6rsxGQUkKlwFxVmHTlbTXkKDGqSDafsJcsFvSJpVx+dsluZm/
lwspNlHi9gKXYW/iJDgICfPfyS+5ElMxREe9nT4BeRf9Ey75hwoeWSVVmDIxpZif
SQAL3d8+tFJKDeZg8Eeni/xR98N0jzYuVjporHayefSR7xlg3l+wB8JkdoMBAs2J
Ur+T7iD69APrpYwixnmb7s2M9ujxUklT2Dqwh0W0qw0DI5w25XIHi6NHrTVBO9u4
MY+cuw8qXGwSVF2TwV9BXGnCNt1T7L4znId8Rw2pwBLagTpGS4CIOH6bzcLhU15O
WzYD2YNGglvXSB79HK1aQ0y8gAI4kUFPhsqGjsv4omMN2WTkXAzkyLoxduWtfKx9
8szVhloeT+9ePAEsPppKEwWQDluDucMmp5Mk14lH5AM3lnQBuG+bqW5p0FDWlW9+
WRYwoDBDN/204wogL/16ZAvU+msBWE7rR22l8axvseF8CaSNR5ZUyhhOeqbJ360b
JVAHrFlZO/srmanMaqv8wj/MDO6KSFe80pfv7qRrqYVWDFWL4lCZ1ll9haaEThW6
9tRdgojW8qSeixXXugIDHVTFFShEYNLvE4aPml2mq8Tpl3HXa25zUkHw0loxlzHV
xpQ+tINY5ph2v+N4kAZANLf6Bh8zjQ/6XBItdd2afFxGZ2p9W4K0sUykQzWcFQ5x
apBkJc7byPrqPuFXrNq+YOc2W6Ws1TC3pLeOSwN0HepuPMAz8TaTn+VjaSw1Xgin
6Pa08wOxZlChBEP6z0JWk5AI1/WA2fkd2Z15rdUtMXOHsowBl5z9e74N7FVbVMZf
K/QvwBPEAJQSbRjPki0PJOjbmfBa/x5etn31IttaIKvvtos86tAAiI/llaLj5C2k
gXq73OWfT7Hd6HLGoNpbYsO8GQ+NlckJRhrb7u0Pp0jhqhoViVw1G+K64Hx5CIKA
OuEuYiuJ6uoT8HIoxnOisdSWIHh6Lgc4Wrgx9LVPZSz2cwbvdt/2avWKNrnAxUjN
SrqJygzn9ccTtabRIsHq0/F/fMO8FKhIlMzAaWY576DVAvMbt/C4dckjBCfnubWm
OOHY0Xht/GXsHJJ7wmgjorSzxV1CKXqwpPdBG88DZqtG9Je+75ILAgW2RBTOefIv
kKhisfZuuOIXEBx6auGZfSZrXu18yQ8zt5xHIzY6qgdOkkG70kdZn5G9/rLm7Yxj
fN/E3Qrss/ayDCXxHqEFUFz2deE80pgjArCIMMakC7PtGOYRjV4sE/aXRlHTwPC0
gB0/dDQe03xeATMSWdAsuS9y6q9p2sViFcGo1npm145LhQBJMX+iMsvF/VQC4h/p
0hIe49h8BvKSGx3bX3BS3sQYGeK7uFBZZZk0ataXwnDH8P5k0DEAb3hQNzwl8Op7
v8HZ4TjQvBci+t7Q8jbKtdyPuMpSQPlWFOhmscrNeCAbi7AbjaChIiRVy1Gr7VLg
+kqwzmtF5Rq0w7SE9vRWJnvRPC0T+lfXwpLSxy6eZbQ8S1+uNzDXYp6MC2WGgZPH
Bvf8wEzD+iePvcHexMTqeKgR51UxAxpBeMpdmlqOOsq3wsMxPwMs/SAGSc+f23JF
jCmwqEmoho/SdIHMXaRJ7SHKO0hglnq9h938tHcgmFAPaOLB76iG43YdaM8VcMHM
J8NrhBoPN3utvhVVJwmHR++P9SSIM3xNgOdiwyw441KHS/SAT3eujuv0KrJ2gkum
nwiDfoGEbK8ULQDashM1qQuW35BTF2z07ivzzYoeCLkPRFRALSm1Er967SshunxO
q41mK3wGrPNw0/xTzKZyJj4+z0QlmWqZQHyvoOtAhvsL/yrBYtTEuGFdOgxbeND3
s6ntywn6BH7GZU27EIpSW4abEB7QMf02NnR8v1VdyU22k0Ct7qyaasZt8w+sB+fI
kPah8YiB2rfd0mGutmYSWQ9UuA5vXR5t/J8E5mxpf5ygD0TWWkPnT2VKOrvVfMYZ
kAXwwwdhJwjNOsSmiz9nCA27HPnI86hdmEYUSOuzrnEoikohQBojmRnttZuGqaEy
TbZ3w0qEMOLBTSQEJ0r5TZSlh10Bhu6cI6si8uRvNDbUnuxAaLgWhBCi5ozhwfa/
XUBlRtU9cPx+8+tGPKFQB9P/0NMLq6U6IkR4uuS4kTw4X7sgsl5IUh0hGFp0LSV+
Gis6BA9ARWZbuCfaz6i/1zelW8U0CVHyqCgTHgM36LL6MpnNeoRtid0CLZsNTL//
y/YiXZmhkwduCjWsOJQJXg3OOE6fz/XERnmdlcSqSXlqDMHLsU3mP30g79JkZyaD
9iRMReoOJmZuTovj5pbBtf/MiNNyaw6pTNQdZwc/DRYPmEhCVWA/GfDCeT4ztPGO
HEeoeiOm1xf8GqESYOinzuNqFzGS1fn6bykzCPqsJxm4aAmiC4hUQ6TKfahx3o9Z
+HOeRHiJL+PrkLiY1JVpUAYf5zv/NMx8s0EifAZioLySJFKMgnzPHVaVjAOchr8d
eXjES9jP5kkJQ6DXgTu0waJosqU4vAbHxzVnO+ZQT+e8NPQ67DhCMt+Mi4jRX2lV
n/s/EZkueASqw8qKLBq9MpSaKFT7yvS9F0dAbcApfnrN2pb4cNhVWGHkhQdtYjD3
muQHV9SwF5oqCtbPAJXkFwK4B8YizIWJfn08Yq+P0FHRkTACKQzWblPf7Qw9eFkW
xv6DSXEfbqnBeVWQ9IJW0BDe/a6/JHjuNM1n3NqJOZu/CvOmGIGdzSvzvTNpUacJ
DBuyKXG0Hf4JhGFd1q6dtgQmwArmQWDdgaHmigjypMRHT9pc3S3+wY7+o/T16Y1N
dVFMREc7EsJft3bU1ZQu29S4EXumqW/sWQWTj35fWkEbH3qqFw+WN0LGLZSVHBEj
y7lYhOzcVwkd4OyIG5Il/FxHZ8o0SPLikE9lQUuqbpoy3cpUj1wL8HoOh4h/moBU
a8E4iv+m2uvQXF69LoWBTktDtG4qRyq1hqmdHUQwKgdOG0TVpX3qES2JNh35hjGK
xNK2hQTtG5oP5q/ehAyajQUJ4kyBDKvgqyH5UXcMx4ixM+wsDjaGcaJcZbvbPrpo
PaTXGFsyVZtB8u/AR7anQG9KzqG1H+BA8Cr5AM7kwAsoulVHbfSddBPv+Ena1F80
T/YIxXEnr/kJJiZTJMa4+N4scbdzKRgfxtDhyoGDAoiV2CAljZyiLxXReP+LX8dL
V+PKUxBadla0nD6PkUgf8qdk4cCJb2SDMEyCm49GLPRcVt2ntGGWIQ4JXLQctr4c
Mt3Bx9PMxjZhOSddQv0R619PGGGYIJaTrCh2C3FpggGek6JkswsLXKDZZDG2SSSP
4k0JKsHcQjZcZ5CNMdCduEVEl234hUSpkssZbZy+n0U3BF4txno7Zz6dVG+qYqHA
9NQYu2J7WqSZqHPANHE+jyE1XXX3J5j+g7jcN81OnKuyFSj3ZQwahLo1eefW31Vz
RFkW2ahoiAVMnIzjt69QkYRIZNRF4J+4UmvYgDI8LWPkUgthus2cecNTmm7kv7Mu
U4oAi6O72HDigliyvad08+NXIgBX3nPHrZ6DoyEMxygrXaPJOhMofENQcuQNTzkz
1YfYrjt6AVE1ThgLN5JushOwc5ilPDLbsNrMH5vkM7RudPn4sjb8vhIpb+OAsSMf
Shl0Qk3FOszts2Q7iRjZv/Hfz09ZFiE25OZL2GCOgmcxECNoe73E7b71R4vNZ+6k
/wxAZptZo+CVzAiNs4WVy6C2ViAO6eNHLFds1HbYT4de6rdFT7Bw/dvy6Jrb6hYt
n9FgXgKIKqH2wEiBBTsNNiUFWkSJ5STSM5nyKXHmXvq7xXi89Km3RynoY/3SeShI
4+bj0EVBMjEG/ZQR3TeRwoL6NtPHC6ztzx0faUdkdFkGjhVd2XAxbepiKXw56s3/
s+0goqLEwVeZPG9pXIS8z0zxM26bi1N7UGZpxHO00QX7/B+8I1fdj1QDoQE4X0xF
oXNojzqFYfJkvh3b3hXC51YCJhs27VsJkNMEJig3xLGc76h6Np9BrL4rWbeV20DX
q4yonfGMyBYPMaFQV5ZkzNjxYTx4zLdnozfU68L87ZO1A8Mssei6u29JNegtNkN+
vkrmfbPE/KITKagl7G++v4+75qlLNl9o3XQ2sFmlyEk6+H/nvYEIxKGZXNelQOdg
l2+jlYFOWAAzwmHua1IQJk4x/7R4Suf9hsbLTsjYoKDD+0YQFnIstaNRToTHQrA1
7k3PnEHI9WApL6e3a/g9JuAdw6woA8T+Ud3Uv4HOJJ7pQk3EEBsY8lHg0XmHKfhI
stw3Svov70zmnb7n6gLAXJXh37VVwhrRWQ77HGsLT37WYPZqLP46MzUdwf0CXqis
zryativ9D0bcL13P591jYZQGTsoRWuqS+1GP5HM2XGlKPGnWP1rcGPa0IkpyVJPF
+ZGXch62AjkWASsR8oaF4y5zc08sfTeHnsflRnm3FVBwgFXnTvnZPkhu2MhlkeWx
H5Jb7lV1e6t18RIeztdiLSmNR3G5AxN48kCN6BuXc8nt3f27NqqpX10ZMukLqErT
4wYWlBHZYnYZg7atTEWtCudZs2ICQOsZyZ4Q841Ml33S7zL1Y5gJyyRDnip2NXPi
ZeYIz/CzUF9Y2Q+NU11ubG+1cCi1Y0PdHAeuY4J/gB0/znN7l2CzSJ1K+v+ALD7H
B/0mq8ZmvK1VWnNSzE6/7QqNh7cDUdCCcIhVQ5kGcaj2XGlOcA3smKioHmisU2Vg
NUzRYoTx+dKTI7BpwN38ppkzOLoI6XHW/bHkQFuLKaiAeuFn70j0ZXW7L1OXwix3
4aK5EqAF1fSDDjF12FoE0CPyPgu8aRPj6rYIqKTsCqowSnabOJa5oIrZzbInIJW+
Jy13ShgLneDmauhpdvcoLty37nxVluLbVPHZ64TpuRtMLlRSKdTH7QxmQhURieNK
ayxGYFUJkYk2HSrasi0aPkZ7G7Wv7rha/IAjBfMJn/WjY6WMDgFwKT2vcSr63LI7
ND1BLF/v53p0AikEK5ufrH+KjqFZpdo66OGVF8DDK5AHQtjAGgeEJAZhSJbF15iJ
ASvKnw+10Nk02CWtDusZGUk+f++VZbTArNhdLvho5fsB658KsF9d6dQcF9WN9Guz
8fT8dOdeYXMEJFuTJIyVTlPw/qYOT7HQ7rVyuh6aVPsa9Y6sdAowmw3AJxC4NmdT
+EN79TZOEkqqQ7BPeWsR6YytyXKzo1tVhE4hrbcUHOeOqjNnxR3xQ/bgE+sRgusT
xAn5EGkudqbg1n53JRDDAla4ok/l4wpwkvW8/vF0Uq5474AtXOGCBmlfvR+LwuZt
dtD/rfpoSzE7M0mx2khJQyMXxDj0PVHekYnaZAWBqBRrp5bgmV1rhn1gPYpZqd55
+1jU7xnRMXFra/X9Y3uN8ONfBOPu1U4hTvoLuGO3cUCklEKO4hJjCqpYvGZ4b9ze
rHOSGgsGy3Nj3Euv94VdMnnmO1N8QaPSB0FJQruGfWtegvzTNGugQnXuM50Sb8rP
/fYNs8EpPY8EvyO4IEOkT9vs+zy2/GIw39GFVHvlICssy603ce35IOkW9mgqnhG4
dq7E69kytqeU5a+Be7fOzjoBSHTvMxxI3z2YF6yQuxUalH7DAC8H6BTgC+dhCsnX
boeSyBav8I3RvoShrFpzsoLp9meHcpBBxhTkIkdbsnx34XyMSjW3g6qdogxpniz3
aJYad9MHi8j6L4ovGaZdxoc9hJqGQ9hPuXok/XfIE7j9Yz/GKSqmVHcIVV3LjbXt
dj2A+firpoCdKH6CxvqHfz4TcYA7l8GwTas+ZkwjvMU+VeAcziXQm6FafuUgHlA8
sd02MZMRjaldyUKBdNPMlCi1T9SaIuomC6heo5yBD6KyNEo1TctOKoZ9H+V9KJr6
JDuiFTJpZa94Aza5PqUnKQkXu9WME+q3SgwDoTMt6HwmF9WxvwFthAh/eoUuwGNW
zc91tyj0zO60+xfyK8236MJmhynJTg339ghLGx2bmIZQpVOUtjCaA1whydxqblz3
qZHCTSUBF1dy8fTFdFGzPDIKewUgEaeLUiHtVviDDR3tyaKgI87osQ0RpGpIW/Cp
WzHQciDhjQoEnm0zBM8f9n4Xafhj/BPSHCtKpk38nGrYHcVrcHxt/fWpWEVNuFnZ
NbLOV6J+uLtK7GEQ+t2p25Km2vEoU6UUompir30lm2h+AfWw0H+gccC92vaSgpXL
reRjkyqjKIAq8cnVn96HKruoqzUmbIWrFFz/vwqEW3j5p0+poQG2ihugwSpdlYs+
bj1GbGYUstIf8ji3Wfm7DOqlGyz7GkO6rf1LhpbbzSuloHDlGgFgmLp7fg/mrB+Y
A0EgDYRIXb6qVP19kW2VpCIGO/MGtlt1Z75jMYC4bQIH3uI7FI4p2wUgHg20NJy4
cMPplupeEq/JVng9Ek8lrHiHLQOD4aNXkFgJlgFNhfYXKMeO2e/bp50203p0pHFd
4cudTtQds59VJJGCJUYh6yWn/tvv+94hQiWqDf77teAoOpEbqRAi/UXh1a1mT/jE
f3IWkyKkUZCBirV45SgwSpW76r9C2CVgQV6XMcX/xGwuCGbkQ6YQm4D3tvya3iki
X0sLgmFkEJC1ssLIo3jmIh29sXHsRT1gNMci+XFOA2dCHKf/NwoJQKNrS3BSGNr9
rWFEJo6z/hN3/7hkFR19Id269S+VEz+pBrA+XeOJb9bMCYyxoG6U4SyuYocPmaFs
DzWwndQ9pXXzMJB5B8lFEO8KwyFkWVogXsIy2vy0rpnx+BCLJj6wxpYdUsInWHrm
BpNQfDCJR7wUQLamLI3GP7GDDH9ihT1WmCaSQ0QI//R/4MjeRdzA7zjKIwZTkrzQ
fofTXF1V1FE3eWQKG8/TGGyfPGuUiBTyCoEpHF8j83c7PPvQyqjLy15XFBn/8FmC
NAJyc4yw8twOPXpXU+VUDiFQQmTgGCnhoFbZUuRkYJO9LjkPovqvRFDoUxf/axe1
NiqhxNDX7tLcXDhlsKhEjjACzVAatEmMwQaSe+kjcQNwiCsDIRPr19stE734lWuF
/X6tV2uudk5LuANyPWMP6trmS9XCKwXSaR3Hq9Eny0vMSP1w6IK6i9ctyPfvRCmk
Q3nWYcP3STkPQZSBtML48xf09B1L3bxLFHnvuBeVfTYPEE+j+/yaLJ0OF5B+7eLm
e9XwZhq9jeWA2UVJuH8rW3cZxsTGbfT2OdE5UGcfNGChCTQTd9/b95UqKUUqMEkA
y+xVJ2NlRWv+j4Rt5AB2CfnjzvKBU1Er9Iv2ZgOlBQ/Boc9R1VWUNK7+XGq+sQLE
A9y93Na1xoHfy0DRA/yMDGUhYXHFwvCQMDhiQhmvELHgxGACYTQ0LOVm2Ikw395b
3EPiHmwAHzZLGokkmlPyOYA+ko1bxYhzsL81uIfjXogYFztEfKscIpWGC1+ZAtH5
VWwRbjg5tO74cotR443v8GxI+hKHc+J6exVOn6zkXRTX42ClDPy2ZORsGJBaKFsU
mCajXQc7r0+x00WgLAfuLSfs1Ehi3k2NzLsM5yfIuQXn8pTVb9xHmoCzYyoTNNVX
DRgCQZGL26hEagTsZm6D2QHIL96qHTargUKHNWdF++Sig3qpiLOX0KZQqTg/k1XB
M5sWqb7iIDFeTPLP6yRQqmUfq0E1JKogy1uL1kJ59ATGSqD18XtzDFN157QbKXvg
Ry31q90M2hmMIItitMOnlmeP70obR7F8ZXn3PQIQiUX58nrqoHuiuyOvxTZCissG
1AQmW1y4wS3iD30QUZhJMR014QwMhtQLYwJR6IhiRAsDvO9bRSfm/gVPh+pd36TS
D7EkJ9HnIolioES9WPsTDBpksaTHc7WUa43bMc84lfP7CdL7q/Pm/ElysuMobqLU
T15BPRlOIT6t06MFqXKTrwDovwByuQN2tdSLJGZptYE/jLuj2bZ+3CAptR1hkRPR
09XiISCSrN72aiDT5FDWSV4a/OvE75dufzHNl+iW3KVN3GqGC01pOTPc0quFzM5y
c2HPUL0GxVy6D+1cyC4/j9Z4CYyRy/DkAlI0laGf12+KqvSkQ9ZO0OaT597IWtKi
1YREIHERjfg9sI5tz+tke24tFoW92GAy3NkbXjNPJWmH/YK8MRopqcjXJKjbzTrI
h80eWon7B8YCM+3Hs9DYCEY9Pqs3XRB4hAGIUTMFpKyD3m9RsPxRyEGL4X4BINdn
upcPG0qF1+6FOeSOn6l801tzOfoEqj4QOJtOj4cBMhMZnVzwLzPjQ/rB5MrCO3Xy
lLB7X11osEnLoJJVJF1KjFwcwTa7mNXe6TpiCV/bmSUlmoaJodDk5d2QtziToH1F
EhFdkfnkMY0t1ZXxnjJz3ce2kI0rUVdmXR/et/BU/mTw4AE6p882An81s+T5Iasd
vnRKm+UW7vl/+Vp+59j1DmsWfl2U4mM90lIv2uah3X180teTFKiw8Q4kByeYobq0
5i8UE5wMhXmllNNSFbmXYHMA29E5EwnjjjSiSXLxyZB5o1u761+4je4sWfpUVRh6
DZdQne+j36HVDZKQPJBvZO1M/gPdC4FiRIujf9na8dAoilyNPA2sfwlHHr8U5orH
+gRi2M9SZmQutKAPC/wW9vRRGwW93bgDtooc+8U60Z7Lv5aXlStnMLZIC/LTwr5l
Tsn67CeCfIQdzYCrIie9ZIY/998vKRj2a8XOj5JiAovN54eOKhXLHJ9jBSjSBBh9
Yg9QDOrG6kDwGPtJSEPPdkRr2VmQ44rW/lsaIQcLG6JaUEkqNSWbGzi4f6e+ktyF
gW5bXCfdlrrQLDGfISwcas8toI1nB+SzqMcRZVT3WL4rrvIkZUd3x9UZdzU/ghCS
gPRuXgIglnDlR7SMMHfhh8Ym+G+DkYJNuhYmKT+psOd6Y1BvfrqnsWx/9fvbPY7L
T/bBr34gOMReR26sg10rG2Ke/Kml4izQXycM2n0hWnhZrt8mvBbsW7A3ppnK0Ys0
lbczKKf4JemWu1JTgN4e4KBkT/n6xkNLCGx4n5qYlgBGK4VKNbIw0QC6g0Mc38m8
Fmh6E8d8LfO5zFDj7AhRCKpulNYx0fWdCy+XnQWpC+5OYwRn4VUW9Ffa7dDOZuRH
cZD4ZgCKu9W4VJY9WR6N4K8Ok3KIhLKZkH1hwx8YH3vt2g2VFkPgdZ0U24qmTyFs
5TSUf+B2lWArDTzs0cNd7P9woNfGYqLbJo/PyZOGmnbHEJRof4ac4EAu2VoBO1Mc
CQ53U27ec0uN8S+vvQcHz2mEGLYaCXe/VyouT/xyyaBcH7AhodkqEBOup1cdBhAG
Wt1rvoCjGjOAnXActdV+tUM6uXqshiPl6LIDeNBKK+mcmdvuuLpRiRtmlRb6F3ly
D09quSXSaqbHxxuZuM4SnSKTbVHneYRw7PUDOMmw29hkaSPXOE099l3n4hOgvMlU
FJs5nc4yO5MOrKE4fyuuQ+d+/57Bbt/2xTt4Ozlpo3074P0MWhZTNBiLGX24fhTg
ybGnfnwzRm/Z1CW6pZ7wtmWiFFAr2G2bdB3CYN0vffm4qgIGXUScuyCDp9mh7pWu
cqLBUCOhrqo44SmOfrAxO0NDLwDzu/jeewo6j2E88Rv28D0r3iCZ3Kekf2y5m+B/
MACazyUxc0aWRoa5VCJthFOXNAI+S9VRIAxLpyz/GuCiiD/CBBu7pVL0n/YQuTRH
8qT04oXHcqk8lUU1yEfjuIxZ3ffP04vjDaL4QBBjb1C/hj2evct9wUpsYPe/bQur
KaDzN4WZOBS+Fsoa5uHpu7utN/pL+8/ZQ9w5RTCfCZPirG2NhguwwuGWnpA/IXiS
EmYYxr8jDr+AMHU3/TPJFdjPhZBQwiC0B1uYY82c+MQb+DEyd0xzibFJIs6Dy1mR
XwKSeya1u4Im5aK78CejVJlV91aMhpRy+OhN61nuSb0AL3MrHko3lIss2j7WClwd
QoZ1hL6Y5vdu8o9R/J3IGFD26tobD6FOjrsxU+zjgXvBS3G2vwQ0UF6G/jzsdD+2
Up4RzpinBkR5G5gS4NqETR55afpqhen4kJA2RcGOL1VfQ+HCa215D4OaiPy+0gb0
n07irLuveaPdZioziRGI0OlwOechTw4dMZXDDEjx0I5D0O7ToB90os5xm0fz396V
WpY1V4J3SyOSxeg3tb7oKi34XKFHAJ1Z210vo07Hy4gfockFPfJLSFlbYGmkpNuK
vFwV2jRCq60qww++1Z1U6rIYd8Kz1hiYj/XZzZKrUtWwOCfUmw9Jwy6TcVqx1jgc
R4EHGlkv7dN2jKt5ZjJCh6SBrxbiXf9DQSgViIRMIuRAUKTe2Yld9d/NpI+32i4n
r8bABqR3l6sVMspB8wbp7nxESUOQLtr/AQunwHBMN1pGMw8ZWlmks2UjGQHrdevV
jtUrfZTPjOxW+2JMC7UhuJFhUIF4PqoBev0L+m/tiCoB5XULhMhK+hqJ7Guhi49n
zespY4DYBY2PRc40PaLe+YS1DRmKxOKNu78WfWhcHmCKU0ek4TrSuuHdApPFMUjv
dbMYmqGKf378ejuZndAQ1OosY6NoIrsy/lJULmQzgr7K/CcvsKG2x8xuBNBxdq6D
x5NtyT/E48eBp7Jv8FE0RN9f7GgyPNrngqDwfz/Cf6oy6M8Thqk84pob837E7wTv
Bu8+E+fhHo8lCXPcKCwBx6tc1UVeW94E5I7PUwrUMtJbyvGA9yWLdsyBwxsEs0CL
UUC3qnQwHE3FKsY36wgOT5vP+P3uNNeuIKh7nxO2NemmG2RLnNFFyJXjtrUPh11H
oULu4Uh5Lh4x5y1sYBijmA2OUP9WPAZeCdEi9PRmrrKGE/YnrsLJId3EVVk+5MOi
fkQFFGphqTp0egmCelTbWOdLmxVpN8OxEfnKkil+mgJZQbQKzUgmYxunw9ccK9d9
/nrM9KeShU68SQTqAo1QlEHIv3NmkT19AqfJlaCMCPihnLFFH6hJyCa9SzJO5Y2+
ALzPdA8u580ItxocTk76BK55Sm8w1fIizMkgcDbHgi/MSlzjuBz44DVtfKwXqOaZ
SK2t/Om/QqLuBNdwA345neOJF/RsTc1RNZvS//fRO2JXhUX8zd2jpWro8jDll+8E
SYcgFL9kZrTawgtpSItUm6yYLkxnTRbJ3diWUumqcDdggY5f50YwvRTVecdzRdkg
9cZoEWEEXTZnw+8NOdU/s0emIJusxwo9d4xVR4xVzKEI0MAxQEP49cx9DvuguCvn
DVaNgBbkI170Iga+e9IAmFWUon+Un62teqBea9ZOzLukiFYmGRnrJDiqE1d+Y5pt
y3KytkmijBpLBJHX50zDDnZk8AOj6jRVEcO6k4STxzJfKlEs6p8Ce18Ag3fjJ1JT
H/M78gNqA7o3gu+71Lz93HBUu/cN5ZRrJE/h0fltLH4LGnjKBY/y8nv2WcGP1v/e
MQk2bMwjOtlRuWoI3VNixixLe3+5gNgRtTY1PZ5rkcyuDkpUPRs2T6DUtRvxwQH/
kGq+g/tZbxRBUP119g8yPW8VABaQl0GDIER4j+vkoNO5RXkUdW2MrSphWpBhQaUD
zrc4oreULcFGG+I8aCqHHazITyafGR+1m54+5Q1VqJGeAWd7HQ2uHx4ReoGAeMbY
jzfeJxHec/MAAjb8FoNC8DagqHL1VN2hAL9lRy9A2Kk43hv7qW1MeV7/KKgZjb/E
MJ914XHxascG20qOoV6/OMUIGEGCP45bR+718ZMsHISjK/3n5Ns24CmcrKqTlorY
er36yTnuffAPaTqXLToy0rXPqGEXUdd6WZS9VVvtM/w2EqQoW1+K6v/a3ugzUMkX
1g1oDYdVIv+AZZltCmJyShI90cGCr0uFXFuJsKQiqI66D6U0N5G/0Ov6vKSQfkhE
zMA6FYTCsPtriX96dnC8Tp6COUCGCTcgTWoJgsE6c4raVK354a7FVTgYBVfwkuvV
h+0kFF+nOjhDtS5N4urLviz3naIrfQxRu7FsgoSAbE0XoArQivBe01cjxxoQEPzl
khs8jZs61PqWRXKcN5mzjOgS6kpkPAzBpSJuo8JYKE0F9B43JLcDRWPiPsX/c4hY
vFf3ntIsuEI+XqX4pdX0xXgLzBM5Wn73UCzuVZxqHmQ6GK9atgkjOoFORtx674Sl
nwHkeyGWVGpWczRm4f+YLcXBgSvK0yZykvzqflyVbLzETZgC/kkLh0sbqvB9nsRN
ffvvz+uXycVGZtMzmYD7KpwjmkcUJd+y2+R3VmieIJTJ0ogiNpiiIi6nbEk+3EeX
G5MO6vkL+f5y3J3lQvgO7MctKAV67rrcaQDOYv45NG75pKj92uZmQHVr1/kPlwQL
5YqRHhQ5J54SKvhgHXnC0sTFR3FKHtJ+pCrMThr4NKCL/bOV6TQ6JhO9bl2vOHa9
TQFvzeZBagAk1Lu52r96FskJ7f3ro2AmkbGwssVW3cu0g4xm1n+XEtoK+Rk97Qlv
tr8O5PI0vzW2jnKsW7939uTHZ7rnYl/dlVpdKyTN/IhiJxYtWCCw8x8ltzPnDBpt
RxoijQmNP1yzS3yWdgDwPJ5YY0zjbfEc7ipR1Eh+wTWhBgeNNIUi/XiQaLAfSWZ7
D8K4n9tibtGxQF8kzHmho8C12oxLLMkN44Qizpv1sSGxcCujtESi1OSyLgy5WRxU
HMIQJ+Z/sdFebDq/aNmtGG77mMnLmUnE94r49XAJhET5pbJ5aZ03HloGsXRreyQf
8kt0bzBsKa52tVd+hdGnCpmgq8Tqc7r19eNfg7f+sWyL3UQY4q7Mb0V1YIrwKqlZ
o59jPlqsFF4PKGGu5fOpvpYGOCuf/57NTQXfgwmjwXd5T0qS/D+6d9gEbG2dyLbR
31XwrnAm5KPQH35/DfLJFOh+4xwyVN/4yHN+nWdbNRF4ah+kI5XT6EIr5/Jc9xrb
XOVKOo6FAjlEfsoUd67VRjO0Bl38Oh+6YZc2x3skyhiqJWCki8HulF9S6xLSEiEx
w55fgJoVIWpl8XTHRc4iSEJneTgVrcp2a6Xs/sROgq0nc/jnmIg6pptrC51x0B25
EV3Jxl1A2igeI0vtZlE41JDobmUuVOu0VvKQ6uNgyN0sLOT7rrGj58uMJOCNH0tz
sDkRDbAT+icEeEuuhnbeQ1qO/W8nZHgVINE87dIBZfdlerSdasmd3B2Qu9PqjJpv
mQ7+QCUfEg1CkqyVT/ahZ6xmbcGgs6dzXUeJ0N/jMJN6tHaW/1/KETvDDKBN5fJX
/y8PFBVl5FdHZiYJR/7SzotIkzG8aw/wk+YV2jPBuUg2RJ/ZeThQ93fR0RvL+wzG
kloRn8YnkM0P9vUq5r8fYZ/EMZmzx6GSHG1H+Gg8b+kfS29aD7IGPX3KXrqFkULb
Or1tyKcsdor+3+PzYp1OUo1GXq4eupwOM60Kkur7Zf7gfi90XphOzdFX1LRUAOHb
tQFS64KYG0q5hayvu1xxbdmaQqEydUaTE7b0O3zY422qXjOn3IVVYDH0ZMsZOCMC
dl/PzIuwae8vLm398hC5YI1HKjC1LeiHD+gDkNxZHFel6vPfW5pA2YJwfkjdGn5P
+gjQFtsezaPwzIUDJEvF7U6hW8krlIS2P1c0FC+xnbfidpxtmbmyjXXdW7VwGVni
c931LY+hAeI3fgZDYzJtL37iixOAY/Irl5JP8U1Dm05Vjj9K6AFgPXSm3l9dC6Sn
vHRoxCA1OEKNiNt3Vy7J6Cdf+96JDikl5N//R8Q6PbmgQ76bOrp11kYcALU/68dT
2gj0lhKJyjwsbKL+kib486M1k2sppV7qoF24DL9+l8RdqWKTJ5UpykO+26elHuAV
ZQ8EsqcTGDWA9vfS4bgVG4xmsGVIjz2ij+niC4I7jjP5COwLq+20SEJiUlCBmEAu
uPGXMIj9y9myyWKG+++BfHVyCCwWsvTKntNbgxS20SqKWIiEgYtQsDLlkTRW8LCm
/fbAu5l4beTracNWSZ5Pmhe5YLdOY2f+ykmm0yJxsfzX272CIWS+ftpb0SfbUdz2
HvD2MGLQfYO3TaK705lTsSf17i8T7f1zkV6bLBI9YabyB9nQI36EFVhG2uLttDiL
sNTbWT25nd24Bbj5/PprsidMd5DLGMJLhHs8d31r6LuSXusXLWw+WRGQGQcILrLU
zetsHrVEGW1edtiaQ1gzIl3D28aJxt/FNb7kiOpgPCyGIptQlybxNaguleGKan5/
MyQZeewWe1B0sgFgLuV/xOSJzKDmzezvSPp2ZRLMM7LRxjrw7sLnVlUyZfnVIMwQ
RHyD/KytBgfvjicG2j2CPTVcLnOLXS8R06goBnnLdThYU4nC7MZOSGXdI9tHnwVd
zfnyAE1n3mkjArMEtB40lGosEBI4lpgHLevCiySZjuWpic2xAatzWTPhVUuMjIAg
2SSQV5vwZu2UuQUxYDjnXh+slTeVjV1u+CtAS+ngNzh0JiIYeebedH4IZDs8CKro
8A0+qAi6SRs99MMPajnQQ64Ep/0q7AeIOW6ZYMljq2ghIQkJBUr9K+zkUGESTZm2
GjJVEwmY0u+IOTkAQWW+C7TSXCRXLZMnCvOUj8N2BSiaVatJZOqrMl5eJiqqgX5h
TolTCBShIOxxUzJU3qpxMSvKQQtkMy9xMxYaq5q8iEDj6uKGgwqy0QoPxUoZLJiO
CPmp89COXUcSf8TXM8G7NJGyALjXGXNMn1o5eEeXP5dRjQMCBu/Kl2mCM6bOVwtv
mt69QyEen23LC2kNhKzf5/uv6haZeUUA8oV3gOV/lf6HZrhg5PBXHutM5rlTmD59
uKxt29pdQFkMd67rBnWksGTPttO7fLzh51ZWK40QAhi2KU27AjT6xZEytCly29MF
RiEC1veqKDuZA4AX47c5uTVW9TxSqLBpPCVOeT0sNOdSR5yUjQGOOGfESPU8DNto
e/kpJ21h1h9n8/uTMerklvNBESIhu+rJxyndDSrYvzdmQ+168efsx8kwsnVwIgu6
wBmLgWIVVSdGijhfvzHPfiiFbnMuNoHorYAdmdPacH8OaiuzexzKlxVKnNq8baP/
eeKl3lj2Ub77ps4YcW7pD37ZkhwSY4pGbWJpTiU1n+egG9wH2M0AXUz9kYT+KxOP
naneCo5crSEGt7lN7fB2tKthkKNzESxqIXofBHlvWf94pDECDCYahBHfXMMjJy4t
UvZal2lo9cc6J6pkHbwhJ0fuAw4CAWLpq3Kt4wIFiz44xJU2uQLAzwIFN1owFGLN
js990JPb9W/epQFFTrDFEYJ1BeubLPWuGp89VmaLxTwlwDY3/qKWoz/ERSjbb4Zp
Lm2QNtO+34rymXOEvv8i9C4wcF9tNBymu4Z9DASEFebMjIsUmeN/56N7Xfegue5Q
Pjv36mhGwQ6CZDorFTyE9xX7MCPuPgPJx6gi7l2+LgDROg6zzHtFB0LFqovXgTd9
rdzEU1dBEfscXFNU/A10VQgmZl8NB2gWjyqP+PLu8hx23V/7vJmqlAMrypLFG8eg
fWq839NdeN4tgLARSkOEhI9jz9ZThLyRpBPzN6Nb23GQyLGxlFqav+/Rfut31dyI
YzbUkPaMHsMlGkXrYqDvkduTU/zQNTwgcKbO2k03rBF/tpoMpTa+aFpsxI9EfxlN
n1+S+e6cGy7VPWqRS1dZL++criGDTi1BVzFz+2BrRq+1QJtv0BO+Zm70BpOhwHay
SYGQryCu2xDggWBg2bPghqF8icVPPqq8pgIog3ltRvpCDewkwdECpZt9bjK69yHg
f8TBqRgFG3Qjra8ZRoRlJnv1SlrnGVUTe2f8S+SSA7zrZM/SKR2QC4DfgpH6vSq2
vjngODThDgW3FYhsgT6w+flfsBQ37fVVFeYWVCC2I3wDBv0UHWvX8tHyaghjrz1v
j0N6h6c95I+Lf6wYidxn56ck1cm+fEIyeEltdKsDTB3k7HPmGmhonTrKrAAm8162
kMk3lLN+x6TIkTVPMtH6loJPJoJ958xLz8EcJ1GRbq6MnODqyYkApdw+Db7PiIhH
+tpd2dT2XK1mbSkFnrHQi31jCxLnhBFNxefWBz9uoSNrECxWUwQAkw8TL5etNSUa
Ac/tLp30H5JNG4PLIaSpX71UfbOBdkJtINu/2WMUlZqFJ/ZCTszhbz+YpyUYIYzk
NGoACtNCeDDWnv5ZA+4TVx6RyB9NTdyWqsUhl85EL9hbyxE60wXblE3tWrluo2oc
5roeANp1cTYwBgouZpUt8RyIjtWNX6sVXDRCtkCSyxgz4G8Kj6LxWfYdsYsnulQd
WHv3v0+BcyfJPQrk14qmpKlbUN0zRNsGbClF59idzhREmLT4dxrhTcKMtg2Ihrbs
qCcWm316Fu6Byf8il3Y7Wfmp5VJWARRKktkboH808u6z/v0x1Uyk1trV6S1y1x/f
V9yoqPZ6F/NhatAylT2l8FG6p2dNSzBy5iJmWBcfoUE9V15OUenhJi7IRyEIaqJw
zAwoVjZ6qm9TVOKW3SAoOrdUCCSOcRMIfYhslrkZvUTLSmjtdvj/WLwNYauNngaG
E/a78vnzA4ZQknp5xayY9Jr8NJqZxAWsjCN7zp0j1+gE8k2MOfHzzMBG3uaMFDku
YXkew0MxKbPfB39VjyHDy0/Eo7f2LQeRgpkmuSiXdHZW/oRSodMEIwK81403PAdB
nJFUhkrhZgz2z3BvAZ5Nfozp03YdUzyPzh7dqsxEU5rxgJD03DWk76qzySGJRaKi
xxlzKuTbXxIKk3P7cGiPH3qSEEijdKJ2T5PFMcLazlTep6IzpIl9lYM8qU6TPUAy
0zGugd+l+g8O+uqs3naT3K8XLqic90G/VqR5R0dMilZ3WcwH7r7LCX8f3yR0ogDe
EO/CEX03W6kdIMM5KVEiLCfuClyqcqMhfy6YoAstTw1Z7ZxZsRVm2tmr87PGLTd8
fYByrN3LIkee9a44CWNuHgxwW/VJ20B0Y4vHrq4JCKPfYW2jaboF/M4IxIgavinG
sBOWysE1B7bnAX+hwvrQPzx6d9UreZgpsYlM/B9GlhifTDGBHyQOlD95Uhm5hhRG
RvRcO5Z8FIYUnWbjz+vmOu5qKyTXBBknJD3KM+GqIIJHirW2Pz1reVpmC6aclSJw
aokSAc84Rm7OGGQOATaEzymikHgD8SNKda6nJ2mYZ3x2DB+RuqPoq3lMAmj3aWxr
BjFjPqafxz4Mf49ZZmx/3XDQVgBPO/HU3y1i0fXELtXBI+CKyGERhlyKfN1q5ScN
+b38NCM7m3J82+tIUofQutgrpv3WGHA1k9cFgnvS0LuYsE3uxwqKv+8/HiKFi9kw
1x53AJWCpv5fytqCwg7dVcIG4PkWlunSpjL4Uli6eqfuGbdyEPdumaE8kX9fJKE1
Z0Y5DY8nsxGXknMxfA2U+Q/vHhS6flui0NMNFa9UhLQF59XbEa4azQxmIj95iau/
EOUDRCNWwp+h+lbuIETdFnS2qQoWjExFBq6XKXtjVq/hXDHfz9tkcKSvgEpQo25S
9WJ6wrO2Abz6ckRc04HrYH1sUiqPlLxAebqkpY2f0LQNTfY5JxushcDGMB6kck+L
p/xt9mZlzWJFKGFjrhlb39U/B0N1RuMquxkGXK0s7PzV6Z2kT1550C5gbP00W0d1
oCoabrxiaIlwywiL2RbkJEc3jJtct7dnltYstw7RjYHTsVmRFXzkA5E8/5diFcWq
fNijxePGzf2PaKiqiI7ecKtBRi1NUqw+BIjA3paWCeZ+wj6jJCoWICbVol8jrDY5
2Q12DyCiz3SOkSVRK5nmpxROZ1ia2zmWSq84h0/iYaq8/DPmPz/G9kJVnOIbVyWw
EH0N53QUE9ByAPSK1PC+/Q3JEU+5gBe3sk4IqrjYToP0oBBpHzLW7mRfLhMiVkxB
QDhq7ZQ0QciNFdEGqFFtGm8XI40SvYyM9juswU7aWUzaq0WSMmetxnnUUu7npIO+
0phSDUN6hQCe0V9vYNIH8tiJ74Zj66oH+Z1TjLicqcIUmMuoX7H535frlKMzZT45
heDrNuYvwjh/4D9iEzYLbBKdLh/IkFKiwFH2NL8/8TxomF3OdTQ9IboBQDshrYFs
6j39s6vJn+zkv4vFccliSQETal76+sMWKQuutVF63GkcadLtCspvIxgRXhyZJ8UR
XcfXffALKlrGJLlLVf8OOqL0qa79wXywK4F5cFfbCRvFOGsBQFwNo21D9oYuRXor
vyKbRr8t+LAJjqs7N62sDBZ4A76vZmdqrzCCTIFAHJW1k+D76Ww5dNkK1osFpKHn
KAwob6e20i1yZnhof9Vp5L3cYax2FkS1uNXq04VaZyOeVesBHe1J4zw9hKREI/Si
VWt0jA6xhnF+AW/txJOWv8aDtfu7pKpO5AxoALu5fr4G5Skgazi0fZ8KVjp3cles
pax9wTv9RlXpzOe+Q+RHcpFvdl5jNzS3YrdMx500BFlwZd5/17bVtjUCjSuk0V+W
0h8seOPfuUjq+N4kYD61YFezISI66/UeQy2n3BEkLxZkVg79tKcXiKtd/bPUf/LV
B35BBmjdZf7QZhuQ+PsCEGtpOS2xd01sNjlbIlq4+ziChdZTMv1ueJcVPS35HzM+
wshaoNXrSNkSqWi6meUtBFR/w/0AKcn7emgBG3rHb0r42NCUCDBLuVEDU9GVL+Wn
HwJlxr9IRA8HBMHh8YHVGStMaOnhbaOhuWcRjeoP4QdoJm+EJV89WrqxckEdQ1b4
vWUXhk9Ko1yJeDPnoLDq2Js9DMylq3/5l88c1C4Erh1VukHi2BWc7z62FdYHJI+P
o2o8F96sQ0jzF2bEhNP28OwYRt3lrJDl8DUyYhKxRA1escjk+ifYSkJcy4jWo7mC
YWQX84a4fJa/TjHQEnhX6dOopuKOvbCpCVCnpuDf4D1sGs4bYVZxSnIO96rJeyYQ
faG7Voptjr7aZlImGcMNZq3PGb+oG64u7pEwzG/Qe0t8nLXWcr4i6KdhU5eTeQDS
otivADwY7obh4Prs9JEFMWoDuyi5hEkolnTzXMXzKFwkYnzcPRetoyJqloMZeEAj
EgRao6yaGDXBNj+jhHjneCPSD9f94X9FckmQY6BM5kE2IbzK0NSgVAVq3C/FAv1p
Thu5QKcxzFGZP0tq04VqXKN3p5x8EykEynxf7V3Ox25/QSLmUZ9B4upt2I7adS/Y
QveswfpROaqdvyPSSiGwt3FmMe0IFrx48/e3y81QaX5LtWXJiQArqMu/SqyRshZe
t9vm1Hh+xeOW2YiEfCtjcnUnGqF4del8lmNTL7d1RVoSYjmd9/++dJwjeMSjiZSB
tpKkPihw6tMfR0S+kgDROF5sJmrm48yqbrbNjTlbCCYcxpeEBNbsVHDBEqPbcHle
qtLHVzg0m0ypJtf4qNvbSUUM4e/q32qRHEgppgYGEfUSC1g8TMmkmnQNIZVakMrN
PmjW5SaMLyrk72ttGJDp6LipzXi5xK8EgaKxtMV9q+VmfZhViOnskee8eiQLo8br
qydOmvB0tFa6yjhT/JPVuvxJqES9bL3oYcWak71UuHts9SfQIogfIBhGV1KBu9HX
hPqXp2nXrxR7CRwQocZg4KRJJXIPbc7BXrm8MrL9cf/qhCufyNNVsP2EekQkTr93
Yj/ghVyxRjZrKLtRxcvZ3XofK/W+V7+p+MoBDyTklWTpRtG5Xmc8f3ztrninq0+z
WCanZN54U4qfzPTx3nX52JR1Y/vkHJCeB5auxKenXhRH1wT55hC9aOW1GuH0KyJA
BsnMJGbGbHiRF/rletYKsmbNYHlC0wbtZBReV4tBXzay5ZA3U4e8hnPEAOz7kLZ8
j7dRZi+4+J0e7sL/8b+2076jk9d+uV9J7gjAtEVyExmqAi4ICKXN7TtrHKXM8ljm
1JihB9aVk0yf6N9t+2WNm6MByeG9zTkl1vv+for1H2bcs7elB9msCFKXR8U4EFRQ
3OiHOPJDhPJM9jFrUTWEV7PEA6MCnolIJ7sr1pmlgbQAuG/FF+6/FepcKXuQ4pIF
LQHjyp5I4yfmUS5LJALKp/fJq5RSz/V967cX/U9cROa3rYcMJojOEnjhCsBp4TNN
FDdiPH4NKEXKxao1imK7Alkw3HwpZSxfO6vbmwziU6d8i8Dh+T81d2lz+fUE+HN6
9jW51MgeNbeao/E1NuQAvanHUN3lUojTYLRw6poyCufoHf2Wb6WNiapQ3SR5+b8U
SKnTvhUb3/CYK9KgLVH/SIPodhsvijsRbVKr7+K9cHuxfzTLbSzQ1ZCToeTYM8rI
fMP1VFbQxwRPyRDfCJ5IM3cEfRo398wN7bvL7cZ7aZtbc8JXEGM2iRo1NDd/Yv9F
C8iQZQkXQ3eqaiNGHQqYD+vSzxdnUT5t96ll8NongnHifzWWIVGXMssouJw2vcs1
yuTWbLBnMSuYfD8I93sjwNIrEzULIYeD2tpjOKFOgzGQLSnuiCwQTr8jMfsNfKat
4UYQ0soZ9BX/0BcT3YQhBC34cY0IZyzl/0l/d0MkRXpfAAsnUD6QIB/e7BP41V23
6EXswJyQV/Q/RmgTHLlt+952Y74QnDCEy0BkdRCsiwJJwFbMSNU00cjFreSaUDpV
qlF+blOhKCzLaxjXRUkZaZ4nMrOQQN8OuBKHTTEpLmzteKcJA63Jx/I9guYibDn4
+HoH1XqDP03DAHQql0ip0x6FiRiO15WTJ9jXbTf2ok+HDFHvAoixrD6P5e6kFUAX
jEzL6VOLItd93jprqkrjAcy/PhvtZIe7SA7rZFfWVdJFV/8PbfqyhQyvlTLG3M0F
iAkDdNfUOnQT3+y8GYf3Yl+e3Er9v8XKYwXwyxyZ4PQNrNlplqDZePkeIphGqBjt
RVJ3xuRfdKGxjkm+Fs35AXJKFaRIuEKo3KOmfzoSyFnTv2wNqtJu+JNfwFZPZLIu
pqAW6N5zjcXmOJ0jeYgFINOpDI3ixajtUxpVUIR2yM7bRpGg5qLBE6VPfXIJk2jU
bcdXvMK0hdErpkZkGcVW9Q7nTZt5/teRVOdr87C6luZppm/A/ssbVwLPy3NS3DOU
gtP4TFj7Dh+xd9f7O88BOAZyvnWW3pSy8yBp1qtvCWm/TFCjaDN1atz8kNy64u9x
BAN+frOFTHIfocl5YfwEcVeF2tb64P8N0W4besoDSXGAMC7GPCpNXWNlzy11U6lZ
Cg7Z6vZ9Ks5HuMR54bzJqUWaHm9LqWGjYh2L5boNFM7pCkyIZyhdyoG9zpFqM/vG
OhLA2KY6o1M4s4iaNBfxO+gNjuiJouaitutPRS6lps5QSf6ei7KV6JZ2sTUBrbej
Y6aPRW/l/eL+U/1yg4fuvF5eB//IZ+/YK+HmENdvDTdjDJDG2DwI+2E1/evg1rAm
o7sI6cjRytm/l4BwiWcDh9TAhzgvrZQxyjqg/iQUpNnjPTRaOojCW3aNqjqehqlR
9k29MR5rmUoJult3qSj9uwkEEkj5ynafdrEt/kopZkFRgikn1XTPyCj4qe6UVQwf
UdiY3Dvlo0jj42yKOMIGkQek482WLthHGWfiHnxYLrEROy65nk7ipCx/9nNkrH6v
qt/uiQ3qK+8k0p9hf8xtkL8JXlunHA3TWbQ/tD8P0EZqQPhEQhOnRsDVEzw56VTd
P9EqXVQ/Z/99ZvbyJ5vr+A6UeRw0OSCNYQU05f0PDv0lbV+NxoRg0OKMeKRrf7Xz
tyUEtYEkuxuAzylHOBvOmkpHCwK0jIWB77qG+YkHnkfvpadiZIl3gGOf1/Nc+5sc
OUPx0gxYc3jRh/bABj5jah24ggL37Cbad8IrkFH2T++oIk090UcFsI1mgotA5paD
2IMBFJPPpoj4lnNZtMQa8umPEEPnzkTp/O+KTy0DcDy++APFGs9UjG4GVGbRO2Ht
q+TaiOGUlkoLkW5gSuvLgtcEbNtAezxOJ0+eYSpDBShpi3QDvdq1eRQOtGm7bANs
D6FbxrkGBQDXIPlTn0Y8tqBCRF7jfJ/UUu00gnPYVvB9vyc1NUXp1kA5tnon9iM0
W1gekdB/NwHtD49IC6DoLI+qjIRC8CkCRKzhWBnR6NE5o6cWQwt2FD89QIV9OjuO
C1LbV1dl05mbgecitioxq2o6rSa6sI/JaXln9ByZf+h1rEafan7uLgsBXeKPi1z0
woZG/R0aMwslXmlPldDOqapwKHKDXCCxd7VCCLCirTDYDcbad6X7lJqnUQPU7Ui+
HOMp/0Uv2cq56QdhQQ11HZ/8gksWm0LQtJT4SrN5+K7Hsfx43A5xxn86iQrWut3Y
EUM4eRyJjd8m34IuipdWmnCBWbGln2HuTVtYsL5+98jovV3KYlpwCHzCxXZpwhjf
hdDJj4UG+vQKtnfNjWL+D1NpXKmk0PvhXlpzYkxx4pKAbcrHZhc1cQ2h6g7bdVyA
wdjkqHl4hxQNC+K5lFzrHBhDQW9HqNIQTuM5LRZ0JlcAduiZl0oYpI2YGE/K7Xba
2q2LVvOijyA8uQLaR6VVdz3/YM0LWM1p3O2ESL8Wba1QIV7gTX69vtQYkJvQFmBL
9nuUt1iNCXxrhuGk2O77PSd6qMQfbq4RGjoj97vkQtooh/zL77Y1HmZ3FYwWDpvJ
6T7M6R9oNMWuAjeigBopJWiKfiRCcbuwPVnLZ22kVsUa1uNS69aqSwXfwrz7uvWT
+855OqHEF4oeSYVPDWnrXkq6aXTaBNv0PsVj3HPurax8TsV7wyLstn4QtvLyezj0
ac3/Q4kAfUIVFY9dGLZMBOsbAoMKohfDA6NpENabKzZWVvtabXcSSUpmYucWw/4O
B0GA5K12+kQYuhd0aC1YRd8hoSGP19GVa82frq/1QmHqG8UeeYZHbJyvRU9fqkKD
Jw0nDNPIojWac5c4gJ8D0Y1cSNklAXkIPBUPACOu5iMk43wFaXGXD+MTQarlC1Cj
C2LBW8hkpGiaxyhh13wMsfqhN9vYJ269jhUFbrfNTpxVsXlX2NIdIOpcCoB24+T7
wov8+Yrs0r3qBeZtxwDI6sveHZ0j+nGKjP7IzXSQdie0tEKIfqT67lLwyNx9Q+Fm
eX9RtCrlnJMvPmPTAyF9uQmxgXF0bbFrkoiuVGFwxCiY6JcQXy5XdZ5rZ3hafkoe
3kuZT3Dv7pb2w5yy367Fj965sK4nvH42NXZBZl/1uaE1Vg2Wso08saXd5WnHWZRD
E4SDUnwI0uCv5mYoE8XrHAAs1iByTSSWQg67VfWEhYRzMBgtAhU4lSjhDFRgwbjV
7SscGJbIhA8tV2DIx95tJAVoFjlOwq1MEeRYUkqSYTm3OJ+5UlHSKiJAHGF5YUPw
HbDPGFXxbH04yxOq79UA2hxPgvL5FoPSKs2/MKD3T/BDAbo5ksRwTKhUE9aTVEFp
LoRyUFHkkQE7ueCb7UQZpmRi7vKQyGyJPOkrp60xaQQD0w+c3O3ShJmfxTjBW5IO
So5u3jRNRh8AjgTCejqfXqehYYwp07zs6nwckEbN7btWrnozNZzLaChhznK6KqGK
MYrgA22vR7yrrj5t9ioT9Yt2QvgvGJylV+BenHdXhGCAvMqx1wPx18diE7tRP5P/
ZDy35ufslaVq7e2XHrpAqvBkXc8mTsV7Ptxg2JqtHrX+pEbMJ1scCyCP4GsXxKbl
Gm8+H4DoCGCDdRfnVsvi2F2osOrWq6o8+OIQDM71pJhcJ0fhyKNT6xk1Vgxxt7ck
Zesg6N/+Lw4znSdyjRmfRgd25ecvrppVeyTFrEeGmz6xnThUf/sBuhVll4pm9LtV
Gkf0QtT18idqKV+bvmQdcVT3+jpGYTi70R1UjCOhNTaKJqvy7vGW+x2fXBSsso++
SS5Bp/H1r46mnO4pchg7A99YEI9TNkhVFiX2tcW/2PCG9Pz4wpqtmyZ+/Bm3HaY/
ZJw5pJxDD329JEXDfkh+mNjr/UA+WPxTfjHxiS2QSRe9cdz8EMnJa/GT48ZO+tpm
WzWOxwXsUJIvttrakUM8H/LtPCGUW0cFdNGUh/BUBDlL20/KjSBw+rNSbm35OnIl
8zV00xlxTeiZi+idpYJCfHAqJ6RxG3xbhvEJKUrr2cx+q9bmWk8lWV22HEmIzlr3
5Zx/vJ+J1Zw+vzOqpDMc780J/dJf9wAyJL0PbwyvPAdQgCiIuo37ZbLBWtrxAdYF
DRxRUliZwlSYrG5OwpMUU1+y6wV5VfQmwxRxp9mMGHdmM79P7SgvpNd74ElWKDF0
wF9fsQKU3K4CanieIpSWnjsupCFmWl3DzzMrCTKIH/GvtrGJGSk40SjHfjskDrnl
s4t1apv02r9zYM3gOFSbeUECpgfMG6dpXrjuGCyHVpxqCx6+rBQtf9UOKdsunN66
IRJKTUHC3q1SkL5Kw1DQ227Yop8utBTKeeDfVLdXbRw7vW7S643MtN3dNKGuX4Xq
TAtVZL11nQI1LreCfxQA9lYDyzguGPPc5sG52MNiYFewE1i95pP+6wvRt7md5Uqm
K9KmDDdGA/l583kilr1gBPKZQxRON9vuMz8YWT+30x8nJEuhLdpxsFDoqKy7mkE4
Gr4sIgf3oVludM2N9OKgrZJJ3+uSCFIXJMCOzSjT1WF5HoTiJkdcmd5oDpFAHftQ
CFbX0VZQW0iJfbZFEs4UzESIgELrQ/7YEGB0+0vALGPBam/HEsOM4K3iQkSnGC9A
GsX8T/5FCkdRTPvk4fdNQRvQIwMmbUUdUDzEZ5DEA44it/pe2iQGs4YMrQKrp0XD
3C08WX2Mvu021hOjmQcfNrpVWYXa19UHAzB6tiPGYsO9zvtHPx/Qecstl47dWJL7
RHk5IPcx3y0dS1KacpbNgdJGWl3K3qqPg6IA5ZszlIpHAu3XnExLPly2ojNl3Cqh
AFQKeWIGvnX6S1AFRQ6yORA/rnYRb0fUc5JuAaCJDBJRO0kyLYoM937yCM1jSOl1
sJ29SjI1UpZhPkJ10UGqxZrn1XvcfHIMYG84U7wSX+CRuy35TeCCbTl0LsHLVItX
yvWqOnAdLVgWvMhGyo8En9IMWCxdjRwWvzmS2EQE6ZOb6Zf7qJwkoYRUoH8WRBwF
18SwSJAsCZmd8jGg3O+dczc7ppEQQoRQfjS69jGyggqoQIDw73hahYjLvTKwxXfe
rY4yEgf7htQqBL8AvWtLDocBGfo0M9DZTBWD670tC4rGHx6l9lYpXokB5oefmQoa
Nbrc1x206b9sJml7V/nYqciw0djhZTYWlK7Pb7HAk7p7W5yGgF6iws4nPaQnN8WA
s8mw3/yapew2UjC1+1Zfx+R5jFoPi3CnFZbFr04aDCqy/IM9R3CFeHZkKJwh9SLa
BLRQdHP8KEoEG/fDqYoUKyIL1pb9iLljeVHyP2JsOLjof2Sc+kzbCetvLhsGd/FA
2GDDC71/CnVYruoxQjN7WbUkhpzo/yhCWPO0UKL7/PH1uHJCZ8DeDouzJeMpHUaj
3CNku9l3zdqDHUl/xZJ04JwNOA1LMxvee4LI1qtFFrHZoC5OtfswCviWGCIpxF9k
vbvW9jQnxRawn2oz8ZeAsRI2tCou+IazvJ57GmfiNmqxi1dRlFwQGklSjhRRh6xr
aiJ6JX1H2w1ZURW3INGIdJPKAZwXtO/8NGPUca1FXhcUMjW1W9WwBMqwSij4EUa7
gtWvYs7u47Z1+no6oGZB1VYuQ12smBqZGttvG1X+xWJdu8EPku6wc5xPehSgaSVe
g/GdCA+QPOYVCLs1ChA+pC2xmjGzAJgUyuis59/JGSsdaVYkUFwkRrEV6hRyxK4w
6Yr6J17gGEmA7IHOernxAc7U/zrqRXvnFAp2dJIbBVld3+LVOB8lKkr6iGEYQPjh
DJbHLVi9O5r7X8JvANb1Htx+Fm+tavhgxASXZzDTbj+yaDtaiYmxzlawymiuCLWf
3DGnEYtX/pJvN3tUV9m+sMorAhYsX42QBI2hg41BbZRvRxiNzQziCIpiKYM7RZEA
Om/wJaLbNCLISnprZEUiBrmdcDZip+snvuR/Z+vzwWlY27T3jS4VB0aQTZN64Det
eKUUVK+To2/Rm5f5do6LraVOsNhInD54qZU2PkZ3nAQ7/yp4pUFmo0iu9lkAgflR
aZu5SoKX5070DJxEbCbJL10TBDdBbmoHlPH7ZxbZE5CYilIK7Lx8Nhiu1vlPEfVp
kKqAcSki78yU03VBt7TtmpJLw44cqbvOGehYpasW9R1XFByJKo1zN363XcJpoXFO
3phVAChNF8KRxsl/dpRQZ0zeUp7WOvrXoQPt/TemFMzrKnMW4jr5sdlsxqw7JLma
wLbSevZczVkS60T8YvqwcIQOQhjp9jh6dxDoUGgSANX5kUGZrskV+xhS9r/LXAxr
z7xdRceZVJn61eZewnBf2EFLNtgD9FSfsomp6jwDJu010G1FPDePQMsG8Zhqac56
XZShBhG3q58iVIVs8wjCqrbZfs9xzqSvjXIzHnsAi6i1NJuJY+mb2NUCtS0yElIp
bRQKm0t3giFhausoLehKN7cN34tOGH95FIPK1Zp7gU6AEitPnczdpcaGssQ8Q05s
eJNQRg39iRFnjOAjxklQCv3sRGANAkS38H6dm7dJnFqKQnE+JjANw5NBJUhdX6Ku
gsZ4bgM55kDm4cckN0myYOBha/giPCez9URtv3t0jKExoCgv16NH9wDWWtoIoQO4
vGcA7ugDB8kI3PoStA/fdMmLPyWkzFhQJnQzLjk46xBEZ6r2qrKf5wjAXbXPBF/e
3ESRZF1OeKqfB+IpjV1Euvvr9tc/zsFSe1dEWQxjMIJbyD2viO4E86nUPdCpQMsM
8POiXKQxkes8e4o682qLLl8/lIFaQOSum/7LWhvMIuqiUKWv+nkc+9Z2OWCkkNtp
8ZVHNUUUsoT0UPColKf9R53fASg4RqndbxtiDf+FOW6xVtUoU0iPDZ2nEvRuFLsH
dc10kI+g/SvXvsIOH7zp3HVXrB0GEV8pz+mJiztLjvr8+lYsBkH40JYQ2YriaUrv
Ulwx8IOZtf8ti7PsmhXaoJGPorq1Wpf/Kjc09LeHwVF9fl96rH1RcDTkzOxGBzFQ
vFDrZOfhdVJHgQ+VYtkyKrtRwEoXrYpljGHiT0YSCtI+7JV9nlbOz2gcmGlZjs96
LqXnJIJpBlmXE3wqMvGoi15uOUem/roE30WSFXVwc8ygn9G+CxwwGg54ux61krGr
T1emErzWOKYY3w4ign8dO48+J6k4vr3kT/OPIvEw+PxQYvzlGCpUOFvygsln8xQO
Tht3oL5V19G43Z7osGLqaH/CLU/8ApolAllehEXdURUDq4H1zDqZwIT3VcGNXtaV
XvdAQmpjlk2rpaND1PGGJqk4fcOze0lgZHAkN0w4fqSE6db0mFnvizLyeKzP7m8T
3F7shMmmvFAKJ6BkMqtDR7Fmw06InF1Gg4qU3kAjUYg2KXrbf/Z/8Ao6uUxuSAD6
3XT4PlB1w0W2NmkCWRFbVWL0mxx5wZN4EMDLIIdk1z5Kregw1JgndbFSE/6lYkZQ
W8lSmJ3OaVfQoKnFGe43966ecHx+SPa+v81juGGtBlgsX0ELP6vaXtcv8qvDCEoo
cG8e58+tJCRcIZm8N78xkBfCv9G9CW/5YImbnJn80duMgogG6lG6Yd3oH3kcX02T
eAdToiDPe0X5rsf+1pEK2h+xkWO7kI9clHdl/7zFmuApW2TWeVS6s9700Lpz8hIG
8m3pw0oyICGdcBIKEe6rI/lJxLGJ0EwAYSBaAhIyhi3dzvTXhF54phN4oyWuEhRF
9lcofcqPx/mU/6Ou/Jni92q0Zs6mqGpThSeeQHs6uFyEtIUDPyQpfl9fb/msqBr0
AMGSeniKpBWIdzzMq3BU7sbOkYya2ix58KClLcNLl0dx+3wz+4mDrhjPQ15ye+Bg
2RdUPsT6nl3EGfl9j/eInTGqqED7yhFhekLCpA7YKAxaHkz3IsZn8aQjqVECAKUS
qWfyVw+UnqrB4MukI0+H4G250NJJlVg407Es2NpMeQ2os6epRYW608E0nyYEpD/o
bGHUHDMwlSzaokqOqwBrBlJksp0UVI/IyTIc7tJTN2ufsjoNLtFDLBkV6aNUuzhs
XO08MucyueLZQ3tmL8rPTzNKqHT7wLtXeKNRysyQkPOOEx95ct6hCgOb4yC8eLs1
vcpgp4GCQNnIL3AFe55+0kxhwqttafWEB2bKFYi1S7od0PEWI1avHnmhyA4qEE75
SFsoO1XRGEmx149AfPl9p/pbgSuw0uYn2iBBKCod6MwsJ22rUQKzPSxlcAwHgCkG
5KiXO6+M78OCVovm/50/kkVAAnVh6Uogp8b8MBJR514cB9f9qUIGFurKEbblwVF5
5ptbNyM8RINANeFtzOZEBuQYFPENKTc1vuyeXwczl5fw9LmEjkcnUtWbJdBjt8Fh
tLa5iwN/eJJ5nMFiNwQ+AjPvTKbhDUaw4auq3Di5W/g38iKp3Hz05iqk8JmE/B8v
97OiNHiXi0e1oiVfbFlDnmr9GEs1klOi/1ze+Tg2w0x07r+q9/a4amvjqlAXof8q
CJjDTvTO6JnB/U8mS9+G3bA2nMkOErn1UbZkzns/VkLw9jcIVT/zDnZCzsLSdALa
Jc/qsv6D8UdCC46AvfyOtktVrfu+RKCqEgeFtuctqjjILi46pjSO6FElLnpq0LEk
wPPStkBVtoEUM/dkeFwaqpH76Mbaq3UAlr75ARWRbZAobuwdxy9K6grFIjkKFuHy
naTLb0jQPic9hMvdqbBaDogQ9C6AII6odm9dGp7/xwO/pHztBwo7AqLBTg/hV1jd
1fIOhH4lq3Y/KCWT5vgSCKYM4okiZFKlPY3UHK9Nz0+CXgTKJwyFlM9rkzCYdIaI
FycoHDpMOdnZFlarXGuKDFg2NOTXikgQIKqkU8vUUoYZ7xiJJbRLBulK9+cIe472
A6DoHs6qLlbkbS7mttEzui/p/Z3ZJW1QKFgSt7iXeNEQfw0iXuc2BrbcNwxAdgHn
txL2aeaSsDoyQpxbwoNS5wNMEJR46/oMnNbSBAWYPG03ESmU4/H1p8vbscFE4RhE
wlEUlrj/GQfKj8G2xAQss+vufqpp3X1m0Pyhri7X1nxE0BupM527X44YYsIUJc/+
jEn7G8bl9B7Nvzpc/mSKOLgFOnfZYPmKk1qRcmYtb1TGYRgEvmxpMxvt8RLOy720
gkpl6rXBiOWL/iB/nnNM99Hx5ZsPIu8S//EtyUIU+0/iJ5KZPftD48W2EAZxMCJy
zUtxUXZMTqP/vHzTinI2CKtqup0UMFOInsyQ+ipfnT4v60S6qkGAH1TXddoHy4oe
Yz49nA4CqsfABbGb2N/5x3VlSiCArMVxrzMtOgg4Y04Xc+aREIkh0JlRKBK7WpnW
rN1v//TB/6JJMFukqNhhrTIiWPuHUccvyKTnyly30s1GTH70WtukDXhEnueWXJWo
HwZFM9kX3v/pJcBDZH+YhazP9zQ85eJNg8M8L5R6+ezQ8jpfTwRAQ6dt4Otai1Ut
OaccXniet5tnhn/bKM9zeuszj2bcwgSCQqTSB5vgqp0nQlrqS+P8M/mZYdK4ZO74
L7vcrMdy/feBm/d0M/49GxsGKidj38BaIrDyJD4A8IDFOh6RXhJsM8Zgc6MRO5Y3
5BVYeJevmt44oJ+pHjSROxXmgHIzp0iwvAQtHopGGg4cdDZw8oSCfTgRywCEMQtt
wnT6NLOod9jWfq/k4wB4pFKh2DOCJjQcw7VbzpVXTYufP/cpkTzb6Ub6iohU8APy
TQdhmz/tbNJI7hHGiC1eCTxayt4Pio/WzIXYdq++52k1XxG7/PKLYtLssGWdHtsn
fSd9gNXTDDNqGO1Jk5MB6xrlUBt7tfQWePEP3JHP5bEs8Zhwi+rtJ7o9k/onPg4x
3eGudAsTuiuPQQV7o+XsaPk8nwSUPc8mZIgRuasKaIpyHQ6pHtccgpO8R0JXiL39
imCy6BsbM/yE3dM9emXsxhV+S/b4eF0EtAj2GtP4yBxRBPckP2umg/Qc6zFjCSSh
3QSx7Z8BjXoTnaw33aqpJJzawLjwYg1rQaRZJ4o8tml1+x+5xHPlb+sR3YyHd8z4
7Z8ZMEwU5aQmyM1rLO+8+FdORaiwXhE/KcNfAahewAd7SM7vaKtna2BZfgB1ZUJc
B43bq9htA+qQLc0fA50D2QtSyBBskgDhsrZU3wGmE1IkQSnxoazfZRWveNjgGlgg
tJoekV6/oaakWMmPoNIH1LEHsKInUkZcxvbTfcqo1hNucckGjYCb8jJtgZyMeDAi
FAMO7+4XlY/bGtCUPXWPTZop47/en3bpCB3ApihvPSSOQMCHRC8Tb1EjShM2Mu/F
bIW6ktuftAQAVU32VtaU0N0Hww+OQOrE4TtpTVq3dUi3rJLZ7iZ8+JDwduxJQd11
JCuu3/dOlnDpqRu/Ln3RfBc2ALKYuG0lUoe8G9lztYiNvh4BIqQBAMUbpfUEwc2G
4SJdv5qbMETYqj+/pqmgD2b/uL8V6e8CsIzw1GVAxC+fefCs+IDEpK6utIy3fblk
PO+0uwhIfzLtFFFAJtDZlsg+x+OOkl/RBultbGS7o1Z6yqt5/Yz9Hc4Hsv5487Ne
j4yIkOsk8uLQHNOyXGIc5CS02ev20X2s8NlcC6Lww/Zmkvs8uFMogXZ2gRlC09pO
FB5NJYxSnKCWJ8FCK/JeAaHnmcBRnb0wVaaCtVFPVURYofSKotxuWzAS5UccOVNL
MD039gJj+EOwUQGh9GPWBdpoLDM8nbQdON7k6/SA6AOHxEXTcN95OPBx4BxvR0F/
AD16znxBPCEadm/ncf26Ioj+uzwaQj3Bg2CN8slFTIyJE3KPX7LhsHpHh/NXPU0E
lVCAZ/w45/rq3vw7Q5kHjbZtXsSZRz/ct+8MR2J1NHx/WM6OrT03ZScBc8xy3fDL
daYb3bGKtgHCkQjEziijTf0cMi5KROUhym95ocx0pN1Dj8EQcrcJAiXpyiZnxWgu
lEm6v9kXmfwpaUaXilKC1u3mSxOxCjD5vQFFapoqSNJpoeOD4522t11E/K6Ih3rQ
QFMLCtl8ueF2l85m0erhhXOVhWjmf6/RtExySzNj4T3nNJHfJn1pG8mWuT6rCm1P
ZvBX/LeBKbWzCkBI3vwj1gG9arpCwxpSWt3oEdu7V9Zhxd2RWkbn8FGmDhNuYs2v
FRLmbaOEo/qzmAEsPh7XUaMiSXv7eRT8F2qCiKecBx3FVCIcMzZUA58bYTJ5zCjc
qPIeHu6MX1txscL+69IYZp8zspROidvxoxPuDTqAECA4z5GckQkwyHjkujVuFAoX
kL5nX0CNbrqrHKJPS0kbCTO+W8wNgabUc6YEw4WdVEs36PyL2O/Al2ZD+qfm5gGb
WU754/cn2ZqjaIVjwOLXP8eIzOPXeNUIkMrZtOIDoaENkxFD1Gl8BUXlAlSLRqv+
1T+6vaKqSm8Io4BL9ZFmT9e/LGNkoPQjUWCdIwuJzx8lAS2/lj2wi2Hf8GCTj9Hh
s79WCTsQ3azAX38h44IjxIlKAcXH9Wd9aCcLiB7CkDXMv1O1B822oHcx83sUq6Ks
97hMQEEGvQyP+EccPkVO+UTCOd5DfoDH8Kzud32LdLBa9NVR9GOxBaoj0dzYYu8H
OIRog8q3JpOVRrILdgcwO4MF1milw8byuWJ9nSQKW2qlJHafSce4pUY7Cq04AiYZ
htO3WaZnbL8lPHRkCE3gd5k1XyZQ4HWq0X7A7Fpsqnh8/0sHBfJ8KCXwKMViMnnK
ydkceytO6m4tG9JCFOyGw5ovSNoDWgGVUcf6LiC7w3in9CWl98htMdFuCSN4Y00a
B8tiM76mVwcc+KJi14LcogigmJNUseKbvaYZY/QM+PKUiRmU2NmUYPa9poFJ0kWh
k9HhONrcVY9Dnb8RgnOs2NnwCfMC/jnabQVNLjEhUK42uoP9AQWoCFE29pU/ZQ8U
QSCS0JIQevoeBE4mk3qzCUHHEdLU8xTJzYEWOh/4JWCe90weZiMyI5w5TQqM4LB7
tw2y0sDQu7b8XlBtmpXv3G4HRjesslhYXA3ljJN4//tjoLEoeNuIhXhd9el/fKyl
1ochRhhCLi/y0Ol+mlUUUzoOflzUE11VTnlGRsYxHWzdQSmEXgjkryGq4vMcESH+
SIhjWnWEESKKrJH5JnfC95HhD/wgqmEgO2CIX7xuhsW1fTwEJUGM/ooeeECqWCJZ
lIy36wFvxtL6wFsHCkFc1ZbUZ+9F/mvFySeZV1YHxzHTdTBGV+PZugm0zq8cIMwY
8VrIpsygd3BQR2DTww7L1TSi6aQhmAkPl8yHXn59347TSRnNgjhcW7AmbCO4yT73
pPzNw5WytkGh2B9QrbkfVkxD1zzOFjnWU9N1pgEfIVv9qUmReJaQYzsrb1fLWg6+
5w7nQSv8wHG0U/ZCCvs1E6ZkSWzEi7C/XrfIbD4vOZHbpVglP+jxOS/nYwqKZ433
Yqw9F2NWPoM6PHhyYmXeGsrlLLq6lh4p9KdZ8k/g3vVMqy1MWVoMkxVB9S0BuL50
eZ+522fSVKm+SnfoF61Qjl2VY40i2Lhz+JPPvM5Sy4/IxkF4xEtf7sH+XHdDSIlp
YoIcG8oEP3N68BsCi5CWRrLB0llrP9lx8pt3KSpw2aFAw6olABpu+ghhB8BCRSiT
H+WWCQiYMRFO64EUuO4jG1xAUO4MCFtnTl2fmNb5IdM0kQuLVCJwSg3/xDvGUuzv
m+9G27DEs/Xpx0vwLpuhLGxN2XUntL4qbVC61hmGvzuqlm5XxaHD9Pu++wexLWt+
o1VvMOdTFQlUhgsaVkg5bo16fRpZmSoabSpUghjcr447zcMWlRiJKlq+Dhqk6Dx0
58L7SCPgfgPSpnhdTzbGIIuJDtQn9LYVucrILcWZ9zbJjI3zZUleKL9jB7frhpqi
CnCk8hAwabSa1zodcXsN2shYrBVEgIwaGuny/GYLEEsefzDEWz/bcdC8wIgzgIk3
kty4ws/Fv6rDuFauLc7hWxdz3Ca57CLUvS9GNdQmqXMIw4NDNswIJED3ywXOTbPP
0juidngyzTAbOSclBs2D+y8MYxTMDO+/ep9dCol/t6atekap20018ataPcuTGTKE
ntvY2a97MHW48zthOBd7oGHBhsZins3d1Tl1dvgZMYU0gSrWQWbj6DFNskfi3psg
aq09yeNwLJzRlVV4DJy110SrAFaf3eVJlvnc65BT7z23H65Uat0/BuFbIEi+rcp/
OARpRQZiWT6kq+4ghm9FhMF6Oe2G2xhT/ZWjxtjU5YBXMZjGVI9D/TrN4Ir0dhD6
FtTxUGv5B41EsBHEH8GoMhndbUR58hNxXxTb9Fq6IncX6anGBAJS46xa+pOh/QNE
fI9nVYg99FtPi5u6eV/tnVfQ5FdrLYlVLCuMRhVQzP1H7qfQldIGfE9rKZ0usoWc
xm33gTRQyFvYrKfkzzhaf2GW/Umb990aSxSirt0cXy8fBmi006+t07JSYJBFCB9Q
8waSJauJ5P0Rh7e+KmMNrnO6hQnPqxwV3Qv5FSw/RXtdxYAO0CRvhS4ot3Wtr//I
9Tj8h5p/P6BdEpeuHWYnZJ64PyTA3RmyFgWAdgG1fFBGAvsbPIs5k9mfqeNL6dvj
P6RLK6gQazDrn2xqbJrEttwUhrd/Jpy9XsjzegH7QjRDuNfyb1M/5uUMja4H7lNr
TxxQEczrvx6LeHgM/pks84l7Sm0MyxcvkIt6QGyVTU7gEMyVWttcuGnKjM7FIxUJ
IML5JswEpKupXt4k1NH0GLZkLl9GmU49Rn4T1/Z8rjbcjukpmpabncznVjfYqU1L
P7udoYZhfyK3NatHXwA0gwPtuQjmfido/P1pUdFtjWkFBZbRPVnf01ybMFEn0RO4
V25UmMITn4VFcbEgwhfp8uS2KLElkSsC2ktd0kA9nTYGbBpBrMArxIE1R8hJlvay
jr281kYPTm85vR/g+X6yXz7h4Hjw3QUI2OjaVvj/zTQcY97sfDJ4de2ZVp5qjXms
2giMtxnWUM9xp/7MIUGJBZT/LgpY0kYtohm9z6LxHYHOB9WXWN40QbHw9WMvQvym
cxfH18KrUjdxlZbW37pooQdfe6fgooekzTvg42bgvAx944ON2vlRFSL8/N04eeyj
aZrPoKlXyuq7qCibTNSsZnWwJncm9c9HqLFpcNCngArubVyU8xsHvyoAGb6Dt2Dw
VMfaiL+zHjsb7gInZ8Z2TC4MH7yR1il/1jqyeVUZLlXWzmhdW2ypLIPkzj2gUWnZ
xY74/H7XA9m4l4FNF984WP3G0S2H2UOnU4VSKrAyFxMoRc/HcEuVIVutAFjs/SwE
98SvRbKXx+vArE9AIh2wkP7xBK7jRlkGz4cyd0rV36rUGWlbMrrjfFm8yCuo8KGX
E7fSp3M61dQW4UklZvxxAGJKYDr7IGkOk8U3QcRzv6Kz4m5ozDinwUP6VR8dOJF8
0ov9SjwbelhN4pVrtoIkcjS5t0nsa6vY5hrtwFj0hIR1ZarMG/zzlc2CObrPY1eN
mssTybvxWVzLYRmxA5Nmfsd+VR9S1zPbdcVw9FflbxzXVbmkyo2sdRs5gu2p1g9z
GNFqPfvNOyrjC5Fky+BnYT3eF+s99vomF0gj7KsxZHGcCJ5LQB3lSjnc7oRoFgkb
LmyTujnoR4JkFHSJBLMLElgWIpZLhghbvITffQEFb2F+QKcfHPUJN6TbG+1dAkk9
pg0GwAo2mNjtuzYy5c6L+V+dL78CnFqVpCoiyW/E3yFp5VlvNPVYCvSAgg5wyP4b
0EM9I6kwNOOZJSjg+8hpUX2fjsUa/dMqcpgUm5QHj1Acax5GroC+1FKbtEpPLHnY
xxlvk9v0xZr5CocUBRzKgPMiDqV92U8vbD1/wVnTEs+BCSotFsX3mkpP6q3jnZQg
BoQGpavGzJ5//gZbASV4IF/g1rY6Ukg+31SkyZL8WTnopTGJZnxxiqYng6D4Blg5
Bt1DL00EzRrjWKAPEpZtf/2Knq5GU3PhU0sHk1TbcUWYjH5QaHKDafkd+Wad2v1G
7BoqYUuh09wEagLwZr98QIZjJIteHXJBPV4CGE7/ANOemhcJQoUvp3+aPyDweajN
goa5yNsdFut2tXYXZab0SDeo4D6Jb+RbhgUHBVVYYrpMEFA6yQQMrg2jSnQ+uEVi
AOyb4UAWJpqwZtR1T13hApK7PswQWaF//L484PD4pSkraDDvlvQCGiBHKyIpq7oe
p7ai17KVV9SZ7EeMKp5/u2DzOGxuH0Es8qV2T2f4WEb/0wZLnTWB8QYoq1DIyPnd
85W9BS2LHZRbS/UhjGUEo/ohSMQQd+Ca7KjIGh6Mn8ERiwFqo0J+eZ5U8PYcJjK+
wp37bL+FkDEsPvJqmXjhkwKU0WA0dMmPJJt4rKL/PYaMAvmUXI71AeRH/x2VBsQU
JA+o8Fi4uqsH3EdTnhlH2STFkbjXGUZMuEuRCHrksnjqHyfU5fkujBg+DSBVDPPq
TAydlniLvEWpXBoUFgYhPtlrTb9CbZKGwp+Wy+PD9eFLPfxKLbQwC8wqt78fcTl6
+s1cjf1JTYusMJbjI8+facpN+mTJ0adN5qZIc/+Fz5+OigrcdQdpsph6gDGoCT3f
wS+HYuhA+X/HnRiRnIRTY6RMqaSyUiYpyeu0uVzoyK3NveKSaeNg+0PCjr6A38Z+
4oJ4yXYBjJ1uTkdIccfw5a2FsbGIaOVDp4a2ZC2sgvokhnyrypqn0Vq1PrZLO29z
ipbdj7pKJgsVaucDwDGrAyHbktOp2GKd1CiLevHeQHUvCHVEpUML9+SO9M9+X4L4
AQuIKlU8iirsKQ5ADgFzJryO/Vg70rvcoxFpn1JPoFJ6ppseiVVdJeXMi+A6NpJw
jXsz2wyCYMOyd8SCfyF4Xd2gnlpuEHPXtk/Z/OKr9uxt09KQn35yTv1ceFNliAUi
5ODD+djeq2aMRWDkAYTLcLHaofjVhiMebYtYkpbpE6dm8Ijpyq4aXykWElPgaUQF
JRsWQrY8mCPtfVaGJ78Oy2vKy8qg5ySKEDhKG1G0u7FCBCC3NkWBIJhnimOwg+zU
qwna07Jbnip9fJitV7XAlgkWzxzFcKwwTSPaEp3uUdeMVQUVMginC17q5PZH45Ru
d50i2DknBvQGWjFNwGv6Ppl3optrgAaxUmJ57rDLhrzwEBevngwvf8LhgPwVOQoo
Ufh1CNReFP/n3Rb+E8rvAyP9PB3DwkM11o5Y4QMEiPM7HD2GssCJCrfc+zWxniNE
cCYuXSQ2QjNR0nBk9UPZ5QAyMeh8aF/Ygmq1cETUpBv1SySSZjmykQ1OycYRSMc1
2+retvwfJnK/zsXjJQ5irHOMX5TgS8VgOJBcrXdizshYgWxwJnCCvmRDSYtFRJyc
v5pGndF4hM4HvtUUDB1xQCnQsVX2zpCkHF/ZgkcF/XTTHiUYAgh2WyUNtduEFoeY
IjiloqTu9BvDwyOPr5DthKHmE27LJ2vlljgZTlkqcR197fEXHgoc5gPYS/mBjwTh
+cVoacLuy9+iC9cLXHVXulymZE1uUjV4ajAN/oLdOgJQp2p45kbYeBypBuB8iv/l
ju0M1NM7cHYlgtBCd3oYoqcA5g8rQ/hTqYLHlMSvJaBK0FGLc89IZso9byW7s3mJ
sr83CFDu2qPn9uhXcQhrviZxCry9fgTg8Nr5ydm8yCyHfj1dCil/jUfl/uFLq2Ji
pvhG9c+q33uoiyPID28FrKSbZH5aLIGY0uWR3gUEpSFSmEBjBMHU9hwlu3Xf5qjx
vi9rv0mn7ZutlK+iigcHWm9HOnfL1u4YTIUsrOm2dKcGPoCPKkmdGQ9pvRWpKp7w
/kq4+xuf5nAP28UMCpbCNDFNm9U8nHEKW2oomrJxg57IHCMCTxa6ZQiPwWUn8cSw
669ep6Q5pw5pYcFS/HtJqVMNVNrAweFGNK70d4ACEnwcXjPJtDK/MacCzg6cd4IC
nixjX9h0W6H4vesT0Eh739RegDUOLjB42nEt74iY6AgXmwMxOYVk7WB/LmBFAhMF
JzYYa5dvdpnDq8jezbU8CLB4iw4gE/c9gXRfK8/47Fc3kdRAFjwFVOWHmRm4xFUH
lUMDa+2emkIytV14w0NmpK88kLDtEIafCmzUdFNgSo5GYTuAm7nrRX/kQvG5WF1d
94CA/CtedpqtiocUJtB9X6uWCHU/gHQcG+DaudzytWyPKPl6w2iq0xwDSrYFODox
6AKq6BDt+zYuQVeYykolzCtMMAhmeevqeNq/GG3BnKO0sTx1VcN3XJV2TSZHEZFL
Hbav8sVsTDU05dr6wubm55+vI8znaqZuMApflBv0fC8Q5UaRx90yt8ifzWJZOGTi
/Jy2pSGR1Qm8mJe3pHQAqn/5ofrpQ0Cs06gXcyjGwDKhgyX81D0rpK01nSA9QD6g
LdgI5A6DXxuvMzGyWKEm76OcdLqTKA/M35725PPhtrFbSRrNa/bhV5XvuTslMmpv
7qEyEI9XRIY7g5BwLAWWYXPOLIK6FtdAMCo4R2eR9+Ovnf0ydO/w/BkV1zuW6xYL
RH3GJeGIAOMHjrfPyl/VvS++HYC74OYZXnyyA3sOp6P7aywRzGoArkZ8/aYbfIuX
QbyyTP6SftJolwKyhmbyG08WMI3L3F/LidwqOLGKIBaITvo5tDLOkMtttdIx0cK/
hRw8yOjbnraBFh1usLRIjTFa/NnW/j8Xajf0g9RmOzx9wLGMKl4Ncd4awpexjExA
f35sJTfZnzQaWtQlHWPntzCWohCil2bvMBgc5ubEBnWF29jGdlLJ6pa4t+mI5DOo
gbGoVAGhVmxV7ypB8rkhfRu5g+wgjvVfCUnbjPO6/yeMjPa82Ftr+u+9KTQ7WKJv
VSAg8rBFLXBhS0mcVt3Ee9IzlUqnF87RR6DB1TeUZ3P0sBT2+AILBa+/qcphxJro
dkIVLDilnmBuREhIRFjTAyBBE+Xo8DL0m0DFCbMJgyaq5BWpwfohuXgbEV1eChj8
cpRAxlmTIoEp3Zlng+qe/QWBm4PqYcyeDKYW0uMeYXgM3EY/f8RR/P5yQ24/Mu39
6pBCpCXuCbpCHVT5r8dD8tasQ3PgUf/1uJrFCU3NpJRmUtIVFIJBWWxqSqVT8npn
7kWjWuEKpRG8SHW9KejGOVbCZmG40RC+wh6WtBtLBTpwSWo1+lxJ7JyC9SZv0ygB
GUxzNx6XjLKRrSzomPY02Qx1t58vhSprxflBljRlyi+TWA59jiyVSYs8HNlx/Gtz
1CCtTC9pMloB8s80kwWWYIzxAA5SSS4fgV1Of8mu5CBf3O/SBjNhiZjc3kjlQoX7
IpLQ6oCTfeYVvLxR30OcVcrRoxxiqRt09TBU3tCOMI4gUhNCn84xLcG1pEEozNkM
u48ba/Hn1PGpxKrRWPlbQCQ5AdQTqwum9W00YJ38OOTwMepNyNqkWaaLCjh5Trf4
fAroB0hZs31CQnCqclFEJMDrCZIqVZmQtQCYxeXcp3Shkb8f5EyhknvHbLuDmlaZ
Zymwsvkt5w26iwywF7fLjz8H2/HZI4lYer3XGx0AYDCTqSAjeoKq0C5QeJxqYm5m
EY4Pi7WMDn6FUUQbUb0MXHpe/gBKxTFCeDrIZFYkvhRZlQJd/1ni4aVeGjS9YGXz
yU0dRMHdmUQZ0iPHwA4hDZzlJI0g1LPAWgw+BCZP8ql13plJjnJYmOWvwkgAtqMS
AqIwVdJxV0T60nr2E2iGSv+E25KVKfcbiV+8+138Dtjy7wy7m4QsNQobpWBLga9c
fuYr4ujO6E65ineWFgF4xCjOo1QotXDR6BsBRMuq7EP2CgYP6aT9G44Z4Rg4tmsD
IvL9vy2m5BwUjPre+q5SMyc26zyObbdE5a7nhlV2iojbYG9Z9Sqp7Y/ZMqbOkp3/
saQ7PPD62HRvNMEk6GHAPCwk6ux2zx3of21GthaOhlGqpHa83MKF7g5JmSpdJXtf
e+Y8XM0IDx3UlxefbvEH6EWKEwPccfBbqHu5hdBrUbk1UpV5J18pcL0vQgEWjGFT
eD9KnGIPece2an3IBaZm5C24nd8vjbhoeBFNtsr9Ng0r+nfHOVZgv6S61kaypdpO
n0QRVfluntQi76cR4HEgSAtfMklle0ZZM6X1myak/zYfUFi/L6hp09SZHWk2BDm4
OmdyZVkxx7Q5OaVOvCRK6vgvJRizN+L4LXsWMwWn4E/ihR8wPzlTsvG7eUuPjuXR
wrytg3FzNDzwrlMjZF2elIpvB4Qv4SFMoW654yPVRnk3CeO/OmV92lo+9hhsFpRW
ykGUOjEnJp8+5Q+9KCvz5ho6/+08XWQwGYc0bp4KOwoBYaylXGaxDqPGS0//Jlv4
ASwkFwEDYx0nTfkh+q8czZTbaaMZ6uM+CG2ChtIXIRhqh7c0pXGmJpDmRT1btO4N
wWcLFOxh/E3qshae68DS+q8gfcNqWAwYIhHk0grpYiYhI+QmGTIO2ahVCsIBAbBn
09HHUg0uVSNAm6+9/W8WLeF0SOM0yzuxVyHbPQD8R99o2Dw+byrsOeVwihFy8GPs
azawTDUNNqX8Eww1kYHb29VyGK2qhLPqSYYQEubhSDPFwrA7rcoKNdkqxgUizzfv
YycN892Kyd6WhJtq3dB26OSoHxAIx3OGN6M+eD1Pq0CKxAYtI3A7dd2IyqCLlodV
/yvgBDt0SCCwmKyJOXMCiKxYcZXm73oT+F9jK4Oj8XYXeggbMGIGYmzL0qUzFv4A
yP7hPP+MpwJOdBFSyKGu2gDzs3DqD74Y6v1cOuRuRJjsHbfSTwZXHoWzyB881Pwm
uVkpRNSWJklrPHdes1qko9Qc3xHHAoY+QhQ6nP9x+tZAR6qqFMPjtImmHqneysjd
bk/Phs69vpBtyiDiAsQHd6faraDh0zp0CbH5KF38guyx1+v3sfFi5gEl9mKl9PqU
tnTwiXm6FdA3Sy2GKAVClIQESacUvLW0MwasmM8e+DjKMnisvT8EbERkGTztY3/c
s55ZA5j3DLPtX/iTXoyBYQp9zj/h+AhqQnTeT8DUW2IPOqH6Jd7+yFkRPtfcYHT5
C3VaGXT8CUU0ioJ808gxPgPMHVKCxU6fNkGvmX4FZqcbiLudZnGgNhkD0vCJ4/rG
gYdo3mbJKNacRbPzxeLWGrRGAEh1KC7riP7CvB2kQ/T3s47Z0j/ZHcfdxXHOfKCA
/dAE4mBGOwjZeGz2pZnLTJjIy0la1Yigo9sRg41S4rH7yvBk5sPS/3lesHZKWT35
3SUMBc3JKeog/Vw3UgqW1eJpqicd+s41VgE79d4d0rMjJJaNug1lTz0rwCiuWSfq
0Gic4KbHkjVDkJm26dqsSrvImOJX3O/YfASntnsQVAUVaQUg8nqUOZ8XW6IFFqkk
isbY09uGeunf5daBDdMjyqeGa+VKXSc27ILY2bCjIA4G7NuZ1GaWWvQ3Dw6DPgyR
bUocNAt79SxeKa4Ugp30xF+ACxGDJo5syvBHjgYQQigmqmUIAESWtI5cM2B2cZzS
13niOjrvlNf6RRfZLQjv4OQMmcfcD6tMODSwUR/U/QD/uTfLX4Jm/MpygAhho6ej
yDZKN66WWNU5PmJ8NPUd8BDT9yGmoxc3kaGzGGQzuHANE+2njyF1EBd8BEPwq/2k
aZUEnRF2AwTMIpyQLHthxkMc/L9IxzV8VCRbaBjxjI/Hxtofs9aNTO3n6eZzZOtD
o4lo4mz61JbYEQ16RrNFHkeE0ttdP4vjxBjuIgRyB9WGzompYgOqvGYVgxjoUe8V
bH0Ss+TwO/mNQFG6ZWbbY4feN1m/FpQIErNjZTaTneZUQGcKEktq8sF2D3/bxQmR
b5zrDRHNjUJpWJCYSLpLWBi94jk0xbHrX+tNTwo0Zv25rlW1lyRL4r+odkfSdX+p
sgS3+zBD2lWUv+VbO4O30yX+QtWz5C+uwb9qCNnzgW8fQE+0FkK9/kRfp2QQ5G/1
dB1hIkwwgGl3hK6EkuisnJzxNCp+pedhKdMTATOeHrkxuM3y/wWCV7Wp/PS/Oe5q
iwasNLxoazVQAjjwyFZav4twiF6Y2c1Fu7Db08grbAYILALnCLBPOLpr1DpKe9xE
0wxi7PdoMu/+uOXGS7rFEN8FD61ut/Fg2cnpCFllJJr9nc4BCy0mu3sKsPmMYAzX
EINhnqDvkWmjwWUQc0c3yGkdAfZP+QarlitO1IeltNKXRCZrtqlnAuGZ7GJobEbE
AhCCmiuZoexeBpvgaDDwPOqLsZd8/CZG5wikfXYfHJ9doYKWvaTolCRYKZl2trMW
CFqlgpwq3sMKI/UqQp7Y2BxwEfcajin2ryCul8t3Vv3i6RX0dIM0CtZoEAfdBg7f
vaGgFM1UwOtb0KkKcgN/2uS81CzCvgAcJXaaUoOyANVETCH+RY51yN8SPmSKuBtM
IX4rhfXvHsKLviZ+MjtiT9FeoX2zosRrMzlIKDdbAzYvGBOaRv5M/7lNy7rnslPR
NcUb8UwE5bl238ZVEKh8n1tpTGBcN6rL0eTP5OP3IM7BbfGTcsQdJrIYdH8J23ob
+1LgzrqyQm3/uQMKo8Q7x62y6vYZo1/WMxYgZ+LmJ4UftUqFwfwzd24cZSPDj+W/
BANLrA4SqXtAf1HETWyF8WAGOR6M1wJkEvpVD/lv9MFo9f5qS6xI2ZwQEh5CRSR8
SHVTvh+p7hMxO5ZxlJBrudSxcAsnacJVYCko7/AARPy+W0C/R+1jH8fjklHFsOQt
lSVMiazTmW7Wz2PaV2IJFsoTuz1ZjANPF26IkITTJRk9ZpysXOU6L347gAN2aAma
TwJrqZJOxoqsBrbrFnM84X6cX2FNmtI0vehd9nWXxEHPI9DxwHPE6PZ4tHz5/dek
dmzQCRUlszZIjLSKi5913Gxb6BhcRc9wgn1wHtu9TvRStFt+cdA4CKfmynXStnEE
omcebELBwMLkBDOIQQGAFVwAL3GawIS+v7tm7HpbvECXx2DsnBUyiRaiWMkOu3rP
r6C5uFXsv7d90ZyfN+A3ne5uzYaoH33nH8wH/NzpcpqJ9coavTl50foRDHVZ5U2y
hP9xJD4ZmUj7502w/JluwYKU49M3s6vIRRSj7WMm3CvN3UIDZxFTtLSfItpVut3N
ioNkzlWrJqBY2typGphsnI3qSWm2/dBh3msazKV1F1MtMEwDCCtYQ6GD0Gg/M0c1
Ny47I7DGAdz5vT98NnQvIqDshhLJVa1/HISWBUQg7dyCjASNgBcTVkLXn6izTlTv
z8Y0R8NM0boBOHY2HdVgJFDYpKbgQ5irDOIpniYEynC4lLIUJMHR5YXeNZN+4txA
0Cs6b7o/Zt2lpCNF3/o3xXi6cl6SFe8oiYLTozZ0ggc8iWX+Af0cSBBcFbDtWoT4
Medz/hEEEawLCyXjg7mNCwbnJkEON0dcnBFSxQCfuPxy9X9JuJyZJJnqQp7ib1Jt
x4XDjdPs7pqWYEqoAoKI7PkAYHlzd6h/qtV0j6A6OjoO0cKTTLzL+Uf73yYsVEvl
krNnbnos7XB28QhqTjaqMDiXJYe6i87ghpKF6Q6PpfcadKek9cmAZhwsWUD4s0PK
BYlSHUfSvjfvwb491WmLgKl9sKNmixiHcwpyDMgDll+XO1OsJsxDKj425tAM5BKg
m5t1c/0+2eUxZI9xFHaTLtL4Y6F+N+OyJOk6N5YnTc4BxRyc2p53SjXqLxVVO/bx
NKg3H7oM+bx4mx5aZHNeb0ESZXt8HsLYe8fjnhqFYP6ISOH6xaI1wSu+qwRLeS49
/m8IgOV4JQhsGpUoGruuaLEarRZalQi5JbeRvimWy2Qxg10Sw+xQXVgtx5JN+rcL
3ZBCE0btfiPBPyS/a6vWrPbC83Qbr3wmpkYWgD4zEUxGxsOfMddjTq3JKtekjAUT
PKevIowpqQPrrjgFT7stzyljbVhDJNGkC1SAHyFWu70EoxSFJCb81u/NHlqKf/L7
RrBnYWswOpehuLkttfa4bdYQKhR2HjHgLrAZRlHT4Z/51qTd7Ke2xGGbI+8gnglt
Nb3dCH/jLclrxJ9D21buqnnThULJPsqz31T+1h5qYSY+NQGfibfJ4WZUoA+MXKwb
XeGF+ASYEY8g0pHn7KyeSMMVXcGKi4qBodV5p0UEjX/fV6J7YQ+oUqDB/wHohfZH
sWpWObye58ISxfTRuEogKsmBf6SIgiEZfu6vVAw7nO49bFsB82RhhEz3I//iVvI1
8st1GLSf31J214PIzCCpIxLRhNN83xK8SlBel9kNELw69GbO8rxRjcPVaQKQEzm0
UWmggO838WgeUkbK73DJYrcuKHh3BBn+64F4Nlmo9QTqWFINB3vaIICzR6zswcUx
oLIfTIhVu9TaFypa05O6mwl1pOWBxbbclUYJ4uDng5uvkIJqIcD6CB4AuLg4QkSr
21khgoR13WHjNFBRFPnI3Z+6AiRn1toqtJsJyoMUx9KFmCq6KFh633IDDSdbH7NF
dnz9Zkwv2aUIiOEr/le395cTHPLfsiMWdwmAawOO4HRCPtd+z7k2ykaBbfLE54Vy
xOlEO7t3tXkvFsCBD357BbGif11Cmf+0mdM4CsEeaEYm9eXFzkJRGeRFj/tzx2Cr
rI/RT+Eljw97D3aMINCj4Las4kg6wNyrmXWQU04e5fa0gbbZxBtJOEUtGA1IjoRp
0hFUlz0CCPaZ1NPp1sYtCHEiXzAzyvdNAf0lEVgGh7ElgLFMbxipSM0mr9g33Zgn
RU35rGlXCC0LwWuNpapd6M/ffNXDk3lJacnWBjQQRuw/vyKqHAZFWV8cdkw5D0tt
5E1yI4TNY1/l3Q5xsDJJB5nwjF0AEqys/QU7mjjOlzx7AGSAUAmo4vcwrh+TzER5
vTnsRh5N68gLL9lOWvdHKM8sZsSmQsg9QEIHUD1fzgZijJoVzO0A4b8Gj1CY4T8S
Y8+TJp+ENY/NVUoTUnFyv4tvdfVfmSZHV+RFDy+HokCRVSuEX6QhPSLHUUnB9X7L
xf0G2og9XRbJ/fyon1W/MYGjXuau9Ccdhqo8w5MBhAGe1l9LLx6G08wRamPpqVLr
Shs/iLMZGBnMa/NKRsgOA420Da1qK6YdhBbSsztDkp0sZk/22FTXc2osPqCrmB8x
9cbwvyMIJwNhFU+aLInKrShj/pA6ilcqNvhSh1CELpQQ6EShb8QD62EgqXmKWeWg
jZzXeCfjQv1aR0xUJgeEVC/ElRDSXzy8wX/IKSCc7xZwGSJSitXeetEtQcj1aUaJ
DULuQ44zNtmuOiq/Da9ijykrTi43L/ykGVuSEd0IeFF1qN7u7HUFKtF0LCv9N6sV
9rzlUufIELSHc2j1K4XDn2CRzZOe87oTTKUXNA32jzTyNS77OixAMiH4sZcajZbF
U8S2IBZss1pRZA5pXh4Qv9mn3JHVKRXQo/1FsA2p8HC7VtTBvmhkMtxbFec1kyxm
L/k3rSlWSoVtFtxZYJZrJyvGpRESR+B8RQR+AF6u+WFGoRYhVK4FuvvFMAm8kiTP
4qGpgK+dPeuT8q9hY8wTugV/Ryjlzf9BnAeYHso+RXWUYZuzbN8OGnPIgSdQN1ie
1wsadGWm/yvbMqvKRW5bnbjTowLtrX3kLbJDST8AHcxsP55BsoaDoCvaLkALY+K7
DcJzMovb3ry+HRcWo0czxIFL1YN6ZCjMKRtdUiCh0ZRPBkh3X/GLLUUHRn0kSjfM
hCSBSawClHA1v3DQ1R/zuY/pDkHdFBl/8Jx2VFKrBvSYpQnhAUE8wDynMsOwW05E
vtfqBE02BoMgXr1YyjIUDzmmcAWuo73jVdhmwIBr6c3Xo+q+9YB3/WL0seQf90tE
tRhDXYUjpiVieqf4HPbBhgVLFzQw0HrNMw5NmUwJlA8DRg6dZuln6FgpzH6HzQIw
4r9BOCQXzku+Dtvmnj9loH2D73nBQlYuFBQg2jQxFFLUiGHW6da5h8+x/Hcj1HNU
59aUvn0ROQeXS7i54G55ayYf4g4ppVbdIWCowEMh738Eumjkd348ZcPKrlkLTLUv
WmMggZfOa32ikU0assq9XVOaJcIl1qD96Hw/8RjVTEyEhUlBHPS3HH91JLEsXbfJ
FdzeSx4GnWfDawAkMS1hMbD+Ha4LQvymQ8bYXzJOTcCuaJDYnHhcq4ks5ZqT/VM3
Q96Wig0ytZIbpXLV8DvXGziuw/qzflNJ6g24JbVDlRp1YWod4UiRfB8lUIpz3S12
yxQRkHqrtm4ShbsM4LuQZ1oS/Z77ZTW7kftJLtCvMQ19mz0/OfLFW1XOqG4ajXJT
jwLgeo6zZsTFO42amhpRFFEb98Pd8JaUnYtOCdf7L6KeibNuHukYPQCZu/RUNhOh
OsTeEFpg0qolL1VVlZG4YhWmqKeWkWcarCDPa8gS9ysPheETKAxLKm6wLZCTGtAj
9jtteLb9731Z87o/ISUKgKUZEH45k5KsmqW+jZedRBGoXC8egm+R3BMgCc7wwEj7
5AVOwd1/nxunk71jhnC2BA2zTWxR4OKP/pOMGZYPlFMrBm4935mT9O7+8oOq0O4V
vOjDjZc7BJQkOcAIDQ6N23hDjoIn3ved2Vow16fkqXXRunLXsvUD2VkC7mhAcpfk
an/9cTCXrR8LZFTmNAYTtNSyjOjU7K3qidFfGiUOCnq5x8kZVK9wm5I44Gr6WKoK
ICtj5tC0VIPscGi/Ugh6gUWS12OZXUhVs+7k9txAXcehRqi2/8gtsphI+Earn7El
OEIL2l+3y34m10HRht7D87p+TvlzNM87cLEfC7dm/Ksl3uHdffds2EN5mSXfzenq
AqupRpXMLDcwIlIayIWfE+RgliGpJfBDnArnsC/i3d6nwgs0yV6tW8oWiINM3767
b5xkM1NciR1+LqTh60ElhbQv8XKH6neCIqpoiZrxQmFQrmWdFFf82ywjgFMTmHCx
aC4FoepE998ADB51t2QQLAE0eN62AMYzVqK6Sm1vTVuqkwml+OQYCO0F9dX9OIwz
sQTsmQ32/OZMbEDeQVosS/T/hBF73ZATp2L4mPcqtVIyn+4AYHIBKeDxYGPSqu19
wUfjhoQTdIUJAR0i8bZvBnzV6/hit0Cx3E31NARCMQkizTd4mPvl1WK8ptnSzoev
8vyG49aM0whOyYYxSFHNOqjr+MVYZuZlcs1rMfW/Kni6OBUizgBAxrcwxrpplLLU
I09/J0B5coaSWaf8F7do9L79Pp7jTWhpXVSuJGOHC/pUKaPV5tHB/lWCqKXGdvQO
JkRuQP0QU1oJIFsac3NFcbqjeKphfEShrddqiTCYPY8BGshRFi+TrEvxqadgqiTG
bo1wM+7t6V/acJSprLIJWdPQ7kODq5mAUs7CRr08ECljYrH2TPJXIt10Hc+9M/rf
PA0SL8xO8rOtAoCZMBYYPAoYcUqAR49g4VEN936lutafE6cGnWKfV0Ut0xUsOt3n
0ZCpcxTBLN+j9vz+FWc4NL2TptuWCf89yyh1HGgG3PIRJg+7k8ujRwW5ymy2NcQ+
4RIijXKAH251EVlXc9wvFpYSv+WKVJ1qecgu1Uibyrcp5MMQUmp/YbM3lE9cQ9X6
87u8JJ23/+oEDTGw+TpHyyC1mnj8rz1u794dCIhqGi/hildT7kC0aY2jhYXwphje
6S6rOdJ+rNwdOyzGWvAR/NX0eFBlj5bBQGIFIHbI+YxhJn/4+ewQACuRK+JlmKsX
y4Q02J4VDUKhvxiyYRppatW3/Si/kG2R5OHKiSkOyYvhV98oWNxXSKMCT0Q4J68R
Z36xVrXb6jEe5Uwo+/W0XBozUmQmWKPp8orNV7JSP4idAE6iGCyLGNxxfr0WDWXM
z70sn2cXZRAv6BRKhrAl9FsKWf7w2+1b2U+VYf05mVCcEr+picLlaKj1DGg/CTy5
44lvwcq3pZrvDQ/2h1UYV9x+axKWxYLWlHbBoNFsxwribEYrg+WJG+tZ5LjPlWYl
/gMaFJV2hZiOIkKYU4J563zGcPPv9iJFjqpbA7bm0A/Ytj3PXkh9MwwJArsVBtpm
sVSNQjOhF/uZ2jSG+aE/h6fZfVQVIuff2a/wW+9RXWygagI5hC5vAdMLIusDbEzf
VZxtFwbO2zFzVe6aXhnCbuOpAyK7O2pu8ATgoRGE6p33RHQck84HiPo3OcHZz9DK
+m7mLmXebDm0EshOQtHjL2g9fomuy+Lj+M3cqmNTGUZcrWdxPrJyIo7Gwr2fyShK
TQe4qFGRZBnzH5w6d/4EBifNbDo76H+lMkBy7AqOelsKWXY2s6CchlmI2nuTEX83
vCQrS4C2J9c2RWH5k/4B3QjDBTCR54tNJVCRcYUcoZ3t0+twdceVTSl1jKgI7W8K
jjW3Thfjlp0zsadQxTvaHc1ZtBtwRLk6qyc1/d2iH49BmUldaCefdjs0FWjrnz8m
XB5QNM5u/adirzxSKon+g1pHax2iHDRPg1OxKkEEsKi7QAkZUZWihKocFFOM54zi
fIUSRDGsnHbLaZjydSV2chdub6p7nrvSLMqpsOyR7DdHbSayeoO4bPWBUJAhbSII
K5GKkBc5WpqI222RWb2U6EpYJkwgjj4z+RWF85KExYKyULEOGeyEHaxl5wrpG418
3xy3PtpVDmv5UYAwuHc5hjXyV0qwgcpV5H+bh6fo8VuMV4DMJLkXBTaTR1TQU37l
gnnSEwGkGfK84RSWf16rlnI/ljo1sEPTEJam46ZYdJQNd9lSW38y2hbJLCV5nqSv
a/sL3icU7FcgVqcjdZ8onkc+kNGUlbexdMsTlLmeaAs+R/nayOMgFiXg0Ukwk+ho
cSac+wZj6ylictlQU0vO+HYfBVibY+IQVAgiDyvT2WuTVYkLdlEwU4iWGkcNkazg
S2PIaZq9LoW+d3FpxCN8t626HlW3LKDaLUJ9QLEByuVHCSbsKh9p0mFG1LQPuFIw
lDyoIc12seYPwWk7+FwowIceiq5JapZ28Xkuxz/uS09W2J+NuzfQXWbPslvUeyXS
niSJfXho+cEm8/yDTEGh2l+ICID/22pXylEird6hac4tsegGJ+l/rTWm9PxInJrF
X/Hf5vM0hmvbw8osYB65oK7pvEbaJbnOH2INF80XcztWVyxg8MiHegAcUxh9kjFn
M9YwqY4Z1az/If3Ueu8BnAy4TzX9q2kKRs4r61WOk0GX0FIwI2BCmTC9Z2tFgbkq
9nVWHOZggqdwt/0adyEcbIrmZW6GfpZDhwlTAuJnaGTGTY49mCNYf+O0XxNAUBNC
wKVYu70MS24Db90aISP1WEODyT6sqsC8Ctl08PNdkge+1v69WWVu8B3pWAywcvh9
ggyGpmU8AEh4s33ByQUJromAh503aEYlQhYLONwkmEsBwDtBN/66MJn1OQtd9k+v
dNBwlJTLAG95fEHFPQHgk16Ae8Pni31LnfM/DZtXbEdGqN0YfR3qr/mabsLtGR7r
hy6Ka1EaxWZtFKENfNCau3OvLMdG3flcJuRQSDwCEmXDRKELIPjMELYOy0wcWzCj
s29qWlQoqpRosnxLHWnp1dSMEiXkydvat3fXU8j77hfbBK3py/SWe11apxoc10pi
UMlNYBQhtnLsSvIJOfZY9pu0ei+O0Bvizok7aXRLsmt9AAUFLKbmYsRxa4z/JMlK
a06DoWF6wSSVCVHo2miNfv9KInBAM5FQN3kcXVNCFKBDNaNv0yVUWf4+509XzxwN
I8sP/M0hbQPbaMPjbnsZ/9q/vP+DleVcjQ7xthdrV9/xI2iYi0ENtQ5ORwYezVYM
TEzFvvH5h+TMJJ1aO0izRQHUZSUAgUzVre7ehVhjzBYzCUh7CGFYVaZn0KX8S+IC
VFxbbbwOqazK2q0JckCXXjRL2mtjE+rfa+zEkJAo1isjqXubN1Iur6LUX6ARBS3w
waEcaOfIOx0KugbPwyBy80lbrTtR8g9PDq0pQdYmFvsbgqddop1TII8fdEYkgpn7
QXg2E+UgvRpdPX6JAUkopp2bVYtRcX1wNWjiCBSUUa3BmgrSJLiabFwFQdwS9fgk
Ap6nRcDxtx/1oqNHh/QOAhGraOAjBub1kkkkSONqzIGErvfzBuRZlyO/L3req424
EEY3/5OZw37boZK9fpu07uvwdERIFfUmq99w1oDHBfM0f5ni2ncN6z+8GFIKqtfJ
2/cgt2ifZz6nqMhnKinXI8yO830djbyDYnG6r9R4vMI8B2f1B6133RaIpS8bjvom
pVazXgrZY673bSBvTBegRpIedZeyiNOqy+6HDYr24QR+dfs+IixAu/sx2877Ir50
R/qPwLK515oUaap42l5hMG5ZjRartzouZ4NJJS5HLaMsU3qUyCwUrF/YgAc6nsS4
TuA0FHsRDMVn0K4GmhwZ3sCrq8AIgE22nIhiJbEuNQ28xP53xpuNIZlOT0ZLwijl
7pAqmAQ3t03PCiMzKrtl2kJ7d7s5pk79kK2yBEZM+FvT+S8tW0RxmkeCUyKJkexX
A3WQZvPkAedcT/1uIPeipjAX2Kad6vjjd+XC9TFFzWwrHuOnXf7wv5ixwvkOdRx2
fdCVhtq82Sp2UfM5AUjGhPtgAsr1wThfXMCdYT+LP6dDGCa3HW+d7O+dDQ6sEJQf
9Yh9x5whUWmafLXG1QdKpYWJyNvQUumkdgTRklXgb2IdC9pLGC630C12ue1aCYCQ
pole6g74hH4QQCnb5w1y9ZqGmRMex7BJEomf6LNx8Yyy20BXAoZXETWzzEhBFmgx
N4NR/G8h7b1zTxJYarc8GjviAHyH38vZUTNfly92/ijsX+RoXDiOTtaIRmF7vvTQ
xE5oXokKqpsQ4e9HU21epVyp1f08f8Se1ukzFaUOhPRrO8QHNrAnFfdQHEOWIGBY
`protect END_PROTECTED
