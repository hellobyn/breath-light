`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xb97R2Fb3kgaq4eg7WcXp5zGFpP0abIzfTxPsaPX3/OpZb4sg0rZLhKVUMg3TQt5
CemV8rvUrbnTaUiD552LU5OLspi6p66NF0FiJqegYyHMgGgPp6LE8S3bbRF/LTqA
Y8/OZ9aD8L5p80pOvs9ceMgpZ4iamBIZvHn0qa+WZsIN3WpClloxoyAErC9Muf6h
yCdIC6cnyep/5sM4Py0wbxV8IwXbEvJLH8wGfr9+SWa5VHygd++0ypZWYH69cRU2
GVLDVJKcKcltyIT/2loc20podrTrtbXvB6dhZySYU1bzRu9G3aIOja2hTr3bcZSd
G2nLJuvyRVRO/B1/ZuNEm91SdaGklBcbj1HtNW2WUsUSGmQDc/AK6UEMaGSTHohx
Dv2F4R6lI5RmKuEcO9m6Atk7m7TQba1HW0rNkcpFxSCInBZ3U76elADwDysOvpQM
TRjuokN1pTEA+F1hdus7cWTUfCEmLmd+cXc3RFx1jLPjm35VwwLa7wgWsNas6N81
i9rc42VMqOrYCX1neFtDBSfxDp8ci8tyiPUUiCf5QzZagYDYrKrGwxvEx2U/7YBU
Dkxs8aehJt9GQ4ItVAYgiUPc2enpsMuiagXr1sEfc9/U45ggkiCCuZcregVd7B8N
01Z/z/uobzc9l6KljwoLIPRwwcsejH56ilPJdGq+kPsai7FTHQLOeWPhAYaF/boR
83Q1tWJcWml3OL8RU9ouefrbwTwokpTo6nAlYm7giGWRWpEeotid9kyD21H6cJ2y
86Q9k4ph6mO8jcFoGkPZ+CcQSc7hOBnw4PtZgXhrzMOCEzeAucqyVnkgaNKFqgUT
sBvAECBIEtJxXcbsrB9+ctGND8PaLdo2I2ID3n0A0HVnj8brUo0zKHhFhTC8AegH
3bNn2yohWVTO0LHWVzRqf3Q2wWDGMbGSuNQDC3X0SPfW7ewRyOLEknN1MZMeElF3
`protect END_PROTECTED
