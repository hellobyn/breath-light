`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUNZv09JNTaqaaXE/mXrowqBkJpp4fvkUZzAynC8A+VYOUEl8EdWN0pVQjZ7rD/u
tf51UGvaz10uQWueTeUSSTizvZdzoOKPXPX9DB1HICO+Nre05GBy0Sb1H9mpLT/p
qj7/US2aRdyacTmBrQpETEejtsaqSugQe644jcMgfJsHaf7GZF2cGqhuvc51QiXV
zcal7koKHKLixrKOmmeFffACGgoQo3BpjnU+QLe49V6qLS8holCqb4CfkmxNk9S3
qNeO5eEVOl3tZHpmqyN0d0OYYSElnHAbk9yJqr19S5oKDzUm72287eTqTRZsP8Fw
pGZ9H5U88ygx6/Jud7Efs5vnv3oB7BnYMnOg9bInH/C1J8Ws+s4UyZPBZX1TeU1Z
i5+kUNXcGyocZUu7zYUTA2cS7s6JCNDXN0REEdp0hlmnghhFIankeL+llK2HV1/5
ptQhJcJa3Xd2SKv76gh20p4Fl0j3zyfV7d6tx6yx7P0bKwMJIowNks2dK3VyMbEa
sCJ0E1JPXwBDdklFiicrRd+/+guqWfgikTGmt19FfVXIhaIDJlF4Pz+jgJWK4UAy
nFW0r1JLmkkIGS3QTPuOPiM/dkzItiBqEumtXtrNE6j8AUJG/bDkDs2S55ufou5I
QWmitqEY394C1XQUC8yePSn0Sr/Ea7mBpPNT0l832p5EzmcM4tVu3d+/fkpCe4+z
uMq2Y4k5m4iCn9u6DmVFjJ9r4G3OwO7lT4JgvS6AbydfCJirmWlBSWMS59wwXx66
XWr+p4GuWGlEaUbclUxrcg==
`protect END_PROTECTED
