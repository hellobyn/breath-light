`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNc/xMq9kFd/fRRXpHLP5U5hmYBVWvL3XfWXwXRUDWSvsBZ2ptYgMOc9d4Ynz6k8
PSXlKxe1ykY6dSTQdXexOLOwF2WJChypnBKi2orusFenjPh7xdms4l08cHcPAblG
J+10XMFFm+exFh1MttQW2/Lgl7w/3GN19nA/H3MIoF7JDOi8HHUo8FdLAS3mU4RS
BvI37Kxmp/dir3Cb2GoLMzkCHBqYvKdYvuUk9TIFGbqvFOO/V/pzJGFjl10WKqOw
J+CuL33S7q9f+Lp6+5alBoM1FisZnkKIDniDdA3w6+S9wxPSdmDdyBD1Cg3/yXf7
RnBiLc15YCE3c2733+etXkjp34hI0zEIwDWy7sdfa1BOIpg0nY6SG7reurrwqNnF
TWX5oEofQV1T2EFNMqCN/uhMs365zSyT1lyUSTme8toi2MbCgW6ua5wmbdP6AGVA
8YU3APM3eujk42U4gHcaZdH+Rum1FB7SFfprSNWIyQCV5tqqItcn/7mPg50w/LlZ
/h5QDy+bAFjQoaYc31M2kdTtCBEDZYjXGTqcAw6dJpdFb/Zgyb6V+KGRzIhtHZ1r
Jw/bCFAnVCRz/Pf6LkpagOdQPqHyQHZNm0ocOWmADLlQoPS+hHS2WIACzUs5Tlny
N0cI9EsgEoqQi6oHSFfmunKn+nkuQkd8Ly9pTB+BCyu3o2ESdlwY8F49+depTHca
woIfz2WNNh/ynBYfPSL5M6corm+9kdu1BPGjJsFjmRS5NJCNWupCqUtnNlIN3i2c
0G/PTLKgfKaDm7FvgRzl4VTmeVsOg0UgJJrynBrBRJlUnrnvJlhpHomVaazIhWJf
h/zePhY8E30BOmvYEnWe1LMMKM4/ppXplAmkOdnaW9bnicbkDZ2wOFNg2hscT3t5
Q7QazcH51VdrACJx5bAyRut6OktimzyblQtErNvSznUwD5Yoj7jF0NEsaES+2hlr
l0yQXG2DNB7MGyVnnmWOtyTT7g9LXG91N4miVH1Wwqddsllx6Sac8YW15hXm5e5d
OuLlHRir1X9OXOTYnYjwVmwGlgPwaVd7BbujIV3pWPnp3CQlOCZgDff0E03ue48D
PT9quYpcvMMBPrVWBqMq2c1x5SymwzYQNUK7bvXxbTmZjKBthQz/zbzwnqSxKQIh
kYyc6F5/Abk1HO0waunIWyf1izy1/YJuf7VxpwDkeqQfj63FH+uP8cC5i8cBUVEg
oec0v3fQUMtrI6wHs8clDy6SG7+sKLhcplO6rSaZjxM0yu0g41U3f+AumuJPKs/g
4LVc2QciYDB8XFn6mKZRoGOIhcwBfosALOjLM/Fvzb/XQuvJWObdg2B4kSsAla7N
Z8azlCf7sbpSVsfkY5NiUKvP1C3MGbbnhVFIXAQxOrBLht4ocZrhLnYMRIFhpK0s
t23f+cnm8RjQOH0ZfUu3H5gNgYk1165irsH/m41jVeW2q20C9lCd4zkP4wu4CzMw
tfLzTUfuhUisMwyr0mEnvS2L2HvkWYprXKFbHzYFQTZeQ/0C+8jYHgKf+YddQvYn
Z/G7k8dlGFnaMTdrs5XwPoTVo2MGoZUbT6zKihSuShbqnGiCMSbzlvfReSOMQMiG
pFqbXQby0aXnPtQS8Gek897ijjxjaCWgZXxr8S2EPQPtpNdLT2zDrmpWm8EmsVAZ
Cpi/MLsJkVfI43DVa1gGaFAq4i5VwWexKFeA8h/hOPYgKf1B76CVvWaiOBcdHDbv
rvn3KB5wp8JitXc0B1hp21KxRMloKa/QYKkSXIzlGPHPIz7Z3lXhyOokN1zlW9Tu
4qF/CuxQqXcEYSzYUWAiauh92/ktSzGuRz++AgdD2JAHqgo6ArFsHIMR97u/S2l6
KoSMOQwZRDd2VTE+7fRS86ARhL5fjO5I4diYjy1/wvAzUw2Im+2l2TuqMZ0SX8jQ
AJouf4vivF7tfjY4ugcdFB0HdLzVNYM9ZEM5xDi1fIw0kh5rgmiVi2dQTUbTXF9z
6x1w2EkJnyRgcoGLyAgVjhhxyWKCWPIUo34mBXjyG40/5/Jt+LEQ9PwdWaSjfpiK
UepGVjj69gky7GuG+MzqCLTcjZGpYZ1LU1GNx5CkrzeLzsCtQyOprchGeNdBt1j5
bA05imM67rZTeCGJ0RYTcn+fQQrHvU5coDZjEabRX+r5pyU+dv0pfiRJX5e8PZ1x
OOQogvappVZOLNKI/H6KbkSMZXJBBgztjRnss35Ych2n9krv9QJOIr6kNLasbpZF
Yn66d2NCWXQECkDY+aIDj0B02xXW8gjr24MQclN1XLKS3W5xfdWM4Iq9YpmnU6qu
tJfd56ZiRxGuEVt86htnsFXMHW5NWJT/4y3Csxt57/Wj6TBP19R8tEqKhCEa7jnn
bPEk9e/25SZ7MuGOMONZYTBRm6jxRzVfSv432iwdDhIFwSZaOIZaU6m+HWdG+ekK
RMUASCzTek/LF5iJ7Qrhlo5n6APi+iGpYbz4fb/IEvWxDZndbsuFEO7LkSnZGwhZ
i33a7mOSifkzN1zimZ9vQpwIQKh+eEyGAMJKZmvWG/rrVWkEVf003zFxaNtZu/nY
BRzbUhr/HZNoWfcPRrp4kUdppCMPQ55E5J8D+712cmLimHxTrQXmHB8bdfbz0DzB
cdw2p2fz8IpCJKe/nGhogXTcJUxv1+1wtO47pjCKCmHv7TZom6/kauKyS6VOA5bq
oxY26k9WqxAlP5Qo9qC75aaZSXPaRROVcqILcc738w43J5eKCFuSkMZy6H8dja3L
14APPjgRO0ZE4ZCUQVL5L1nL5162ohR9QE94ETv1kI4mPTOaxt0iC4FgczNL5sCs
yoCVbvd8/iDGDOMprlBjjx7Ztn8VD9veLzXOXPBkE4d3++vt5YPCUr4d9PluEZ/f
gtzWxSpNNMOMnTO1e42+mqL+uHum51yY8JxN5HP6TVoNhOXcrRR5wGoaWgA3oBJW
voyvrTFBEDy/6vgponHGG4FjgOIKVtciHGfUWIRmVleMhYEV5Dp5vc5Paf3l199y
ilVDS3xBzD08jrmC0epf3osAgkjgsMYVDB8YYIg7LxG6T1/VJniesnHFa06hysgX
qH+hIxZ85/f2LtKCFEQexItiNgFuJg5ad2PJs2zUQ3QwGhXmy+0SG357OWHvCW/r
fwtTfjXaOM6dOeozr23M5durKnF3OD55/tv+4aMzP26H3DJeStkaIgdM4p9KdwLn
ngg0PMmJ3OLfErxVMC4CpKThIDZUc0HdSaGeOjlVLerel2tksDYuQM4wiFj+hQdc
KTUQpcab/kd64RKJzkZPMUYrDZips2zv/6WolaPQIW8ak0iIcdh6oANTOGicGW6d
2I6fq6klqFdogUFszwqVnaC1vAX8QAw2y972xelYVgCBo7PuvcDuEqfVc+bs3buF
DPPO/B7C54erGZPX6J92W1rsoQxvaWPOsWUqn9usxW/kcFhH0+6pXEnOq4BdcuCT
JzdbsToIyWaOpBDlRqG6YD/89JyFAuZl3OM32tk5VFeQABztCIqqVy7obHSB5t9g
`protect END_PROTECTED
