`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FatoOS/5pLRseFkd5KB2ndF/zT1ujLuGHKRndefwU0gZJskBRSN28yqozTnkYgkj
myR4jXpm3skZsp7vayZcFUbSPpWfCQlnxU6OHOSWOTBnLUHHPZYjzASuGCYsqMel
uaww9H5/l13vApl3hgXUA8dE08U1Ywq1zF6ikxT2zAD/VVayoc93LSC7KWXSwwX5
90ymYJgjolF+2GQPwbRKVCtRBD3+YB8HqX1Lcrjr19skK0UGY6kckjGlc2ly6Xjo
EbuAzrQhD6HKId8BDmNGTNgUGZx+fGTQjGdbMJHDdz10klIrJnWanBdbUza7hELg
eND0MPv01iCZZOdetomX0xzlSazplOGwGPp80YuUZhUHcYT8PhUncARwEOhO1SSu
V393m0DKWv2j9UGnofIxxDKix5SgVUxhUtL+ndMN3o8kLg5lU64kRnQ85zhsJgmB
b7PWeoEJrXJv+7yUY1h5TCw6RFvfAYg0dpAcNJlqbK+Tva42WOVQczciUYhBmk1B
q/bfob++iu9kpFBOKzv2OpjqbIoWOIgjePlRNFvfHDs=
`protect END_PROTECTED
