`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JSslrHtK6wzb+YZAjMEatXCp9KBft7QY9U/iDykuf0nqk9RVWwSnl5Ii2OvTQEpx
E1VYlLoAjM4oAuOomrZFAjtpgt15JjRlwMvEuoljx9JpaHjjkASmSQ4W+L7OnORU
snWQ98TrxDisF9FYKsGcPbteVkIeqI6pkABPuNiNojRRWL6n5+SFLg5D44UPbNQf
NIvfRQz1CdVYlndzq+nLRgrJZaudToLUdHWTnpUusMO+1tXMPlWiKbS9ONl14oh6
Au5JCoq84y71X6tYN0RZWVtTnEQ0w221Gaw/GMxbUjgTnUG8lCiuBOZwAj6Ijrbf
/XVmNq8vfsmMrqpNaxywm42B7PprPd9YOr0wFe3KyaNsMCvr1tFidwVPd/iS99TI
ae03AU+0B/ZLHljIXFZvamKRIGOFN/Sg+INcK6zg3fWOznKZveuWGl0uvv/nQAIl
mmvacRucjHxJPmC/COz1rhqTc9UUIe0EiO0OmOodaN/qLpPCDwyA2metxS+dijxR
aFmilIgHV7DG1u/e2BJMQJYgG9Y61Sky8wnZlb4WfT4epN3BlYtbT+sWskMaoh+7
F5hRTwMCkO9rNqO3uMWTtpMT099mb8cct70wxWxEgAahDFnKztksWPcS4LqK3LJO
kGNh0LEk5tYcq6ify1g+Ukn6iEXWUwU74hMnJhlhhqNWeEwH90i0KDk28gcs0LyI
6tp8nRLz7DGk1IdMmptizaf/itqggnVfS5tC+OJJJwcNN/ls2zLd6/SRRqwWUkYQ
OqDbt1alqlmlpeu2lFkCi1t6zFAFIX8lgw6ZJ1Iqyf6RH1kybftrQ7sjKF1t1B5E
J2ugoCl5IlP2y09pTuGZQWAbnIf2Wkllv+pZn9J47Xu8cRQp5a2rhmhh6CabrXXm
TBK4TWzUwk3TG6YOOsSv8aXEPO/zRw0moxmNGA6G2OPZTpx6Y0IuCGlG0R8sulJF
nUfnleO4W6BN3wGF8XL4yJxaeHkf68PD/muSBeyS6lalDjt0GUtpzVMW7xtVZfE6
nRvjgKWOUfz4U6KfwqiwOnYQHWkvy6U9nPcn2JAFHKi+o9LtEktzXddYir3MvYxL
IS1BQF3nKc1QHhfqzTHPAZSgWwW4sP19Rgs/Wmg4S7hPWyuyGS3G0tDmtVbsD9du
cpvOXQUizJZEzYW0V7kaKXFSdnmlvpth4vXDneesgHocEFq5FA0PFvjjvEGZ+TlA
uhXnrqoeJFtvSz0+9Lm32DzmwxvvHE57I7SjvBqyYXSf7Fcvlswod55r0GLl/HYU
g5KzaCixrbSVKAxgTYe3j9DZP4Px4POeaCNhICPKir1rADDr6uzzlOcRtIUuBNM6
mL+3h76hqaCorzfhIaBaRwDFBuODSflIOzaTQQAErHSfEDEAbvUnNX5205Edf2Vo
PKzczA7bE1XaqSpY5JZAZ93zJUS4iBukjuRT6pqcb4wW7P3eyqDRTbxapvou55Md
6qwkGpSENHIIQj13SQY2SEbPStRYASyv81IY32/lXWeTVRZCXSCEzGxn7jx+3nDs
LW7uUR6r+fIXDJTGYXJbhP3Hyx2DlmB+9awSE9DF6yDXWRAjI9cid2vIgezSR3+K
W45dJwRm6ed5xatCOLAgE/WnvWH6hMvBKa0ITu4F/nK39p4sngHk2mrAQz8Dmori
QLxRLMON1+s2ZaqCc205dxgm+1gvR2ObMv5Pea5SPB6VN/1bEhPwYUSe5kXEhwIE
qcDmlLnoMugnItUiliqUahSJy00smbWYUnHrltHcTOH7u2L8ofM7mf/zMpry22yj
e7f4wr1MZ3dhg0IZKHu5ezDCVWphGAM2Kj4JszUtr/rkOjbc+VtMiKUyD0s3YnJ7
6CqZXEW9EHqDylsyIsTe6dIkW/QUvk66xTwy4m9ZAg+RS9YDJXIKHwbFlstZKwKU
/n3KodpGzHx2W9wzQfVQgGofvP50V1gItrPYxDLB8SfA0e/L97ku7k4+fAXRN3zy
qclXNXOIiQVZk8lpMk6MVGQNF2TyKpOSS45fjIARSz49o2xNVjEb1tyQV8iJNQUe
vDF+xyA5KBlXXVVWjoCU/Dr1qmY949M57yfAtttfwhK3SqiV5xq2+Wk1rLf4yqhF
yqxOUMaeAt73dtFcFOhK4IZ8B6a/b49NfBYKfLiUkHYWLBqnqc6QM3Mx9D9Wjz6c
6JFjXa5b24mrDL8MDkqzZTeC5/TX6yyXNnoQn/Y4BGXO6mLkK0K6vBAuIYcdHhSj
/qbvn6X2K9yRXoNgIhg4gXVBuozozRQDiak6IfGmv3CGjhTAxS+MFpN2lVaxyp49
QeA7ia/zNdZCfK2A2HKaGDYMPaxdelEFpPz257HRVsDN1UGcvzkwtiLT9CLm0Wbl
1snvJwTkCQVPjHM70F13jkY6hH4zZZYTcN94rRA772qc+58EYganvIoFS1HrUkZR
G6AgRmi2rRxBqsV0mQlpb5ZrJJQYudLNKicBXlwi1ltI+sgBMNZ0/LJI9PTWrnBS
y1mlr2wYUUaUworDHX465+Rjk/yYZXXcKCogEO6ZlTwtc6rd0RybaG1vvKJI4acG
JNEi4lGMBdOfaMnByfNiyXYRyx24+ctQ1OmNwpe7CgGvxSS05EFC5gqzfPX8Q5Ln
ExKuk9pcRdY4UUh8NfmcBjWpufJ+zU+NxvCDbKEESaFL9q67tM/iQ6DALAb0O00Q
LOLHdolGBLRqQjL9VlDsa5KmdFKsXkHYi5zLmz77Jw2rANwPEf/NqoczdunPh9aP
m72GbHbZvfz2wAI2cZSeUwV54vpQZLafCQoy+pgldu783va6ZZHV1qEmpuxggXtB
Vmg+waisrMj5z0nMb5i2w9/grpKrHUiIp4j/HNMyHTth6pX/B+W3DMBxRPYpWwPo
IN1km7wkP5M/EdnpsQ/2d8KEVnz4YCqipflltiRnoIjXW/PXuxKhoep3AokpqSD/
Y8ss8KqdhSWpoJF8faNiGaRwdNClAtau9EgTGpT48WEiawFwZD9T1kpL5qrM7V1M
5hPt8p4Feuy5cQYq5AWHU4FGMuyM9ctyJFpfEcHjc9hxx0Gvgir8lme9H8CYyn7A
DlDJ3uhDXw0ntXb3nr2A0g3GiPwPmP/Rt5iBIk6GHG2k9MFnU3cp4U37sEyFYvGQ
SB+hYv4bhVDMqBrqJDpO00GtzIAKaKBjcxwhw6NsiJTOYGbvOS8zZQCwXNkOl/bQ
ytupgEIgTju0I65pzYqFELhFwNw/DQoDFD/PGUD486bjNdDX5kfJGc0fkI+WTWOd
h8yPPjFr2piP2iaMmB2FbE9V/1KB13Es3volJb30YdV+HcjCNbpKVM747pjjknJY
cl5SGDFZ1SSApn2Ud10niWFNdBmlVBLv3iJTLVY5ZOsdBW3MhSXlJ2AlSv/H9opz
DCOb5/uHPMvZOqxvfzCkV3k3quhbXnRf58YhvbgyMOVRZW7wUVcr5cQHpnsroAyd
R6Hb8d1ChtZcCf4D5jnuzJ0rUrm6rQktoHTribvwhDcrFLdik3Yfhsy3X3BAD6PA
3ycq+TRE/7CJhAFvBHjWcPTZMciFtT6d6b9JssR5iu3YLStrJoG7Aj8R4CN55COA
DEMSLqSAffesBNg7rgQV+uRphi4X89IAgJ4e5iRt6RWhT7CIKdk/Y5JX29sJqhko
symKYWDiCe+s2mBqIGJl1XKbSP1DdeG1HLJdvIRDKEtlXCRXTXsBOX3nXDwGumAW
aR7mTd3g7StkRepEHHfxjgfTQFHvGa3URMQ0RxsiUHrfQjX/fZ4KjkegNad0mohm
rpIebFbgBVZ+WD/5bZzxtJwA+K7dFZC6GtSpUpy/ltVPFaFUj13/jSLxmjBukkbz
sVOUh037WAH/3RefW4i9ZTMQoeMEB8AcC2C7Pu5VEwaEXzfqCGH0aUFrRCdYcX2R
hCjRw8KFi2F4zzv0u07GSdBV1KYynh6lJNxI8aQ87J1n7eaWfQ26uZikZ+tylkNO
DbnzmUXKQPTJ6LdBzjXS2L6Sa0kzGTbwGYVpC9OvyNoTXMecMdZmnEBW9s9pVNzE
Hx4irI4PL751xJ9QvRFypgnam/eqiPNsBM7nmhUVtaVRRkHh0x45cbuKdRd/+nIG
R3ZoXbgVJBNMVpEaR7ItHHxlu789PyylBr3nBFqeXbTe7IdJJce3kz15+iqmHkVN
owY79nI+X1a+xJLDvUcCFxXGaR5UwB2xRtDScR0qdzeN5iWB2q5rL0HCasl3WHn8
zx6gxyHn2yaPULGwLQHoNvq6WVBgS9ve1fRBw45Cz4dN43mEX1GbhFwaZ6f5N/2K
Gzc21aFxk6+Q7Y9Ts4pfrqOnVeIYPf8Ucfaa4rE514y8DkV+X/ktFH7AxldGSgqu
AD7j5eIARnOAzrk5z9Vp7jHTQ/JtE+t1AhHRGYgG9KtrKwFw6qJzKS6AeyufY5U5
SOEvLp6IewStKS5fMQKCDx4HdFtmwGx0R3tLK/M6E8OJ+5fA0sYcOCLGZDA147i8
6qgUG92YSqWcVp8ewlCq9+j+YOGbXryMLP3l2B2vGIcD65clZRdCIFxZQJautuf1
yKdJHudmV15JCg3PUsOpssj0MEYDIUVHBLQaSHziUJkjdR0fOuoqQ+1oSuwg8QPF
KZoswYIRsOUnu3JIkj38c08n9CFJmFrvcw18HWkJoX0cXq0yWy0x3+AI8sqfDZt3
ZbKpOKQReXYrT0aBy7wLc8tV6RgLrNgTrHlJkNZkGfCA+6kvV6jhODFTxVNxOWD3
h2Mjq7Jhl3z1J4Q+heNkqiv4gq+FShgEg3j2VjgvLiT+rLmCKEMThp1O9cpbvOXL
Pr1OE8HxoPNAhtNkux7pvVwbW1XquiV4EqjrLnZ+HousUNXgPUuhRGw5Tztj1NJ8
TDgN1Xhh0r9vrfOHayTrIWu/X4wEIwdSwhWgRGOzV2xEmn888s3U30nEjyCv6aoU
7nDcBRnCjo5qcFCwPx11swObsZBYV959mWlHvZxWOP4axvcOFyTe+PTlGBad+5v3
HyU2j6BLqLbPRTUDpds8AkF+nR8ZVD//UcyeZxJfo9u5xag0DWbKtitEepB4LZFz
Bo0W8Wxuu+dcvZ2pN32MliMe6BAdDFBvadcjPFFcFVircHsbFHZ8xugi0EJWUW3X
ZMvJh5RACMzkBsBQAYGcZhbpEm2wANv+Nhc65tptqqIuE7TJbVTFhvBpqSXJNMjW
pUc/zQh0zPEEZHz8wC4VYJqHS7e56hYBy3TP/AIrDlapUWtrAMbZ3nmbLkHGumJZ
NpOE562irqSXBqW3NVIAFI8BDFEJPj22ajlw/w6IgJdbcPWLEhcEceL9FQBUtBZK
TJke0i1iP/HwxUIuqou824l7X54esbzY1WmqhoUx7qplrzfyHYWpcbhJ2eEZWnUh
GVD9cNFl3BhUrrmCvUntdTePTwbPfiEEgDtFqXLe269f549s2n+58mcthH3K/6kV
MtkxvD6hHBAAEjSkbJ4wcK9FWb1aF2a7WeC6AG/acN74Ny9e4AyW4e9mJatx+6Ov
czWALprCzVfNaMfiJhftbU5MsCZeFnT7JS+f/TuSErKuZAHZj8g93ThQrQtAFryl
yS+fX+h6ZKQXsXbSTRHLX3bIBwdyLpPdUtcHrMEETOeNJ+XO3IRTCwkQ5BTcJ14+
kRtb/eT8R7jrFHVQLG+Gk5c9Yzvs/7ouFRBB7Tn8cz7Qc4f37P2zUuTCl0i0aEBX
Olijwu9tRi0fKngZMojpRZhM+oS+zl5dips7zxwtoQ1Ovb68dEZGqPNgzhST6u4J
dm4AHL7422+Dn8eX5PieUAfPBc2dhaqYMudb/p3eXI+kc9MrCKLlum5UKtqB5udt
l0k6D22tQTdwyAY62S4dnhgYCtyHyqUTmHfpJAVEyfM=
`protect END_PROTECTED
