`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNSOQWgvR/ceBrDeoSrVa/EyjzXEp5vjDyOQZM7PpRpYpuLvV9g2aY2rAOQXYUzF
XIDp4pvlVh0RduBN5+cg1jta5RwX+gaI/SP+8uHHlHzo97wOu+4x0rynxEwB1cwY
kVeFrhqhV6qG3JrQ4G2i2Oo2HZkQ1Lv2HJo9NkzE1qOnnmedbUfKLDyT6bnTO/dw
QSaGlgRzjKft9Ndh19tNPG052732v1ljuVEDwImkVrAw9/cYBKzCt7SbBbZZr83K
OsW33nkr2FAr7P+O2AoWcJazSgQWozzut84FEhM/lG5/FMa6FBp0ezsvi937FOyY
MEGztG+1xhXANR7LS14aoKxIJq4fhBIf3pt2o2fvVvKx1p/bFrjb8lC/6Cr4cNVf
yE/XGThFZJASvWWp13u+52hfYQtAsMsi2JzgMo4oc0wt1sg8ioEgk1Fx+yG2sVx/
JwSf2YkBziegT8jekvr2aVOqeU0umDdB0B55LAfVk2/mi9jkpPh+rhgrdeY+5Pun
dTau9MzDJLpxGdXYNwxuUyRRGHRt2WKH1IL5Q7uNL8FELquk0dHxP539MwVNkDob
oBh7b+n+M8e2zjFNKbVFQWnPuaPUO5dnec/bEAZicj3w9M03Jj6gjNVaOCzVNuK4
tYYP/ZTd5b9qqhOBYtw6ZDtuccAgHr9hl+TWBOXNPX16XiTDeqPfOahnYrZEsb8T
fsMY1QrvocqsuL4ofkzbYPdDsC6J0ppcMbL2EW4/bs3XiWOrsMqosMLcczu5/N3K
2fLto+yksstYGLk9+lUXXA==
`protect END_PROTECTED
