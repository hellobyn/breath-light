`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQRTQEF5Ro5mAK2Op31GyvEuq13VoBll84yZzQDdVJyviArhualLJ3b6zyzlypNw
vpqQaVnfgGnLM0cVUc+JyIdrlSUlzbmqx5A20u7m2IOkcXisSO6abolwS6NlRd7S
CjetxGv78esF28ZrIpCmvIE9T84c+mC0t6UKV3XM4oZIBrxs6Yo3q1/Ufa/Q/Dp4
Veqh+SRb6ocT4nYQV6Ry0Gnl/kwiahCwYHvEvOB5vG3Bb2RV6nRilbe9/C+SgtyE
qE2oalrl63h/k/qU6F82yoTdiq0GLifBmwE8E+/VadkvV3vzoLGtoguw1Q9FCr+P
SyQ5MsO49ZdbqyzJpUpGolontHcORVDyB11DRNGgCniAeOKpbh9J0bMTciaX8yCp
nlML2XjxxBKwSEiljdCCu+aUt9q6tX/rIzRQ5Pnp25y8bfHmOwmZeM8SAf0vdL59
JX+gmNFMQBsPRYyiHAWDGwdS7er+uQtkFTAjE6tVr+/udexVQoRtDDmVI8AUb51o
oZCgn5nIT6b1EvDF3ARpKU9pKebk9w9lgjPkOxrwXOuZn+NwV9RkXxLQ1/5n1ihk
6fk2RpqjXUyV8485K2MNoY7O3Fl20RiKONKOqxlqzT8Y1nDmfz7xww12DDMbsHCl
3s7f0Ga/R5rOkgCJbGVv6HpCxvZuortAZw5cPhremNDn7wrGLBoHqz3semvw3520
KgLajAX0nBPAwSNmFdVnxttBun3oRJx0fBNMVSbjXsVB09LLwokVHalYqrLaovp/
cP0fnutoT4QIp9OUBq8sexymna7bY6cLtnqUQzzLQ8f8FJbaFTVAsPClsGO1IZC/
AZdy5YQoC8ZFwXfydhvBpwHC+Rg87BN5eFH+0oo/1WjFuPj5NasZ9fk9mMzoLDZY
i5pno0Kx+U1/gRsL9/mh49cYYMYwCfsuhIceoAZ4isgLA+3DBUhPeY7iKZSbH1aN
cV54cefcvFXvnE4h0Fe0zQec3sgwu/zppLk5iClnF3g3bbiVHE1eJJpedDZjWKqG
oQhJ3wEh+1HH3hUjpjBf6rzXqGkDl6Q/HMw0UBs/nOiIrYt4lBOf0CVoM1pDS1gd
cdF9PHGDTd/k0Ppvx/DwhLxMG4h9N5zKJXl3t4oIAdsuJwiXnl+wIGbZVsRVcNCq
UacNLZdAkFD1GvHZDRaVVkrJ2MRpjduZBlbjP7YYtajnZgmQcQnbTK6YcSPp2BI3
DF/AX72jyOdUFJ2yEFZQlb1eQ/wdtrUMxQcl0ON+q4ReMq6frXI3jPKfNLz737Oh
sLLpfboJ8YpNy9udYG8Z9XjdV/eafniDHjtQvsRHtufonwS6hFENBvCaGnNCv5oZ
hCOmOwKCwEA9LizzZHGa+dhf8Hv0KoTlAGg4Mcix9nl++qBjcUw6T2MvG4Pf6Pg9
+0OovGSaV1qIjBM0SEkLb4GTlEY600SxDudRIydJAWFRHyQBdKX52V8QmOrfA8mW
8sgi2KpO5t+nsl+pDeuh/bIA8UAZ0QwNm+9Ic8oq8KR+rFMDCQjpArJQUiv5XPvc
4UiPg1B36guhotsIV45BOizVy49DUv1iwAjZDXrYsifZ1QKDM9uQvXuVWk4D0bq4
XT5rxZ8qcd9ebPJ3vVg7iUviAyLk/FvjVmX85Hqfe039JLlz5SdwDKBL8z4UWQEL
3X00nMA7uEMfmvioPhUu8+R9SCmAat6+3VTCk8tOYtoCYDqt21fahkv9lxROLRwY
i+MoMuKFsXfuewJroxYElKbawCsqNMr6RnfEmPdOaW8=
`protect END_PROTECTED
