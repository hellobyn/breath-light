`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1PefvrnGiIAm+C/oZRV3pR0c+M88RDCnT7Q3kMhND1uVgsFdScXSdj1xLPIPwUo
9yCd4YFQnP9Sa2C8CyaBBORFrDSXniR6Z3xboB11aRMxt2iekS4nfG88uq6wT4Eo
pzPI6s5l7eK0lIy1k1yZ+to/PRmpPrX0AP+dGp8sZnGxZU+eeIK8TmJ3VIc0xYph
KponJ05vmbmqGGmcASGwv9zD7xzi/Clw2BpngJ9oEK/i9app/DJaFunLLQ2wMhJ0
U8kqLA4xMFVLQ114QKaJLcyZ1NRvH6/yWoGmAhdXJ9zmpYoGu2wuC0yKKprmiFSn
Aj/7Fo2faCsMqgDGSUVeAQzO4S9FTrQisRsoLdY0dVx3u8DIaUAfNwE3qwxlFQRM
PEv0QwUUkY9LeREDUFYgQUpcVWz8qHGMlUPyV7kbqZcQVyZ22FVKdEfS04SCzY/a
x+3Z3sFCF/2hU/aEd6JeLW5CH+Biw6WbpDB5zvALg20R0cKUEjIoPTeUsgxt7D5W
pEYCexogWMv08juNfb14eK51Ai+O6q+AXQLDXnYLPb9knqtaKZWyM5xDNli1NEpe
+PYQ+du2MWZu5zR/ZgF0epSaz2QMuz3YTpOwvODSQ3cv0r0UospGaJEvo4CdeU4Z
YnaxSX0m+QN2u/eD/e1o42EbTLJV89zjuclw+eMweXrv1RkCt33BMXRo4yP+Amf4
2UlTwJ3/Qpi8nN5Fsfu6Jy+hx1bxUUKieSlH5rXqTXqI+LyXgkjXNZti2/uM/ki3
sZdDdCu/DOZG+vL7lGA9psgvRTi4CyGr4Q15gPRkIf7LbwCGnfB3T/S7paC0Qs+1
PxMbsroFfQh/C3S4QGlcnSYnEAhGeW1DXP2mJG7wcDKa30lWIXtNBtMeWtFop97x
AJEwdPnGN5S0PYt6wCssb/qmEYYls65QPHKILymxzOsn9qdWYuM+rmSXQS9oyrWY
7G3ZlrOELi1JEKDKUSVcHfEhuiEs7aVN8vvO1le+qbDOGBOUiF5QzJq2ZfBunGtN
znku/yQQlsK7r0QYqSAX1H6EQmOH582LDhpHZfEhAiGsngcbOW+0mX5K3itB7atb
TcuG1l1fMT6YTz9vFvm/6PlpsLuhnGPWFSx9twdzmDjUpvFMMaBSQ4owTD//pBqz
8ZlPGoh4QU5IM/vtfS+YNvLbz6VofSvhhml+2h+VGHLK8SvPsLQSDwKM41GIvnkU
tdi0wPgXtvaWav52t+buHiqzHy5vzEDKieckeigzaLotU20E/cCDRTK6MpbDMFJb
GTMDSkfUD4czBVdy/WRwBsVzFs9jc1dp03lzjMXiUcOvGfIAQNtUzVXHW5WuWJ8j
xcIv7M+WPKyuPp0jUn/z0OumjqmKkmWNTBzxW7c5DWhyy0vuhHqJbac/14jQ74PN
zpB9CuXPClYEZ2CG36ggrI11tlm5CFm7nle17utWUgfPmdqjbELxgv6sxdn36muT
vtc11wgNAUsDgnnQkG71mDD+6cIpTJPi4TwZUXnliuHXuxWSctwBIbH9iDCDgAL3
m90kyayP8sbllhnXlp+zIvzHT27lnp3HZOEirSjIU7POMrcMvcSmWQDiNyUAYlDk
d17Gpu1xYy9PXjW15ZfI4w==
`protect END_PROTECTED
