`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxNfJlcfbLZUnuxEGu8ObeynZjuT2vv1d3fZ9K1o50jOrbX4dD1ACGzV20Y1piY2
TpghZg/Jv6gFvlxVBbUxFsAOlDaeBOlRzxn0DUQbabsolcDh5G1m1HIVH5j/vMAf
HTfayhutDKXbKL7HuZ3SkG/Tveb43YLekAR1ulLYrKCWQ3vm6zEz11bF04O+ZIT8
vcabrUcFtHlJeI4cppHmf8Wbxp5KjKKSeNg9pJ4phcam8QJvePELATtO7EJspJdJ
zOK+/V3UQP9y5ac+apG0E7610hbu1oCw9scb0DbDF1XEYqxUTpFK0u1JbGsYlYjX
KfqD7X5g16IGblznysS6G/NVkXmyqDLsSBOH8SwPsuvuQrDV8W0QCt4OHb7VTlZx
zZS3Qb2ZBTSxiHEy0uhbkoy91trVdmbxdrC4FnyKviahlMrydgXHYO9tV7SLC5+y
MwsVV6uozASM8OmOWn/QImm/iQUHHuPInR392IMmOzuN52As9BUHj5BhLMq9zwu5
aTvEXIt+kcNAp0PfDyaIj47BCUzNQ7imsAMhwsN6kKhaaK5uXl/7pZmCnZKsQWFc
plKN+MIkMfX/Hs9Dzr8O60nydkQRLRayTQWkQ6JQecU2XGl7GFSmIYSCAcnCWtRL
6GSbS/lHwXr7KfFAPrqdS2IXziTPFCX7R+OB7lBVyLvx7TRSwPiu2PCbaUCcYeU/
BUMV/yer2FOc9Xv0VvUPmsJFocPV6wM8LRliM9LRu9oYu/quB05VRw+qCewVbzPF
MQcIZr3q9Zs4v0aPxq+YiBFgSl6HXr5bwDzv+1d7nZLMQtX6it3T02SjyYjPJIZT
NbDNzSQyxfSiWagCUp1+r9rDxkARR3K35bd2kbLnfoSUrPxptSPj1Lk8Fgsoc10D
sKh6jCpNfOwK3C8t61yzV7EtdhNDMLaPQNc1YoeEFB/8q6x6DEDQE3OzvhtKjFK4
SU6MH9RY/uAlfm9GR93biaInc1dBTqkveau2PPjI7rNdZr5WOgSvQEpSxeI1FR71
38Rld42puUGTAgS7W8PhX+KdPgxCvwahiwfHixYOUe7YyTPzYepK6Bc/gRRt3h+M
lUY/dbN9PaIR3Ggs4luy86TJOrf/dJkL9r7FPxbOJfzn2s4d3YjbkqfQa80dZ/rQ
qInfCd5S2sdH6cRodpcUeUXlWME0yMGcFPmtLoEe33U01nFI1cTMixjnsG+g3GLw
AQJNo8Ov7P7DwSc6RdtwaOfL7urEnuml0Y5IZUOu3QMcl04Vyv+TizbnxRcVrUDN
IRX+Xfr4XsWyObLnoSfbgttG1cNqRhbbVtmgBePyqkCpV1qouFkAV12Vl5+XRSWW
ksYy7uKd4xZtkS/Ci2yNjiX0JUD1fTLkSCCA9lRChodpdgl2aqQTRQVzVyv+FXub
ViwChzx/Vbqf45+gH7D7qCPOdXDyxguwDC6tAFo5HPrWsYb0cutZfoUCsypNgRSF
XVkkIQODTZflaMW0N3nmpDLUd232hx/nVDgzvhEXserZaqpNyww250Q9mZQ4dFFv
FxOvVnY24DGWDnEogjNG79vLMWLjSPTMx58xJf48xZs7AaH74p0fEBsUlmmg71CJ
FdtUZMEAG26XMjC9E+9VZYL44IlmI4pL4OiDZYZr3BAmis+bw2Kcn+SyHP96ur5G
4jckeWAMTJImeoHfBr4k9nO1GxM+ItaXSFvT408FaYV8bZKaBFPphzWXZn6ISnJ0
+c4K3sKdGQGtv7slIoYnO7nD0QPqKEIjj4pTVkP6/wxh/yl7ACAmdBiYOYfofZ9j
RDYrnkDMA0lWtrYyjAuO32KvdRV0/Sx3qe/vO+5eRi1mN0guOXXxv6gJrpuXo46C
Qz9RkLRIzKrAbVAZfZzFXyEDiHnIW26bqd1yNUXoQFEQm5Suzugx59oCVSncfH2C
+MoZ1nWUCi4x3dxp2gu9nCX08/vRl3Z6TmA4pcY2faSul8y+qCXfrSgjGy8ojVo7
8alOv4BlU4G+s4DzOdNlnZ6AUbfY8uJr/EIEYKa68S4uVZxyFd25665aSPWBbrhe
zoRv/Q7UeT2eUIWo6GCJFwcyrI5MzwSX7bBYjeNzWHHajAMC3oD+tPa9TnyHP8Ii
f9LUFdbZJh9++FVtq4bOcVPUyWl08zivWZSpuEsBTWeufhLa1EVxVLHos2sMvWEg
komDdQigBzmu3KAyDXzGa6p+pLKbRecneMwj9jMM8UYU1BLIHfg9QB8I0awiUCCe
BpyItUMbg+C6UWtxCljV1XGvD2C+u7HH9v1WncbocrNXUSoMn2lZlOLeM3KEOgVN
QjLGbpdrCTfj9KqzCg8eK2pbMtcWKgmNm0A9+Ww6FajgfV78LmTljuWbU2QKx8+g
ccKGCvJyOCT4Rbu/h1yNfB/g+Zg2BjMNBjparBT4LcWz62gZ6ryI4Ptkb28O4ToM
KN+38E4ZmUDqdv4NXF/jV4GpifLbw/Vy69Dn8wjtVkoOcduD9UUlH2d/T2LDmsTi
uXAFMlKgPFoS8FRXM1pCs+GxqJ+d2URIT8auQh/YioXpTJs+uWR/YQowY9exMiiK
02PweloqcX0cIXB0pBbzZLIOHS4FRUDdlZrdcA3Oit7tO5b8vHsrVUZnlC33T0SB
upK8oI/bSTpR1UZHIumw5+wk2wQaggud1Tv/ohCWAMNntGNRu+PjYeWExITevO3K
HeGxWw062aipDrNpuT2WUoCG34BXGJ8udteHqoiVxnFJ01XslrDMrwYG7+Yy8job
iunSHHYGSD64KFB42/6ERVHUbkPGk72z2yoZLzQmeuRBGEywrR4Fj3i7Y9ltk6rx
k9febpKxM0saJhlp3ZnUSv8ZA7BOsxbl9NivFnVfLEhJchwEG/6ihjgIlqW55Rbi
OFSM9ebmogTKI4PVC2ogVK5wNUygP2NDl3nLz0qCGq+XTAHYRzqecfS2oxhyv4Fd
s3gkMv1SuI76cjgpdFtgAzxGumIJ3iScidABnCHFKObkgDPR/jGgwZ4J8p9Udw6h
FlMKnEPghu2AFsKNxj18z9lCFo5IMzAmms5NJMKSVUl2YdMMIMZcj2UZVc9/U5FY
j6nNdpMIierJBB+f/T+IY7yQASzKnBLPDUNS6G5WvYmSnXDHlMRp2m/uTfWkL5ac
/PFSFm4AeZlCijg0MjgZvVmNQ3opLpr0rZsw0cVo2nCw3Wl3ac33wkhF2MyzGktW
pOZpq24m2sm7VkWoIelEbZ30gpwlse6OikmKG+Mq114kb2Q4Do3dimu4XdhUtSUP
30wihAv4Uu3EDlY7TxhySCfNNWkUZqxXkGhTXn0vMfx/QY5K/XEB5ntvQKfgq2a/
zXdNyqVyJUfVuOX9c3ChpA8n8JTwgqgbWhWlE/fulQZqEQtLT6cXRLjW/gnp+HVo
sbDWPfleom65if6ZC3WcL5VLsH2lwOvbq7HQE0buUaH0/5/xMKkKmWnfZEob+Yn9
TNYHofzNoE7JqXg5RPnPCwCZo3rc2WAvGP3QKW33uFS4EBGKpuqSyHiXYqS2Rtet
`protect END_PROTECTED
