`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uw3amt1P6M41J7FiKg061aPT6a57wo1s5v7syNy1yMlllIytBrZxC8sG2L1TZxGz
yCYKFhxxGQKmMNAf0uB1IuFMKWWcKfCbEPKyxKpySfOBLqgXbsFAANb+6Tgn43Uf
alk0a1a3APIs2aT3FPkgfPAzY/thAalvj1bfotUfE/xQp8FSI5/cdZBRSz/Lbv5s
0BB7SLPB3s7qlrHMxVNs6VoUSBvUkjV2EUxj8w2qMwqdgralncxKBTqK09RDC6/Q
OZY69zbOUmoFJVom0Eo5F1GZf4qvq+HozdQBklrlAywh1g9HdWG/L/M0J0MbVM+7
AyuzoMHe5vfkFcj6qldvnDGBa8/DmLo67n6SqCJwPpTTAGuyozcLtnZH4Deyp0NC
Ozv8XKVdjaZGeic/hwkK41Nus6xIdIhUpmwFqeYyWrhHd7xoEsZEzbL5lk9OPC61
iAXTSiujUb2JxBU4YItCYstiWXlbT8WMRzIkzmV8kkuQOJpIkvYFMCreRRjsLC80
m8tAuDOW00NOU+2GC1fii1IK2WS2JgjIlO0FCEs4v3Z03IeGypS4IeDkOV/6FLCi
yOeNerjSCu3vyahf/v0i2rFeIw5aIpJDeGpY8YilKzzvUP7wJdHnnkkTretmepEt
j7LSP97UQ2P6fAIYAYjaoA==
`protect END_PROTECTED
