`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pk9zjQMrnjcWbm+lVsV36J+JSs6//mA4sgqBeQwGicS/gfJCywrGfGYEhK/8b6UZ
XNWWZ2YLED4SpwRXLeEyy2t31/PK+tEcbAXf5NxcYUg6rv/C0wMHABKlXJmxKwkH
yxbXvM40cGjvQprW1nPr2dxd9FDED0EABugomzjbSEzhqtUylKxvYxmWhgd4aEq9
JFRvJetd4eOAl0M4E3B12bk7WOSapQKtpo1hYL9PM/H3sH2jcGkOBZ9oXTKWrlBp
bSDvfHkChK4TJkHycaBZxP4kI69i660QR9kNqWVol4zMiTIXblN8YMxqzXfUZhYR
i6HAtgDhaBKC3gtgnoaBTCdKYIUQBIP3abBL1uOqzVdqnVVkSqNCEokZsT1jeqIJ
h4vGIMDgx51VLW8hMMS5yqBVUs23P1I7wLeLXaNuVP9fSz8i2S484Zk52t4PUZey
4cdavo4l96+qmm3K5LwWp79zYsKZoUy76hRb1J35HZZISRp7qh7OiBbhJXBQKzy9
sKtjDQ1/EOHB6XxfeEYLu6SbIbHRA62EY+AddH11hLI8raZdquSEAOK2Dv968UFP
Ww04WsBRL/xpKJpQMvFaNd7C9QVTM4emp5vubY9rMh4NoucPj0GJNW/t5xAcFy9T
xRzUrD2F5ZgOJYAmMybWpEN8l2knmBViaMCXZNRSN4fijQn7ebjFwRj6vVI4T6oc
UVLczRCuTvgNnoNDFckGpAVUv1UOHINNhTKYlvY0KpjEQ7PVvxnneuukdy3WWRSm
teUWKEx8n5LwVkKYOdAjWUw2ahjTImsfTuorATqBxVcC+Xcp7HC2CwaIaqUyp56S
c/61wod2YwBrYJlXSrZFHtpADj88cgaW1GnajVaADxaZId3Q5jlmA3uS3245oRnm
Xzy3xh5oPwKeZn2SPXlhxrhnJWQEgLZNAEyIfnbCowpW6ZqerxLcVimeVDpdJjb0
m1Rqvk9ZWBuDlujfLz5eDh46feLtlKj0kqUR7bnTBJcYv/JLQth9FKFrD6MCXMs/
xOgr1AjQ+AP0LdAw1vXHMTAJBj0bVWEKquYCnsbPzjjji+Rj5p49JvyVuKEBfn+4
TRSDRXzj8pQoG7bvL2EIqCcW780oV+37w+/6CM16u/N8x+iaX6ErCQ6Drdu50QNU
BhbKuwW0mqpmaB9uotNZFM58sOe1J6OC8sDZliPXHUJ1q/WOu4/W+UGzjE5eOgyt
uNUHgZv7QXc9nw3sEToyqRO/j4NgchKzrBqHA1tgDYHFmDlKzvBvXL/nn8xPSb1s
CDMn7ZZF7BU6Il7be0F4KVuMsu3fV5RYBSM7NtLvMIWpkoGNUiZ90Eg1HCI40M4A
/eyfT9U2S4VWQpHcIkF/utOakqHfVBiEBi5bIkTxcGxDoUH9jrHjfilQFZN7dKhC
HI3gmv++pZxmr2U+lLOsRi4MIbCejWxaAN6cwP5DyP94zcxAFUqO/oF12SVAEBIL
/89KfCLP5bQxYlD/6hMxXVEv0GkczT25M+SAw+bHJ7oOe7Cn84ItmUtCuLEnQ2E9
77HrHRjuWVm4b47jejngcjq6PaGxDpEkySmlItIZkk/ekxXmDeyIvyzbJ3h3XfY6
Scd6ettNzdKbnvWm488sVHLUSlgLBdGN9INnxqILRiO0ppri61xNpPdkKVAQBIZF
IQAP+D2lDGSsqV20zo7yVDAI8Rq5mn9s/jWb7/Nvq9c7ACvyOnDB26MF+pjWIUuB
XE2Zy3RBnXjAekyL/4Cf98D+ag8J02qQKSwyM/J6xwjk9CS+csKw1Q1eH0llpqyK
uq4G4sGRzGYXbCfGT8j3IJtlXuQDfGqscmRbYw2IPlcv/e0WmtxRrVD+kpV/t5Qy
6A+XKVdpLLC1or7S4hLnEEPTmJgHs7aRXMYpicNFvVFH6nqwJyT74A6Qm4G/Q1I3
ViRckJOqCcy3fpAWpVlhrvBt244mCVmaXrLDFVS2elcr2KhGt8G0WIYfqWwHj4dt
pIou3YZlqV+em8m+lBFA2EAAr2WhjakEEwKRcb4ho+kEhFd93N2OYwemCQ2vg1D1
WHBYECTTx05wcOa5x76mlNWHY50fjIEFbrFJoQpaTjw3GV7j+CE3P2nC1xshRShC
oTvMpBfAE/x1U78w433z1IzyM1BRTvE53A7UpXjfG3KSziAM9LMQTHUWq29zKq8l
xZkMawYZVl6guLQovRUBJyNj5YHISDfRJp6Tyh5qWBLgKbW3mcURrOL+J/yZ9glS
hoyCH9iGnl5zedUwzhK3aehohQ2ekDt+nlXLJXHZAYw2eKwnQgUcaPsFWRJZH3X7
QLZWsmaII4LSfK65FBO7EiHlLkzimd+FUlbKkK1LjHm2xHGmVsSd5z/FyebFfRaX
DH0WWZ1YyjYk+t2l17jjY9xlMM/kxsFrtQduPTikrejXmWT2ewRN8nbQoXJb2ubP
fLIfNssLwyx3+prOISpsCgKtXtnv+lUGyX6+wVMzEQDD7LT1/hABH62ifVak+Ddr
rPWnfyIgn0uFe/j7X8OXTH3OfTD5p9UseqRBc2OYsq6NALzFNePQSx78ogwtDS9m
Au2bG+7e+3wZhMFYn8rNiwWRG+KV/SPZQ9IwUPM/hHNgkBehH3cboA/552S/DT+G
/HxRtCwy+1wh8tq0gi0M375jXad+aWK/NCkSqs4xLk0mfu8GEqTPThYaX8J/gNEV
sGGvNpNXgUeYE9QzSEyNBDk2VSL6LqbuqX3UfiYUrMkdUI8EYn6D1esEuZKL5Jwn
xFm1K1pm0AvFDP8b+2XHzhLtU5wyJTxUfa3wU16HzwJ3jbP/BqXSWT1TDCAD8GrH
t6UiEjVSTLzcK0gT3QVLtQ8Crv690GrZOVzm3LKCSyYQDtlHu73e7wBJ/7RFCqEh
36gcxSCPg935vqDo75WTtRSOzWfcEYigmjAVHSnj7Yzl4ufuzCGEd/lMmMKdzJPG
yE76CT/VDB4qs4Y/6ICAG0xJ21iT9v0Nke9mdXbeQ3m05ZgsKyFPay6/dJeaAXiu
ilpZiajqjiZr9v3j6298QT2yXvbwLx6IHwy/gToKkYHsGW82gy/0Vk3MORj6I2im
WRTEd8TjMUZWRafegFc2AfPHVPAFj9e+D+p51QMhzDs2774vc0dRUrKihU7u/W1w
fEvJfkqL1MrmQwRACcPf+xO4hqs5Es6dqJxavxK+QHuHWOMR8QhOcROHnqN2EsFu
aC0iLummujLHOt6zBwy9f8BnPIzGaxnU4sC3eKKv7Ukh4rUk111YcUDV6DV5UHSB
x5tbhSmHH5FVXqDWCD4BdpVzQOBGIFG24Nn56Qe3cHdJo1kkPWSzHvktAy33DYh+
/qvDloNKffdp8KpalqCQTNupbm/mHm1kSC3hquHd/clmqo0twLB+oAExz0RvFGZj
gxOpXI6qng/Z3PLnrl3Jpyoy1RmaoL6R6TqTWDe9BL/cdJFAzong28mLUCTy/I7t
fgU/6AhZ8/sVamARAimYOeF1tdHFEG5N0ss0gnNR58uKFi5YZZ7xkAYceXpsRvvZ
DcLr73D54f8gpx0uXDBDpLtonqs3WVhKb9mm/e3+hcJ4eyBtIc7U2DsbIjYxUXxj
lflgBeGSBYE2q0715ecMrTJ37VVuGrYCkXeKI9NJRl5OgcZOrQ8OG5iJ3IHJvjnt
V5Oxt3IlU1JIvQ5raQ1QDvLvrqdFZ4WTOhtHMgqJqxV/CfJx3Ucewjj+FDpseofk
8ksmg6DiIZJhCFyl/oVFYmxD6+e51sfqqXPJB94QXwQZvaRdLkn/LapyYgAoCAh2
fD68GDsMVsn+UZtdUHIFwZCwEpTwvLfsYvQY61g5MFvzhcAqfaUDk6wYinhIKZ8z
xDQdTZzqI/1HuD2XOOgd65mUeFmIH3OJneuTXw09LP+x4EVgM1PW8sRdn5xnUppn
lrjnXDpZfOm+BmL5zGQIhSPN1iONrISZIPPSzFfNLXUpAQhtuCTDVCh/zHTTstl0
xj7qTtb0wgOszaUnOJH+RoJblFTBhbX6ZwHO1ApYL915v/kf+kldp6NDm7Nph9sc
Ybf0HH5kk+UUv6vjHbA220i1kpKNXREUvQFeTZlM3iOU2RBul0OCCisMwLXrZSIG
qLxDrgHjSvTvXlbWJD2sagB7E1faCZyCBswh7SLkwYIPJj0frwyL9westEUIUXhr
UOEc/+TM2tEyynA8DrPKMR3ZPqiJcIgfvS2pOcgsJm8mZ461kqdLz4c4Kcspyuio
aWScf8aJ3JU47/rLJr42cc996JNtoP9WPen6zOiOM3CLxPfEur+RtZ96wnmTuq9y
sNOIzyoteCsmzZnb8AfZACMkcg7WVC2TZzL2MBQLXpa/+24l33/Zps2DntUArJq2
eDNLJGpWJLcOklmBaUQ2SP0IZEzMzQfkucHMnaFxcUpUnx8BfX9n4Pq2yuLnj/ly
89OxyVV4YdBkvCSLUbOsVtdPLvXX+DEkRTNgUUJyDdFbpX1Lr6u5XtyWDMg4AcEy
iys1x02BszXYhXo+Nwvvpy9IMg8LEtYzyHBo8XcP8IwN1toeX/+WQzZIGY0F0ru+
jDgtRHxxLIPNt2E0LliqB1sjqT2vl772pV48HXFu51c92JJymJQoil5OMotbuvbL
LdYDNIFTCqOJg79Zpl3HqJvMlOkQAVa8gbCo+4sow6om8NhpJ5UbvmCPEJBUpAmV
SEHBQKiPPLLdoaKlBffuUwvLpNVTZjGwndVcM2p29nxUDCZQQh/v97CZ3itg9FEt
Hr45JaQOgHCeehcXWILUASzukA+Ui30EgTHLpyPhhoaYklbz2Uf+rEy8ogvGz24j
4tAKj3m1wUP5V0CfrfppFPFUqkwTdEpORpOxfm8OwZN68dnsF6DvCVTQm6mFIhEh
RIL1P/0Uam2DtndnhTvxVLzIFnKzRIN6Yb8DLPeTsDT4op495pTNJ/f1JxWCUVF6
DZxkmuaxxxrB1TYWV73WLA2VikaAS/PVhuMXjJ0Suxd0EW+jmCfNmZJxfQ9K9FlX
w87O1C/IoKeTOPahzrQ5BOXiiCLfkSM9t3o3wK3HaTzlDQ/hcLb8biwvgSLmaQ8U
pd6NIf0/XRptBgbswpJuDHBTnuFLwmz55+E0m07DmLYxAau8J1cZ1BEPQpWd8OIF
65uDhN9sUHlDMujWc0cTSFsor2gzf1UbN8s+PpilKE820eHsT+amAkCwTVZOX+AW
LZ6CI4RngbDZYxmUhBLjD1W8boDyeQWj7BCSwdqmfMJ3bRmMb05dJ1dsuBrPWx81
O7UmOIpqverv1WZ9EU5HAzVbJzhlTSXaFNi0hZDgDPIciP0CLD+nglYTlZrY5iG8
mA4SU4AN3xUQVODRgkkRAr4c/gmPFdNe/jUTGG6f9A16S8a9bUsUF8znUP1EA20d
Vil954TrnFI3JtsTdwRg8lCpra4pC53RKSZscZDUVLN/yPBGP6jTbD3q1H5qs+gg
mr3zeV+S9gfHsaW6PwkPDcderaRU2zU4SPfnDFdjutX13iTt4M0scDwvhzS8Qo64
PFkhc7c166T4or7o6jkClWQJrbJmivBPwX++iA+yTxPLQ9VGiuKIZSo2rLKMN/Bg
4V4bn2rWKNAOg5f9kPcQiGVjDk6DRleVkqvbRhVvLnABu0BcAVOEqurbjdFJkxUb
q0s6vffuKewe46Mg1LH68A43k+rfHg/7SDbHU6v+gy5oAOO/Um7HvhVWC3Fzop4+
RucUG60dV3JEpg5EeRyDPx52r55Tt4Xfydt/jdEtMIdK6vW436h4uKy9AWy9rLTq
6Af1eOi3BBIQPOjZCX6tRVKjuAX3ipmOmm5w8+taIISEiMLeSdoIbSfe+GTN9fZF
22XKKzP/a50xj5ELeR3z2blJDyBMtwDqigutvRJGqNZgafqUzqTMajMZPinrGZ0u
JhtApz8hyeE8gaAsBZESYEooCVgJqq475QhINB8kkstoiVI1M19AJSVbDVuh3LPu
5HJoCl5jNs4mU8eOyzxT7AvLpRxrBoNGHonunIW8Kw/VPZcGc08VjFsyRSaqgK2O
GprkGZvBtJLwuPQXJTMvm4OLlvd9/owmru/JV6//FP8qqvITYK2pH1NjFYfuNeyo
`protect END_PROTECTED
