`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LLEsIJRmSE0nJzGcaZb8Gxg4RtAc+u1IESJoTRdRH0q5cOBJm0pZjHQn1axb29rq
z0TxJHTQ0lPC2YzaMjCknHIo3EUVnr/4QahdBnhhBJkpfMH2D61vdP1DBApKi0e0
RhaSI4ShfnM9ZdMhjKpu74PSPEpdn34RvSJH8DMNJhSYW8IQ4Ya8BJUApDx9IBHa
CItCwqQ2tKRfA5P6dB8V4gfRMr+NNAmoXUtDUFVC85a7Csl5EiV/dykBuPyL6j1R
96Dmeq1EyZpsuY7fVYd6T7i/FM5ih2In/uk97EotHjEkF8uTMwrlMNNmaBtBhT3Y
5rH6pRZMtQv/MMiD6kUzq4VwG51C0uFcIbBZyvjyc33FKNDI8yVX6ImYOKxy1Glc
7or5BImd1qQQ1GByTWWQwBvqGPrx2thRhB9UoHxwB23UfgV4lwwQB2RjbzH/Pybw
TxFwJ/V0H1YnGx2nfFKedOqJ4tmnay7SqT4L8Tcx5hMy7bX6OkCk1aiCSDgi177y
`protect END_PROTECTED
