`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bnG3q0BXzJKfG140Jop+QwWTRgIhd4/rsK8wTPUNScRZ+s2r1Ss4qSPCoOMGF5I
DbD4/d83NGa17WQbVwfTqCq5dRFUhAghVX7ABdXXvl89xcpVCyg5qg9Oz58yXYeB
2jppRdnqz6Y6vfIeVsnoVmNjaxFyhkmUGU4sUh81eKLly0GY1s/44abw1wwYxmP0
JQJ4pSc0bOsapZEHseuWaumn1vLT/ciba48XJ2RXGwYCSw3SDXXqCm4/EHuBJ5V0
b5BHbpWdCWGdVVAGsyNzGo6yNxW6UQr2yJua++XOsSshuZfgaCaQkDuoF6dYRnNz
wrTldxXvbE/GIN1/4BLEMAmQZBsMJTqodwR4iLL78+962cPCetYsEv72Zm6NGizc
abBSACsDWXXB87aNPjLTHRamdPQCI0rH8paYxgWJCXkuKKVqOG6AxT6hZ+yF1JJ8
3XHgthC9z/NUUjUB5/AxBDPDtoHYslR6vZdDLxD6mGByu2vNKLHFJSxmD12uHIro
qszyN+mkYrweMxfrLOOEYIINc/A31yLYXA9AYHlS0SQfP5vLr6QMu9kdb/upQVnF
4OSq+PhDmgLi7m9kDJNdhsGV0+g6eVgyF1ZIY0JrUYxcpSzKxDpQRvKzhb+MYxLx
TTPyumrehTlVxg2LNT2nIfq+4s1qnVc/T49SYiDWfNkC2yfd4yvZCks6M478gEaz
KL29sgzpwzHebTWveWEGr733p0C4MhqWcin+d71lt70C8PM2MB0MowqxXliYgvQf
Bq27dcvZVngUWt1i6i9aAAHkTpo8d4UZDzZEfK2D95Xc4slfv9W6hrwGSgnZH1vq
P7Gb7SKeT6CZeeLZCA7t2sECg6nP1SuqVgMtf6kRTUuVM2jLKu5G4H+pvDq0s14+
MrhrEU1WKB1+WkFVPAXH0BKWTPIv+/1dY+x5KO3kaSpAnknARO/HvOCWjGZnxLiO
dMnGYEI6B11SrYHmLpmlwXA7JRjxlPjz6blJXa9JxgduQHAS8XFi1wIr2NB+RfFD
N2TR/xpljiEJas8oOVB2YXf7C/9wzhxMa8c9d4ldzaYwwcPf9vSiZk5yZHpbYqXI
1ZQSGtDWOJq6WQoU06Kn7zX5zZzLTzgs73qNF/Hd7+5yLdBqb1oN3bO0CWafDXup
8ZJCdFu4pnhhflJKOl5HCGDSaow7vU1dBiYhVukDbz0vkyMAKDKdegjC/LaOn1lR
VXyh2P4Z6csn6b9O2SG14x9Ac0uwQtsjaps8wpzjm2+3L0t8thP3V2gIzwO3MPj4
420uSLsRok/lrNg+hDvoe6FiKbwk33CPEU/wP3Cj8bC5Fm2/zuPktINaMbVT47aA
L9svgWAwKQzz0XAKzN4ed5T1gXr0JL+sn3++ruBZxHMCE3swYAlcIOXNJwNBZn45
YkVGCEEbbnGuhpx5d2TLmiakoTX+19HZK3sRX8K9w359n1bpFEl9FYww831uYS9W
sLsEnJIseMxpbWUKLJtla0BH7jsfwpw9j93wuwWLk3V5E3BndPOkdrSiVze26nnM
Wv1Flov193JTun/Q/c6BrfntVtohDrS97wksQAeK8fLFLDT3Zhog5AsJkC1l1gb7
/zoEKk4BEzv7VxqapmfUYr8EvBwXWoH9kZCbN5iG39RyMiQ1/UWscAfjTvJwEHyC
YcpHFQiCNcrZ10KLd+JJqNccaE/uEbLBFbBGtJoXcDwKUmJDx6IBX7gUwEVEPgqw
GjAsZMgZC7h22ajZ86DJuXJSd88ss4t/YCtlZ7GP1j0XhZNUB/GV9kqQrhjQrSKG
i0H83/uHP8hTfnh8ucxENO5uOUcZlInSNuulXDUazx72TeE5jrSblG7jq5ctzdei
ENykQnrPEnqG9ohj2SX824RyseM07K8c3Lrg8yFV6YKGOrIpSNoGslgHGBQtW7dG
Qvwdfl49ZSXyxDm5tprCjw==
`protect END_PROTECTED
