`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJ+zQQR2jKaxCzYBed6/vHn4yBUjj6f9t7iDRfLQnSrjqXGxBJsK7FObcVxpZQ1y
0GpWhrY18ZgGs7pfUcKUSEYQEPlkvBtu9TLiPFLgnmFfKmdsDg7fRq0AvVCq/LrJ
wfhXaLhtIMIm20WOjLmuDcqkvCwMHnstL0da32+Jf/gubFFNOhZo8Gj/0SXOSh+X
lhCyIjHWkW5hh5ekBpezBYb1GnhNmAfFZCAeoSZ5dLzIgt4inSFtzgRTbn84cX/E
jdc+RQ146z2cL/+qlEuqwGRzGbOwQd1t/SogfrulRYtv6fmdXT4P8z90iaAs3+w9
4nYc7tpCQSHtFjL4WT4h7Ndx4Fl/ZHqrUVN500lSD28BHT3WgDJ8RvT7CoeEikjq
yDDI5+Z4tTU5/EYBbc7FpJ2khXJ+RCoJhbWMOLC+EtpczmDguB5Et58rbxjutlq3
44XXVXt4sf9Qy/R5trKySu5YkRRAe6QFx252zuOKV0PH+0NabTbfO19i0lCnYI/V
p6yrs+z9JF3ZdOqoT+/fOQbWyKkoTJhctePtzr/YZzAZguaprItjTbmQ82FLWaPg
C2vppna8UroSZD3iKIY0NZUBHcY7l1K8qw0m5QdFWbyOGM+1RUfLTJMG2CvAvoaW
nj1jLPVrozuU7wTpZPCUblYcr8/e95L1PTN10s2PPfI2dJGrBT94sAv4FPu4U2xy
GwdJRQVdIx4PjYUguyl5kl6MqJuMtbsYGywrqU+QQzgIIEOYr61xn9cGKeSaLyIG
J9/r+Ho+GYDTSFAKVsgMWUUFKMWUpUqmjNPXBBu3wlfKAoQz9yPyqpmJvQqVtlcQ
jPg+YJW/80tiPWIsVVt3ngJiPnTSgyAXQkiSK/LxUnjWfdWbchCXP6co1yILUWR9
49/v3Fl01xSGN87eLRfWf3sYr72NkabYqtLNgS/F+2d3osLvcCizhe9zZ3pEIR6E
RaCLWult7I0u22z6Ssq/ENb8VI846D3XLaFOm7nMy+DHOhuQ23bHh/B10ONUa/68
Woahvz/5LiuOPW8oh/k0g9ZjUnWoNGIpuMe5qlmPmbYWFQCsh97QKLiUJRmIH+bl
j1krdcgbsgOufXAC7DCt/hRcs+jqqoOJbhgxAE8u1CY86ZZ9eLU/fZKDU2qxTwk7
x3lJNeqRVAiUjrn2lX9uYJc5XcdO4FP9hcS5p1Go438giSaDkEuKIoHEJpR9EI8D
9oLPkujnrum9xC9YEn0R/4hXsMmxGfDsXYzmXju9UAmG0/mKOyqrm/HlbOg/qKi4
XYRfE6lToeTW1L9ow+38IVs5HVpzpddfm7pIj4/cZtL+cwH1VoMEdHKpMGrpIYHH
64aBMTFKxwkHg5vrnQQMEyF4fOBXxWv6gxCjb1Fmr1lBwheKo1n/5fZXW+zSGjGc
RmLUZgrTyIL7cbFpxCNtQ5ALwejaMtpYhHcBZGl6HaUDX1pLcfHJ9gzDm+wed1zr
6DvyJY+bVMP7PhPDc+R5isLRRNECE+uO6eMt3TNf4jRO2LWpGhxhFlGvJ0BAty5y
`protect END_PROTECTED
