`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLiy56fWv7PlwtEfw9V+vKU3mkaLTdrV+3QCHZBBB6qiwvVaPBPL5I/hWt9FsZRn
U2cVof/8mnAVVlXOgVUF2kHfjODs5qQeTlBc66LrK3O/8li9PpuBU9o0qtL2IG64
/X4q1qNZylOTeBZw8Ew2nap1N1Fkyz+2c8tRsS6xpnWZpZdcsb9k8bydS0fKlsBl
pkeNNW89XWgtLtaweCyQ7pCBPjbulq1+UcszmZAdNlA5P3i2faVGnqLnpWvOJQ1Q
qKs0WIhrmOmHF0CO8HuZn2/hLc/ckwTimc4RU7ZsnNs3TdPJTzo42xk3qNAViOka
NFux8ihO9QqhnIHQYdjL1jPBZqk8p+jGBl/uKQWZ6evskpa9fuBbT+hiYNaqKsCJ
rxDBVhZDtzRa/PLXoI7i3CrHW4OMPHJb84UGghwMKXY2nZuPtgXmWGEhTA8oFwtL
6ucbJZlFP77wiR2Wu98bTfcOeTON4BC0uEoo4DxmHzoavaZU5nVJedax4jl8eBSm
ybQ53FhwDwpfcYoyWV1nI/jP6TDfgHVYkMUOMxim9H08q8805dJXoh8YlRszKZqn
qah0QXGaqEzz3gLkEHPQpjqVzZ8BeiquBrIS4Bz4igwC39X14IBq8hyCLepfD9Z2
9gDynGQ2rkqzvVYCVYMyNL+hu/uONEZRva5vw9/LX0t31Cx2rSkvekvO3HBxJ12o
GAdBx84sAtHNLPAJ+oPBc4Iqy+ulaCgCEiY4fnQnJl5TyVDPZ11Zc5MLL71Uz+3y
fFDgY9VnZOy+a4iRHPxf4PkJ+eXJhmVjJR5lo0nXRfLKHSIQy48I+CzDi+Yt2KyJ
s3G1hKx6r55lqY2TnYCEq5vZyEreuyQKuJSqXiqbTv5Xy8vXwc9Xy+V6s7q24ahX
lIumLO/DGbnP8Ffy/Da/TrYhJG17vvaZqDp+xYh+8qjVesq92rLxoeGtF4vWJsQ7
e1RnWclgN960y8nSgpGN3eLJsIHkDQQdU2gxDndHS42bcL5qXU3wHgL2FGuUgtde
hsbfLF/IWRnF1n+1ZNMPylFneEx2oSPFtCdP9AlrGsMtPQE0Cfrs4ITgTIo6dZbf
y4LXRSydJmu7ChPaT9zGHNjnmSR+PpLMkKvGO748hQh3P5umVLs5fT00QON3hUn2
q56zpzOVjgYCMc0Wx8rfaS4RQfIG04t3P2CAbrgU+9nl3XivyQnn4lDAxby32Zyl
waOnh60R4A13TcN6k3REFhaQZdOkTKq6WnAKLnLmFr9VUWBN5dBVivTqsRniJLBX
NZlRcUg4YkAqal7S5f7l2WSj7xg3l33WJmfiVXkG9+sqpno50z2/9EFC3PjUDd/R
ZEOcUh/KPD6nT79dbG/jV8zBkcvbKjwodL+L9HdFmHF4ct32kimF+P1cZFOfnK2/
Ks5fPMVnw+doDwpSYPvzjpeA0bEBjSPKPJsWmcyTW6BlIrN3wwUidds5k5o0pD2+
NsaKj+ynPBtBYz68Inr4r5Xw/UOOORUe6ULrNajlaISyBV5cutaCEwfpQYHhmT//
XB0UkMcSuJKnrl8cQpHAuANq7VNS8akjUGlgkKDDKVg28PIvtvjQiqvtohtC/V7U
HRx+v0/T99/PBI8PpDUc7bAMKe4+v0vI6B3/5SZti+/TBsweplZl+Y4TIgL/2Y/k
IEK6O1algIrcqJmVm2fH1ML/4Kq/VkSeATrYYmH7DoOn9X7eHAMBSySoGFCxrC8c
vtfimpEY8ozRCvggkZYdLJUtTGICVSLura0hUOqSCaCWtZgKl59fmcZ/ioKZg5TW
F4EuTyjwdlh1Pw4MrfuDNK8AquxtndiXI/kmbgjM9G7WqzsIICZwseP4MBYrpolN
uabAnforE6sNiddNbdtnomCB+GfIE6WtgXiS+Gu/UkQ8SibatwJdQNKvo1zmMeCs
FVqgig2pQoQlcyzA52rKFoaidT2JkB9DPgz+IYZwyIT4P4kLVz1cFZqG/Qwr0rvN
fYTkLOnqiWBlMAr2T1h5l+DR9kEeaArs0KGVSiOSXo42wOGjx5KZbFpbbImTMQPZ
hq39FykCJNcBhYmHGWjSR5fqnHEDk8yZw1F9qk9vqr0ZEwbwuOcAlp7G6ShlBvss
pSnZMRLBNdoiDNrQ7XmiMyoRah0X2Sh+NWKVrcLMTGf8BXPLJN3INuJze+noH+02
kDnyp5TfLATv+sGi/iW4rhJuXf76uvamhXsEB/nZ8Xz15MDfcXioAZa60mF9lo4c
jypep+BZqLXdp70MuAkxthWbJyUSw5Y6VRX7CEXg4/a6RWS4m/pueEFA2KvDNwzh
+snUhtLXVJoUpRUzpqJKpsgUFwlCy7BwBbSa+ul4J3sNwvMw9WIfEkTVMeaUDk1q
gGSbRk4Rs8D05TB1B16+CvIt8DSKOoCfdkUxPYMIFRlJVds/Jp2XkspF7PE6GPTM
iq1c8zk1EzCWCo/cwvG2V41nV71r6Saghhkn5Kqln8MkbTwIP/TlmonJ7oO06hhp
Lg7+5I9APR0IMIK6qWL1b0EbR/uGhrRmSRdvkHnfTE0DXrzdCsFLWs0VoS7QasqP
imcNQuYYnmgatuNsXuhEletRogn7+yeutQmwEuWNh/AIRcz5RAqGeMNID8hWjtTJ
Z9erhB2vCVHDbVjNBYUl99+FNHr2KuEls3zzgAQTiX4AdIXyvdotyf9lw/mHkrPX
b3OHXyhAZ+vchHhdC/kQ0osA4uAU7UlFWGvd9HnKcue3BMKOE8E+cTtQg/OhxxDy
D8122OoGvx7412kuALZq05M/xWhR1GLJt8BgqRLAv9dXYds/403ed1MtuLoXUcEC
JSNVEGTN8BO+5/3wDoTIx9wyKcS4nlUKmh9TsF5YbKOgJbJ9pR/f5ZzDzV2kC5Zs
KjZqLU+UpJi25Fio3DX0br9xiPUxAPDZ7NHXGWDbae/EO+UNVl5GWFpxPGNUmofC
7aNaRWDUr0fHfI3jJL2lV9U0ujiF3GDgvL1gMMg9Rr4Xjmn9GvW+hLV76L3q+Zbj
K6ZC3cJCAK1Df/sJRtfAYbZnUCz0ijipJjwTM+H/9KL3HNrS4Ab+cmefb0ZL8Ifu
N2RFRpVDgABRLyWPgaV6Qm/BxEVux069fSqG0cbi0Zmd5aJ6s/qE5cAdLl1X1Kdt
REKN1TliaTFOTyCrEkVOSs9Hd5AuOJQ7E8hAW3Lr5aMRK6dVsexvBmh3DNOI74W7
VUH3CrKalc2R7p2fqwbPyQr/vxRoZ4X/0MU3qY5DmhFLBFlso/vNUQSUb4Mv7Zsa
D/aQoCcNWKdlo4C2faZiHBZONBwgQSfypCTfWmr7Yz7fy0VzNilReejJsLcJoRL+
oKNt3VGzQm/Ksu/cKt6hKKgl+SLzlmDGySrpbb8/QPzELjEOw13RWdWRFAy1X1j7
L6smLUkcdoYOB4SaEJ+72tHHe1KBbrIxMyTSALiBPGwUcN5kdcgMYXwMgPKnBdrx
hktWvKhArqBsBvasDRc6MA51zDANppPp586dOEr92O07pemxXvmjxRXBJka1b1Og
xFTgJUIcgKi8WvUqDQIvRXI1R1vwAHbTbO5cIJe96WNWkxL7kcsDCueDx6syMmKw
ii9MZ0Joc3kqyf3/x43JlZuUZ2ovk+FntCl64wUnS/yoA0LknzAzHvJg7oLVji3M
2HwdyW6hKFnDUDFMzFsa1I5IgdqzAFm8nEtp9KVOUOAFWDkQF8EY5e+1P6VSdzoR
cD41PZJrWuai6rkQSnSjVuAvoulGTu0QHjG359UxPzOfY8ENYSxOdiUde3MzY/f0
OZGnkLOuN1tsFDF++jTx9ml1FTdnyXWzm+YfIevsI8lqhTZaXlzfEEPzGyPi1p5H
Tc3mzfqqiHBgu1QBJP+NLsY5WxJjiJ770nsPo08XcD0ZakBzW08jjmBRTkomhdQT
08wkxtrRVhLI0ByJ6vzNgYNffbSrCtrFqoUVRXh+wNuPeevvv3+UaLDKPL6WqP2+
C1Egaqt8x+zjThvdzkkijrvCyKnpHM4il0uLTo0M5zOngwr96nEOb+6tbTPJ4NfH
oPPJNZ85BpdYa0S3QyT8ZEN3eosUFgDsxg0PXHKTBxXqNAHNhS71Z0d+bue/R8+y
FT69kbMrdjSv88PJMkkmhP95cUhNp34SsiEQWfDDPILv/UJ0708sUufEKXldKNeN
PwPdlV+gGwK8WPw8cpd8LKeIDf6NOBcSoJHUSB66QHB4bS10n6u8IPA9aoDiKZI6
`protect END_PROTECTED
