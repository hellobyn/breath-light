`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5qli5gVrhu/LVW0iaqQIHfhQUaBIdvxPeeviPy1RFY6jmQ5d8q48kdXRlVWAOCKd
WRhv6SWhgtGDcLxAUmzz+0rTMHc4/Cvg09yP9QCNw4P8KojqzXfekAdJ7gLpkrsO
PQ7MSblvBcWoMG3Za/F/04ieid4zP65EsIYqI5D+WpQ/Z/bXBVlqn9m35+2C0Ld7
aUF+wblsWxQ3/6HsKw7vtX4wWJ68OJzS9mFfsjA9+WmHr5VeRyQi48RjJOtg66C+
6C49uya7blC6KPpSNC39Z5a+G8X8pziA5CLafEd8WmgDNKOUp61rEa9x8C+dMoWk
ZfsX9RtryFnNfohniiiW/ZuxgIObzF6bIVWkcfSWS0Sp3H383/lykohtnJGxqzjN
NUPNSrH+iOv7MSU5oQGTtWtzgQqQWK/11+u8lobb4EVTRGUbYjlFcJAxIXrxkLIY
b2e4eJQPOFWnUzjPDdrwUcx3PsHDoAKrLvDGnR+uEvLU2QD+fEcgLtGLU0O1MH4K
3XQj9hqnP0XD2q7ZtJ5pFiskVI4jmHMxi2ScFWAS9qujxrsz80Ds3mimbT6qzISs
POptZ38yAxggyMRgdgnq3lkiV/7fy457eSWtejM7CtxpliI0gKs1ks7tFiRIlFdY
VY0bbKcIheFS4SbEJ0WH1q+qCgCFA4nZE72QR0+zKQsGZ1OTBf5aoaS83GXFcy8H
VeCfKIL6UXvSc/6y5PVvhrvgznwomrwJvISfJh5hs/tO1DTfgz8lh/qMUGh2Dqx4
dHSUib5tuzDvBOCAj8UtWlC4eusgqrgTb9ju2yddoHfbkZWRp8ouODda8XrbPCDR
mOVbTBaBQ5vWX8atWBONS78V/By9PNWkaHPjWdeHVdNYUbou43OyEisGLt3wjany
6KUNewYwCHmj8t/hznanhqCq7nYmWrfJXGmqR+1Usqfb9f/JNbDYX08k25fD4owD
pGNfNLntkWpjzbueREcK6NPSDHCNKrloy82l75gMTuSuimJjN8artZUpLn1uNa34
/Xb+TsDMsy+thqVog/GZ+Ty4kr0LueJeaPMv+E6ZIy/KBHw+aCYH8vVVoukyS/il
J+HPuLhCU23p9Ucfm/tVH30lIrLGsRDACTjiAtqoZ44Fzy3XYiZ/gVMJMHuEHZC5
kr1eT6tjN7vyj58C97KFsajv6XE1UVZIyR8j0puzBgBxHdwUSDyJ9Yfy+0qPiPuV
NfFtYeg2hovlARIAYw6kHnA2Ppn/bClaOx/M3/+JIx7Uzea9p6rcPHVRw6FcmCye
GIlvNG8UPZdTSMpyBPxw28iBK3jk8PlRcnh5gZ8xTjYsS1Uytg89XiySAcYhR9Lb
nX6uiRrxgxNmz8swK4LP8vd7M1HZ27HT9miY7iW9j0gmgsHY7uTGDTbciRWHRI4s
vZwWauqoPGyQIfyBzyywOt+BCxvtgwtEs7UTvrO5rZE4HomlD3l07Zs3Xw58O4DI
jsDWF9c1XcS5uP9yhUDkM0Q8iYOJ870EyT05WmCdl1UPaKZL+rh3g5KLJuQo0fNc
nNInn2l0QmzOUi73rPIwZlOmtVjtscWyiQmdZ3tL+LOjBMiVUs1Ps4FJR/VVodwj
6PEc3E0ZQ5dHQt1ZHYAnsNk2D9K6jeRu7AwUU/8BeMu503aO4d8McLQ3okMDLVBE
81e+nAwfvt5rWWxc0ns2XPK5bjD75EpHsYfX8Ruh+aroLtPSrdHCBJPTQ2xRFiIb
/S+5GvjBsCyALHRBr7U8M1lNxEJWpOq+r7jx0yElW1q4+MmA/8YdaaXS1dg5QGKi
kKJEUyI265vD8N3cMiy6aGLBrHV4QgsF4MXSjEmD2X/m8lD5GAuHvyiDAS/B43cf
SBfba3MQXjujtDnLfrhxrlE8waPYRoh/owOyTZlmT9fv0g+fM9tNUvD/kcWgsrdV
fOAcTunXw6JTnRYxoK6z8OauMmZW1Dm4h7Kx/KVmz6SfcizklJ9ehrvL8dylj6Pj
RD8P3TBPSBGqUD8tXZ6W9w6MlxAiJQPfDNK6ABXa1CCcpN/MTZ2bxcZSQOLBuBpi
QoIi10QldnMr5pnFNtF+/YOvs79CtPYEV5AhEAY+YXr+TXgSmJNhgIBqmJQWa4GZ
TSVYpZANnhXzk1IyGsZP2jULMw+A8qR/VgQEAyE7/kdsAHD6X0/CriEzmQsRcYMv
7J556bGJdg9O8OfoSYmuVjxKVsqC4vc+Sq3JiI1UYjoUHSSrnGdx616p3kEFZ7yF
CF1OEsIsfDugsxKIWeuwU/1UM6En0hYuAS2+hIceWrjakRW9j5Yn+syEDa5UVIDg
Pcb9mlxW+dkFhMbrqSzl6jcjvFUAENX0u0224kFAoMZEQD4T/ZpPaUMQa0bKlHHF
GSFn1OpqBkO4VTR8lEY209crN6A8HLSoc4ZVDsr5vF07zv3YX4vvePF83Ron4VW7
YvcV6xUvhVEhZnzxJxgJTVu24vQesxvabiIkGmJHSm7Bi46gudx4//wcfpR6o65l
Fdl08FKRPA7oqTbG1iTvY2eEBpca6NhHiur/z9pwHLaGo5RNwm0MOtG80Tx5MnoO
z3mIeh0n9fdOiZBCA/YoTPGyGFqLVGV78ycPj+R2Nil/x+ZnTX1Wi/1DhM+FejzE
Z5cHLVYlfjDXI5s9kQ24QxSQYb/yRulPYtPYeKLCEivienbtJds+KrpFUCqDLyFZ
VPe4Apewnb9r9Xp4XGacQamFwMALyOO8CDc9cQft+r6PgXoxIH0TJX7961RRl30m
9cYl4NmUlHc7cm8FOjP+9CgWjUtImJYr6KrBX31vT0mrPKM4dvow32KkNy/EZVET
OdExfrTakrMUu16ogDSqXRRXVO9bwalzxBiFdHxvYcu22T6fK2nZvS+fg6HzGOFM
iDT2EweTum36a8S5VTB30qvGnsqIN492XfGygjLEeSugTcdQKnj+PgfZSYoxzlva
XS72LId/9w3I4sPglvfapr/oa4MFmT97YMFmWyhVLizCb6rr0a6Hy40hGFAZJmQI
XKdyf3/InkVbU0padsA/+EQpxbCZPK8YFMiH70iBWfSMFVgKgWbdj6sj6fG1iKia
zm9Lh8YQpOSA6Xl5DkmgvA4TTfnChrgi+ueUDzmWWdnbyiUg2Qu+pNOSC++o3xWH
1LBkyglkW2jAd3sXkk6OgFYH/5lG5kyAvaBKedIQkhUttLd8KKQoKoetLZIXeT6J
VP1oU0eMlAgG0i1k9lK/ZoaPiDiK/URFhZJyuzbKV8UwB+wEik/xAObRePibX7Gm
654shUkApSJMLQmi2X0g68V5K9CEBdxTPtPGTrdQijjN0RtnEaQvObjYexu0nCIH
nvJeZJSlVuSVV+PDYcjZVkTYY38XtH64euDI5+9lL+mKWTUIVluo+hLeDFNFZiuK
QS/ZFXNtfe+vPLgvrLsdSv2AFhwIfH1jOSAcRkHERW/RenJycmDcnvcxef8tgX1h
anv3YVZA1qCFYL84eqjm5rlMj0FOjHsBx3+wKsdjYaKyouOonHbw5EB4ZvWcZjP7
q6nNzQdaTGdxkkrFjSW4BbGbFwKpz4337ht2ao8Pndbvi1WWCqm9brI976Maq4os
WWi7OhQ+QJPZR3j8AmmvE1UmzhGqTX1QqG38+WvRLiEBTSQPBd7uhFjTvM7bZofN
ggFM7UPwbiid5Wf0JRnVywCdArR+/YKxyM25K4coDxmXhyrij160HkzfgRMRyY3z
SntfQVSG0jDMh3PUxc+I74Umvgd6oRbWbCoqleE3xvbmxk8td4Aa/vqyTHSgCrAg
hhR6mzgAfu1+pCr3uCxKCSnlhB3O/VfwY2No5RNQGruD2ErzcXcVrfD5JBzmaATf
29sTDpqn0tly78pBxdUbcQlKWI1odpyrm1PWbeE4S0xtkQyHrhhj5PldbqBqkAOE
dE7sqtaH7P3GxZIpMpv5W/K2BOloPZGSk0+f355cIZaFq8u+/zelqx/eHiaU06z6
WJDmwpke1OfmoYoTKK/TkgbwxW/r/tUAxMVKilUWfI7rueQ1+GI3riPu1u+dt7Ij
8iv1QfL9r37QIDJVX/5Ko8uGLMnZOaTLZUf9G0TDJR18on5N/FaOBcLlT8z0vs3z
IHsLf7e1gfYuYMinsc81k8OyM0yaZ+y2JVhXOk/NDcu+TA3JWnrFwkWZbHY8RKI1
VA0qUWqSzA2KTWoktK0X1QGLqfSerEp3TBcfRSuDyVcB8BZcdEmod6Ec5BeLT9Sl
TME7MhDm7ac9q+RPQd38OpBl5OACbDRjo1wJvoU8i42jsVRkDZJ/QZWs6MP4rZMY
SwRQaxS96YQgUGZBqhEt6DBXNUqz02MMQlHNbQgn5vtBDuYvhpaxFGGUsiqPoqdB
9+SmZ/W9PMKZjk8RCpZmuIfUTah9iYoAeq9WgVfOTqfKftof/YUXcFXKat0xxenU
9gzgNDBz0eJ9LzOP2pHHYPJrUdFtK7ox4nX1ttAPzV6wvcPl0+YSiotYyr1dTLEJ
hMJWvCyu9XNEAALw9jfSYC4mb6tKISsl01RDFPEcegRb03Nnqq0+9EtYyjGXQdZB
1NDcu3naQ7an0qu9tQVGgf9FgETFXjrTBUHT9vHlzBiHTPq82lOwFwrMcI1peJad
olEVyeQm52rCHfbSz8HGW5X6gTOPwd2/YHXCmt2z33pKMsI1j73h19PHJJCDd96w
nczuQ8N9P72b6Ya9pnIBAcfVaOsMNrTLv357kEJrFg1rWTybOaVuuP/L7ZPNMgJK
k1uNwbY+hp3kM0rkUIA7exwoFX8wOykW/A/qEyVtkoz/Rv65xG6IWhJmcytM0ALz
gn/SQpDEPCQVRNa7CS5gL3TcpTlxtnYCis3eiFiObvh2p0t80/aySwfp9nJT1UaQ
lLWoxZ5OlICmNJUViMI0Gxpt33AuJNvDJnS9SI36xuhZUNmXA8wsKQ9wIjKhL78u
YPdIF8v/mhwvCJxFgtT2Ga1kVtiaPhPBVI7rTOS9D44ujKqDpF0hMVmybHmvu7++
lcm9QyjEWTRyGco4mG1QaMqXvcq+MkIZHF/8nXazy4asmCR7pAgVVezrLnJJL886
+xASQzGRCrpHQCIlYK5K6AUzELSmrJff2de2N06ToE+eOz5uq/H6kORWwIiSWOAc
3gHIWYBPMqat+0gTCk903wHLwK1SoeQDurOopFMFkRH8gG4Qy+LYdSydE7cZQ4h5
7BSkHKFrRoS++HW7uea+3jZP+MUFBYgIs6XYBbdZeEicaBAZWs3csx7uTTrAH7f1
EehzCe6jDv1affMhqqNmO3rztWbC44w1uH3mfOGeb5SzSABYmsK/4kRLCDPSiLSb
naHk9KYauN4UIZpny8yzWzLnRo3vV745BaV9MfR4USCG5npmiWIbYF4YR1wICXcJ
CWc9eVAbqt9mhGOoFujtiwUIBxXt54pidvA9bolqerx/8/5j78++Trf9GQ4hnn9r
Y3MlG1MWAMWRgaauOUw+HvEHHRR7TB5GcyYwU9yHSrmm/LDdmsyMHSqI9w9Xy888
wf/T+pA3isbc/4MfQRCJIsvDhSHG0hlBuyTVnJEgNsqzQ089JOB+6l5C53TGCHvd
QsHBdOV1nB62L+0rXo+1CJbC+oRfrhHX/zVaXQk+i6GXf0NyFI9Xp8KVjwcWzGtE
YFlyBkQVdmpXU1ie727b8hc1+A/piLXcr69sivoA5V00DeOGKSlPwqsXSwmUAZBC
tHLkq5nW4MQ8r+CnzFpSDzdi0A8WFqfat8dwoO2qtqwPWL4z8Vji+R1rMaduwMyN
cqYfRtLg6p/5MxXNjsVT2bASJNA4LP/7veMHVE+h/mvHVMf9coo6HjaThUJSdHqA
O7B156oX1OJCs6zmXBcssDW/VNwZ72w0ZC63e5WaCjqMiNaj06cCi7Fg8MyMHT80
+pHAdW9ZMiysUN9/Bm2oPJb+ahLZvF/YUmTvzspmPLXEFShPdBmjYI/b0MRyH2iR
q9LxnA9/Wk0jIfXOs2+FIeFTVz8M9Y+ov6big0NvNcbb1EqpkT1cyyrYfv2Vw/AI
IBkkawaBHljh3tGCTQ4y72A6+w5QLlULJArzqCeYI+9YHwlL6B/FaEcxPIJWRzCk
BrYMFh009st/B1gzxxMAnacdTX62b16y4gRoYPty3ws5Nx1CSybYdM7TTQBJpVbV
pqRN179dRPBSuxonQ6bZHhqb3E//l8pcooLhzndybY8S6aBmb+fNzFjgKkfUySez
rJXasBfcG7ybTibDmr8k91adftmSQt25WH4abkMMaFVo/m8zXUJZ943mWlcYvM71
crP2gwlxpbPGmUL7PY5iRC7756Vg9BK/uBffbXU4w8fm0nvsiDFo62PD6rKGsOZ2
l4GyS3xBm8S8SQS7HMlEjeOSp8utrvMXJFpqUM7VroSFm48hvhsftSbtB5QNJslu
Ep8wLlcMM/QmYTD9Wex9IuXqQDc5BY3gbJQgYS7nldr0dywXgptVcudGsn1YA3M5
77bDeYblqPa5PZrz3nuOvxapEa1xqAaJxH51E+ZlPD5t70wQzZp3zU1M2d1Yt0m8
Zhu8bHhpOmzVAgyCBuRTbiare/6l05SxTM88gy9HHaaYFvayjbMB2g4rrPjLxUPZ
YZLPwKYtA6GvULA16cG71ey5odj2ibT+ew/jLOutA1QGUBfrw3Gkt8l52a7S/uSv
KThNo5DLTv/fGBf38czNofQ6OFumcc8QTRESbprB03VB7eKEwYz9XvyJRqI7r9pZ
yYXhC8dKOnAbdkff+Do33U6wzheK7iBFQ555imS5AT1jUZJTSXgST5VnK97m0H41
UzHABrWLgkqbMJF6yIxxD3qBPS/e4jETXZGzGgvwOIsSL54V+emCQU9czN6BezaG
j7MtW7jtagTq46/8pZTR/352YbwCPtERwoNAZWfpeBeDQxMZdzt9HvX5qi7x7QM1
bNCXMG0j/hzt80VbgGKzvaovyFttOAXoSIkmLRezQMjRHoXz7r+IrwqHfZqjOF9z
B1ZHTkTLGG+BC4MRFihT/vBO/PTmvfnkp/twwCTGlBhoRKnpMZSKWZ19MUG6wbK+
dwpQCDYzYYTkoMiJ5RTJrisusTcOjpWHc6kRj/GD+Lf/E+bpAHUzNQ9eiM3o3JDp
cy6erVj8mQWfdRrVoJ8JenkjPElD+XbQ8CmqWzJICD9XAINgU6/yP3S3xtddQ9sD
0WDHfygeSBnwomeRrD7Y4UACFUMnERSjDYSm7lVzZKPGcZkNbV6Z/u/csU8Dcbom
yyBvtl1SCywOpRuLz8sBdd38HuonCijQwSq8L10XFd0OaJztypHxeoWqOPEiM1Sb
EyBxTozRWbZW3d1+hUosh063F+M1IDFd+uRMaO/DQAXC5NFDMQlJi9QTV6A1DhVX
nlBRRwd3oRIs9ma0JMK4XKqpeAQgY70h8BIptkClbtNiZOSuTPIB4J8k1AbQ0wTn
mHo3eOIWgZQDu3Wp6TonmFMM+QRXIdxtLWDcXb9o2YDNcRpvENbkChrbZQlO7Tex
9Mu1Nr6as3cYUdWfq/I5nSzOVLM45D/E9o17UrliXeV/pnudNCe3yYZxZe1r3DbY
VNv1LJpRtuOFgluPXQAFsdJtloE0h3lyO4AYu3CPvU7ifeI//ixLyRkpTv5qyRAK
3tZaBSUgvmTwO7yk+BHbcPXkMsaOTKodZCvZK2lp3XDwRK56L8ahhySJmEogUJ/Q
l+uwmJnXBwIw/b0d3dxF9Gb1EDzIkVJbqxntypnFUP5Y/aaxzxBcl1r3lE3LL87f
yNVtxFjDgFJ2akFuxY1P0J7s0XHfFeiBJceXEH93smlEr2hVF6tLFS1Knx/r7leZ
3MMsLTZlpDgsDp47VsVYyFxiHNiYB0Lp8VtjBkZOc/Xu2CpXMuKrHup7a7+JKP/d
zHdddMdbp4afNMmKnY48yOFd/KfBDqH60xM1+0GniNXWdfiETmh5RD2TJb5M/DHV
aYcUXKicdK0G7oJ8PspMSqO/ROO7c9nzslHgTkAlNYnZa9vQAlaBkw97ZFrS0m9o
Rc7cy45AsNwAV7io4H8NyyUCatN9wDdndVNK4zIh2+hzH9R4RaHYUYnfGhkBdDcp
efu12EebVOfF6aZqrUs382d2QRWc2pP9hcwyyGNncYPeDcB8QdsqPLK3TMkXxniF
8Io5r65AGqbB1JRwGD62I+a3HH7RG7NPUSDffUJj4C9/cKll63MXYboTsQyxHrxR
WCZfls/f9ON4pn/BnZl7nBghkSWhRxKolfzxRhlbPTz71PoLKeT/lyd+uX/JXHt3
z+sHw+jJeuKZkM6qCi9XS28xzAoY5VE0gX1+ivNPcPy8PF2lBOA4A8ZjbcowmoKJ
7r3KVQNTPqLR9JDpx2LZrwYdaWoQtPWvFy5SE2k5OowZ1kwf+yu+UNQTcobTm3P8
/q7gcWEqjIrP/zNkFPBaKtcHo2eBmGQxFjEVZlTCv6PwRNMRv+0e0AyUOz0K+TtU
t7x+FAvJwg6Bip3N8hHIzP2RUjcxEGp/6xWEQkZvVAMDDIW/kCgsSLLLh5M5YI6H
4fscC7V39GAKTX1lW6as36d93gzZqgJp0MP2VJHfFj5iTMrjWYdk0BASR4wEO0Ln
aQhseAuWzhgrn9RJvL9iFbfx5FAasj5trsqvbUxTAdCuhY+i9rVjKDAY3mo81BK1
sVJup6vrasfmxx2nvYiD8HxmD3gEKdgFCtG8I7w46E0bzTDYSdzvEieRyPI+Fgm7
9vL0RYj2tVk4MX2VcvErXNlz2BpuWCRX1PGABv6l+Scflv8g4vMUYcM3X8uaRSfi
2/lrT4CZ8jLlJK7Sd91HfMO8gtYxQGZDCqrs8TSS+eaFVNX1BnX5Bx5NfBVHX4xz
Cmr5En+pVCh2mTyAzA4EZIJ1XG1sL6eHkmfFuMKuKzVT0KgWIo1l5Rqj7EPdk7si
GLzg/nCMwkTNCc11clKy2gLfc446lwVbxZ3X1Wf7z2VYIxaNGr1jzK/ItXA/iy05
iyguscJEOg5u1+gZqHbaLYkBwag7jBQV0OsyztmVDJIq8LWAS6cHpYSj0WNA6VSF
lHsAo68S7Vjc4z2FTSnAcbVy47x8Af8A2HBw+7CK23Y0Inn9/VJLjag3az9IvOq0
yHHi80nxDmKVF6ZVSPUaFPDDSoZmhhEJjFWEK0VsglPfPzUoUC61vNvRsNvQEd0R
yrpBmyQrSUe8sqLgK+G82/uufUu8hatU/do5bGbo/L1+0EG31ytMMe7KykWwvv+q
ot0mtQ8OFE6VKqoy1yeC/Mru+WLYlZ+Ld1TqeQ95D0Z7wDNw1CLh6jF0mLwhtwgI
xRdmY5Oharo2iMEbQF6m8e5hDauPmxXTeR79meQUzrZ/JlzvHInUaVVf6Elbq/c5
LT50z1jEW7yIyVQGVeSg7sUdtIqhd3gw2sKYNjV0QmTunJokwp27etlKrv+k/Nhl
bqIEy8FN/giFbZU4htUCVqtGXfZEgrf04LbN8u5RgsowKMhr8qKK2ntaIgddVdRm
dvx4FyM2rdNSWnIPsrBxj8U5xgn/S9xbQUlH0MOCBD38w8hRLhhUA5UITywxFq2c
qKzsWjPZKz7NYjUwy/Nvdh9to/N5rqhts/J7/UipAeBtARONsWtsYn1PPZYt6q5A
lXxLTJEZu8JJ4yV0NRaWZnWmH/zeUcL1Nf4hffwrCPmUnHqGe7pest76B23lq+Zo
aBEw/P8Z+PQWGTu2lDvFxyghwFCx6cxAlGHBnzZOxQkrhrhH3pgaKe6Ybzfurmqv
`protect END_PROTECTED
