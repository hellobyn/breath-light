`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wO7ulv8gsZx74dB8H38fjDmYcgrCjnoKo3PSp/YUf9riQW7ulAf/SpGJ6OY3WlAo
XhHmAJZgKBDK2117aKV19glHPffSooHfRJM4Q+JM19cvIqBFJIYIxzpxcKnDEmAv
rIOuGbSkr+8q27LCjN/ptCJDD+5LD9tKzGdjmBhyYHpUOqGr+Shvn6U0bODidgYc
fIa7V3WtAm5PonVNC2Oli7ZrLch9V5tNc9ZVriOjDf5z0Vm3ktuHzITqx0yrpNDW
iQwDxCtkEcvgIjO1KXOnq23YBuFy6KMR7er0aHYMSI2o/pvu2dJfdDzDfJTYMmwn
IibVnfzl2tGdzoub/59rlu/JeH91n21tb88VK+hP9BloNOyM/LFNEYGmabOvMsmk
X1IsKCipBIkccYYznvUBlk2SUN1zvbDy2ZKqTlM5CGjJJQ3S4cPATwqnGZL7TtDY
g7fPQ6cDtC8zfxF6iGG5S81XTk1ayUwi9OMA/qWgiTBHeveWM5ulXGyK84wJX8Dw
LbjKGv1xr/2+NdxEgF0X1aYJZc+NYeHHDEbyDvvAXr699hAMam4jw2aPshUYZaUe
3Fp7k9tEvhg+DrhbxsYBzGJYf75jcH8HRboBMMbaKEzgXoQRld5rdK1ARNSnsqR7
NursP5R4JKkdmRIrlHHB3g6jHhDKecs3iSRRHxMBWTBasBDEUxs2Y9UY59uHMe1R
klVG9MBwaIBW3MxzWnKb2cpAyBdWFVCvZUMyM1W90pNCw3b7Byt3eFpJXCveqEoH
db2DNUxQxBMkvwnCwEpIrjbUkQ0lMb98y8tmzSkiZKqZE4VYZy9S+7k0SeYqJ/Tc
s2ELkoqGy/uIV8Ck/oF9LWW8biXmxkPFFofmcKd4PDLc66MZHQHksjSZMwLoyvFm
Dwtlyl6pHg1mpSKzNf+xUa2ZyURNwICgIkLep3o0z0hOKU5dAtEvujoZryyxfFfi
DLjReMjQoLpcLLx0c3U10ttqWJXyQ8PwEa6YPEqF1NeOpmwsNLF6smV4/J1XTz7S
pp3DAnqKio+t9txc593Tkw1QfsgRD29N8jXidbLBl9jYopRYs6mXSNYEFHk7aVOI
jAFDOPCcvvlRq2JyKtJs7ZpJkjKdgR8ltTxzwRnZAt7Pk4j3LfUfsajqDODieEGm
D4JQkGppt+05AIJRy3vKDL+aBh5Rd0Cz9NrB6v2ChjM3YwzWQFO8B20mVVyo53d4
4TW+S0kUBO8TKBNEaeGxDK84Ba4ux9vWWjfPuUzXAj069BTxJgC1zdLGIbBQbK2N
ZRrXkO93AkC0o5nm17uEWKl5yRoJmRoh4IzaezAYXB2lat23HcfoeBJkgVK46yYF
OCrlihNPshmDXJZMA1KdLuDnMFvEDtSItrJYvammy9BxcgYBnJL2EY17Uipa2mt6
WAbZHhOzzDzDwkgrwGRMR9owukl9VQCK5LPWWon8v3Bvm9zEFXi7xo/QQfKMcSde
RHgiJ8hpx2YAt5tgPtTQh0QghCm2+RZzSg6Ndy7RM7ZHhbgYHcI27+NqcZaCu3nn
rnC7xjZeY7MPJI+FJIgzyOEhpwA6Mn4KUTDGjiIOwCEZ6XbzdTgHuMO07MJGAMje
+avXF86iHN9HsyL5YudcA4de0BhwXiT8za3mxS+hPsihdCDlcyg2GgJHzVSkUtkm
FsDa9u/wDmz6KqeTrXpdUFc70VvEO2t0zh3lsBzlPm5NG1Qk8v4AywoWqaQXrVct
RPW5rnsJhTRENc3wnQtauAjQA3fYm6wGMHfHuTTxJdyMFw+X1PjxYuUWzqv/WNHb
49VEKoIfF7ZZ7fDBlObV3+dI3hcFJe2kfCWbEnZW+DGzRcpW/42IdSPTgJLz2CaR
OZH+GVjUEmzMtzAcqaNiQuX1PnwgrarMfYXSylJXwzWHr2dnDuU9vWOvYSyemp1G
qefDkvg067zpXltDcLC+I24BB9XuyFS0Z8Ipvor79Rnm8e1iDq31x+gnqCrOQZpd
u0oQxlKH3sCWianBQ4GuEKHKYkwh36ly00Oqw6fYY93d3MIDrux3/pzZtNdXABj6
eLQPbUAOehjoeQjY+rtaEWTNHurtWbdRUIFEX2rIam5TcvZpZhDQK6hngwq1SI0H
Fu1oVEeFTzO7ZJZad2PIUe/9wjNo7QTbr8rF+Xity0P8iRO8e/YZ9vvd2UfQCYY1
aaVXV0AniKAcZ2hMr4ESUxcsfA74gzuM4+6upldubZE/BRjEhEhNrgTKLzqLcJsW
AyLhyHtEAiIxgnI0MfwyeZohghjpYpbaTXE8X9Cm5JUJxBzQ5J9e2Z4SXRGNLAYm
2v5Rvi4+A4rGjh4naq7kBJ9ULt6+AYU5Hu9p3/pCyhIIsO/cMIV+C/32nM/JSXO+
bZEZqGk9ixkxmqe/MFXFHAcmZP0eP8NLZYgCxkdzLEgxla7kVP6F1ry2mItCliIZ
+RtLsXF69aj8tezfXlWzmA==
`protect END_PROTECTED
