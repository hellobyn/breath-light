`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRFVFtyXaJwN5zeBNy4Kz26GK1sjUItC9d423bJw9hbrEx+qZM0QlsCZY5Q/i0fU
WfHOoibn96HySwn/r+bqGavorFdnpm7O6UL1N9RL2IWMbGrZh+yx4oLb8QsB5GKB
4+1X8ROaQjgQcdYFKEnfznSuW7WYwKS87lRO/Q0XXn+i24SN2zfFIULpaj7mgI7Q
7UEVKe0csEcvgIV3OE6WxrBxiCiNktgG1qI+VCC8oWmrmFDI/MlvZHjDAbTmyVHe
D9+4nee3BhtT1OHz2jdraLqp8tL7H+1JeI0YSEg+yCT0yovZzycgsMJU7x7GOpRH
hNJELxXFc6w561l9oh2LfJQxikNWUJ+TwL080mZsJCuk4oGwJcuSfiB52emGm1CF
MH2vS4odMHyS8SES2Muy1rPHl6hgJQ36WTRGkOgRBCeAsDM1FWjVHkumfoPDNX8d
pIpAcDV0tvgLCklnhLPRrc4uHSOSwwhRrR86ThXUBm4HSY+KSGfymTiei+y+/nzq
C/siRIAEgq1RzlVGn0RhnlCi4uXYl1am98RygwEwQFvD+V+TnooC/ldR973qfZhd
qW8WfRIEn1/byVeh8h10cRdNq4MPJ+K5voWdGlhBknpRwqG3SHukwfW38CXA6lJz
Bk/+X+hnRWJ7ior7JrMWoxQfHsI+2i68VpShRYmzqwnLs9usydR/sk8B+iwKBlMf
E4ke9isyfTdLobAlzNz7KUS/fSrR1i/W4TtQY/TiD75dRz2UlBaSkC/caUKeNgH7
ElVpmjIEiEdhqUk2DUGQRj7hwcKZvGSwEmYiTE98xwDkBO5Bj4dACFg1/8cv4han
8//B74DlscpIl+ItOtHOczFM1/DqoVnEF6QialUBud1YAIbaLR4M2UHh2nqqSiU4
BiBgLjlr9X/jX4T348xkn5WjGARr/8ZGiEgy0bqlvPYxhI7XkuKEWqO7fHftxLYt
k8/DwE8SHAFFybZNvpvtf2SOKchj9ZloKq4xbgaKag4/8PkXYRHOdTkmxgDQYRJI
wRB/bM4zhDToMYLECsSMmuDNc0YbWo9HjdIox5MWHuPtASnviDBKWkzFksiNZ+B9
EQVelz5LcZmXzwqB2GuSX/yHaC8yqVpk0GILS+MB6yzzSU3rtV/x4ToeGzxXjqLr
qU7CbZIUZfCNL7Ra5VNC1VORWCDNbmeErvwRHpEpZD1BU+jrAdYR1dAc6iL6dezK
vJaQ6qZdNBqY6zNUr0Ymo32oTsb6PB260UnlqytKElWR2scU0AFgrVZbU4gno+jM
lbdIkvA30XRTNEURiuCPg3ulikm2Vn1IxD4Yvrrk62ggxJgsYE6mCogiuvfNZa1Q
ZVfbyKFu2ALb3/2Wbl11aORPs7P4Z890lTXtSgCRFo/kpMYgZX6ny0IfuDw29vGa
NG9ATGUkdE96GJoIweNf90MqEuTy+OyPQoFUU5zrpkwEXQQFhbkglVYDxjcF+LkF
`protect END_PROTECTED
