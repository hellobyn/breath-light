`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nK5AOWV25qEfued8khkMTrVtA4yBNOVtU4DWUbe4xXaP+NKoN4R1mEDmd2RAFC0s
07eylN6zZDS2F1BWk7UE6TxxuSfw9BVvJfTDFfKZPSV9T5wyH7aOay5mcmYngSPq
yEN7GU4cuiwu2rrJUlk6dBvsYYYCXS2Ejuy+ShUGcSWdQeYxfwfjRz5pZDqLPXnZ
V+EDZhc0U3idILTfOG6c+ymJONupNhEFqvkMqu9ocrfWfIGXjsJRvRsNV5eOxAJ0
kz9qPknGcpkfc2G2e91SgRaZL1GELKCkVpNq2s+qCr4vEBcSB1LB9yABnCpPywg/
asEmhHzanJG6t/MBybiStWoxfkZjRv+1hRpuY1+jtByFHMUC3kvm0D6sYXZUBlDd
qD3OobRTvMM/y7e6xbJEP0Lxd5XMxAly0KqdGDmyvxVWvwIs3/VeOUA2Hfo9G4aQ
owYJVCIr5sT/zeiUqcMTnM/zhkHLze/fbe7jC3dBobNl8rYruYGNuFly64cRBKNx
AIvSMJTSag6bvwWYwbQvUfSJbT+8C4eKIQcdkNl3A5YG9vVYsMG/8lZSvGvdFV/O
rNPmTiwgn1yBPBcHHTP0ihuHegvpVDFY1z82VJEnbwQ1iK4YwX5lqmlGWhQbtcC5
6UfM4ekkAzuaXfFzMyyrvnAptEkMwbdy1d9Bty//PTR+2KCeb7iVaigTKGgedoj+
VJIqSpbJ1wHOKeouyzL6VY1H1wxue9Gz6WMe5s6PDH4Sym6tvWhW3MKIw1dLW7La
nA/cFvDKw9FLbV5Po61aQggtdFj0gFv2GoGcyQCxkstBLGDedO9hNOO7qdN3GaKF
CraLkIyPIzl9mgaHdEs9Vwt5ZW1ERBrJLVDjyF9vgCR7ogAx2NOAqBcYmmLGcNOo
coiOVsKSYb8CbNHqsLCP3MmN9zjTRwmrHwPRPXnjXQjVbG1t57Puwv9qVmu+bfw9
rdWhYyKxBtQSlQ7hYPwOBZDmd6InC1q7q76vDrzwtSQzrFoa0p823AvhfU1xlM4J
iBi87n6nQ0k25PHvAEg58HtvPyfJssVMK7qCxl+V8EosMDyNPAHzP6FvN1lPrIDi
5S1EVjRT+QpKq6Q477f9kuZk1dIpvPW2BtyJ9ZzZJvEX36kOJXJ/arX0pEi5RWif
pNo1erYJf9jfH8e6f/8z+ZPJR0SI5b28xIuLGymXeYeuOSyxGeuBmNY63zslRTHd
uopH8RWFoVowWKgL/OtyK8Xh3K9N4m3JTOj07asGm9RUnXRmqG8D4kBC0fkQM7mu
6z4pNNV6uCNtd5JFMsD8u3SX9ecHxpNPxFn9jRs1cVMicOGFUTguBiXOHVuRYUD5
+OCsg5j0ngLgy8oW3w/ewzQ7ipz2F4YnfA4CxNBjY5HXxkC2sVIRB2r10bNq+UlS
4CRy5A8pGKKuUL2E/vbHqR3GvyB8H++fEBrSqcY920ljvNfX7nt40R3HP9hfyweF
ywVD3UfrMFIvVFDMjM+CFnAXXWICA+YoBItY/o0QHbCPG/vj1kAun3jHvIR7rg+u
6nDcxbAEj6H2LK4CYGxy+VzVigklVWwfnrqYpULs8f+FtwozwfZ/FpBhFEuCb9z0
CskWobcVXGGDU8ir0idrLXtFpRl4swd0itpgvU/JLdm02J32UKOxUUC12u5ozLvR
A7z1f85Z3EIAs25czkxX/hYyMXSbkT+9dIOBzCvhx5xhRPnd+F9mkKY0vZxylzPo
nn4uPZG6H28Kanj++7s+D8dcfqkgmcXDtKlcBDIhRZL2RJY+7rcBG4/f/p/hRdO7
r5zI0Wej23dgEdypcj/+9nH46hbYjDRq7rX/F62lnd74dQJMcN2Dc7sO2YtVjutY
Y5nxL4WivcEndc3IQDV32NlDqyGKbWGDFUlYusX4yCr332ETHG7WgqORmKEPIzsx
QeQozw5eaiOarA8wdFKV6i1Nm6gWXe41A0m7nTEMBrKG962a41NQqH25REj8qAO9
hYIizYtg5SYFjubvcdJ72sByq3tpM2UKYXqhXQ+52ZduIoOr37CcqimFyWhIv9Wj
i7jJbm1cvl51/00fNvCbvNJvODh3MwBcWvxKP7u6BJzXwEPEg0UCLVFqj2slbefE
FrDmmSewCaa4lMfmC/pFUxYdWUZZTPbxG8gPKr7tPomOkfdMzdPDKIvggAt7DS4f
9dHF1W3STvV4eXqoKT6Pkz1RRF9RMQaykxV3y9ZkQgycux2PuitD1Kt8uoR4ZIIY
Yi1q79I5ozmhNF02s97T3GfutIzqPraX80DrExBdObR6W2noOXKjsqKT2miii4yn
l6vCAgsuFMtfkkiKxvXVpazaOA+U7LGkvGPzOc9WX0E6WSeO9CIJRA3fN5NnHMKv
dXeSJVBI69kClihHGdTeR6sTyFjNuDLJ/A0Ph2Lj/2gNB1of8OSc/u+1nl/MZAR4
sG4g2sSEwCqk5eQH/B40hTJgtEuygn2x1lFfQGnQYUcaU9TvpXNqgIDRfnAGYNKw
ivNIMPtfF9qtROMCFAwyjhaH8IH+dsoAjxF4ANEVHXHnWaWeBSlYjSivaHuV6Xkt
IOD7rXXeFvKAzNCs0pQ+1jA8oPUQoBNuTmJC60jjVlJHm9VrtJnLk2SUV2Swl/qX
YqOlSvDb4NU1JrOnh3vX4G3638IXw4eCzJiCVfOeCT2UDVfwvj019gKVLLhYBy0Z
iv+1EBr6/SKHfl7dutyin/CB5poG51nTy/XXsQgcQvgU+bAlOiQsFYiSjFAIXfuG
vad29Fwu5ql2klhZjTVPyhPT7gqFdy8XEduhOLGSioGle14gawW/275GNmNPpipN
vthz30l6QqGOSi2jX/gozxqPtGBWZccaSS36VT9gPf+xcHJtFYlicOgPE8+v+Hgn
pHfE04J1FVYwUdjOOIhA0wzoKdpwc8PvTaF71ooRiRRgnATyRsaDIJwv5+Qi+fox
hfQaBjDqu6GJrVLS3z4waOtpiypHETRIZHR8OVHVtLirLRqrPByupj2BipHePX/B
akBJjr7SvcCR1jNFMD0S8im6te6vnjiUt7KdjhnjBNnfQs0NT/1gQpo77BKWXGb4
QmJA8o+0/pr7hXvfJNUUuBN721TLq3chwU0RCQ4FD9noJD0wqoLVu1tUHqHCKumT
rx4nELI00UsAy05dITPkKKwejPiti0FEMYRuosNJ5xEHRrXgY/rG28gHWBHMdThT
qgFnmixSifAdfyW6Z7nEJMBLG9b5u/9U0v46p+amRGLvGGX8U8pMFn8Q1AlinTzn
U8oP/VUve59eIM9EFEKSa9+SUO3rGcQFLhrJMt3s26/+yb+srjA087SLxJJRN6V/
xJ/WxroNdz10ZWZ9OcyYvCMzkULcztZ9+KVkiWKUL60x4wOLcbY1ugRNk9jXfxzd
5nyli0SQHeeZZXk8GgEXlMeAVQX3Avc0u19Jj97SCB3fEhEMMJ9WELXrAwE0jwpZ
n8KRUJ0nnizrQNbahiL2z8rRuMWbujo8QT5HBpY5r1Fp0tscNQnGP4yMfPN5JIx3
yzlvubKBbFx2YFB6ziG5ERWLWhqQcTB/DHQXdWjgPkzBhx0kQcYA4gRxPFjEum9d
okowQ/cSZ2KQCTiVqS20v3Jdv4qgrNaPJ2rtCKMYQd22FjJbZVj2WTYCRfkCanHV
OPU6tgufzCJ/1F81GRLK4roFhaX/A4eOzMiHz4+k77mAxCUR12Mo8SiafUh+8Ish
T3gHgJ24TWUy/lkQAb7TTqDHw7eutRISHgJy+agr7RT8aPRLcoiL7PtqHCW7TqKl
3jIJgAgCB/+05vYagXaO84VepyQsBdrYhsylu2PciPxLnJovDYPFrb0zs4hfYne6
Vuku7SVKIltsMLkRk2PdsoBydpq4LQbp5E5qhkXVTjbP9ZSKDGujVLqTwNWg4iRI
iNAPdAJA6zeZRqEj9c0M/8AOePfcujASvOGOw+f5aiuTAt7/ixVj5kQLa5NG0JmU
j4GPvRjyVPM9Q6uu9S+e9QkvqgM74XBVVPqFp6g/dff5+oim5cuNCl42A0wndNLi
VcQWJQjnf+kR6xlQDtlCiEZSqu2MKHMrEuu28+b8FDw2+PL3rqdkxXt5wFD3yQrU
JH2cD8sLPnLq8VMlyRQlDETsT3Fgxq8d2r/zaZzfAnHcuGCSJNKb+F8Cy+gzKbEu
6OvobyH3COK8bus7MwaZWysrSG/LfweYJrGEt4iZt2TdwCqUMQp6u2sSbZCyySUP
6WaKL2uCZPzGvnscy3aK4Oyvrxk1CRW8wzCJb5MVomhF7WzR55/GgPAZ+I70+OZO
RYOnSWoXG8FzUGbAEoZc9Vv6Ca5AOKmpqVPgkSCHMDT2GwhNpBcCPeef/xl37I1b
WCSsa+mnyZ1at8qbA8KftaAVWv9XC4cegyy8i/b5FKO/nL07Bo2jLYCRhHjni8eY
n+POT1XZFSitG0lWtsKPJvfkIJMl4goJWkb6S57aOxIiQnA8POpvHImbjDp5DwxY
Lh2lppJLiW8kExZVmv0rWG4KSh+fHHUNLIq7JvrA4qFWQv64mJMsQMtgTIdHhbXY
xSSE8faVIn5eqypgj+gd8kQ8A84OjWPJzCN6q8j4EsX2SZA1/SiGKg0Ye8qarkli
7qOLgEIbiwARthSsKESsJbATq0UOEwnPXvkT5WM84zt5+EANf1wTnqIt8Cg1rS5C
ZH5mvzHIzbueZgIiBWubmnshGWVcluJFFmTWK7O5XjAsUu2NWtx+XYeC2uTkt4yU
cI2/1yR0MKK/rb8cDchu0f9BDyxeBNFf63OSDV39j/+7DjTaJR/egK4a38VHjR6X
8VtZdNRTlZIHg3RqMkI+7yCyR7TgkfUXrOcnBJjwGVF08EBEGpZ5NtgPN41soNyc
uFJnEWJf9HLPqVyWgWW86KSl9eFaFa03kW0XSn+xTpgPaEwXTPKEoJL1h9NfE3wX
mpUhbxXHnIiGCcYayO94Udl0FDcmcN7xuUXZieNfUh+ceMyLU7WY3m0yO4P16vMQ
OKaBCuE8y4zRHaHmqmKS9lfg4tuJvUOcvPmfQ8Rh0PTAKClIEe5YXOqjyL8ynpbT
VwHA0T0H8h1YsCKIC0DHXuuJPpvO/qsUgVWuk6rFQ/GurlmYpsIcPgghAs0r95tC
Gg4l5OwAfgSk9FSw3yR+iRCF6zRxK1qsBanAL1HMZ7mFB+d6mK6V6hdNhNKnabb0
U5py+GaeLHHnoMB5LslwoV0a/F/hX46HiuuryL0SZPsekEP/viu/9PXb4nqyWNcF
rox4s7g88eXtkPWSepB8P7/nkijXSYz+eHBCTGttcCMhXqQZwprT1MJgKRWtQhE2
AID2EA/+jKl84IIE8RB5c9FWV71XeyF+63F9tkMfodId9s7bKZFuCFnX0hE9sHCF
cp1SY/Su9f6ktSNwPLgevPmx9emLptpX/v2AcHtTNhNvkIQI0FqrMMz51JS+JqlG
12retZIXjLMgaZQu9G3g1aSWJrzQKtPqw1vj2x2dp0FDd+1GHBemETFsb/Kq3m6q
rGhe/QNqRlzeVf5B5ja49CzwW3sXYaLFr/5N4Xw10KsaYwMSxX5tKBVH1nLbz1Ca
kLqXjwuZptzlkltPynzii/ddkSy34jA7IhoO0WcpE8m7sp5hwAmmb2DmtWD2BWXU
8NVX00qfcQNXoiLFRWjHwaENlV45hDHkEW4ijSRCoIHbCd6+Piv3ohJgbm+oMqHC
Qq0udK2IG6XByClbP0g9tD+bDm2xdMPr+JkF86KLf7uxq/+aOVwCOs5RGQ1rtopp
GTYnv+xYvRfGQtKCtK64IqG8BPeaWnkHf02wSWgU9ZuNE1b6Z6NGkbobnXByZ4n2
gnRK3pqSNqlV1coIPFRXcXqb//AoE07dv5q26LTkzbLM3CvnQ6B+Aj+o7nmapiwD
EWysZLkNlaUYHdEhK3244d2V7YhgK8wq65u4p18lgiIBSG89uURe0NfyDTvpqNsn
U+HoVDmQODRfNAXHTnoMf727pPtilri0U0rn6+yfQfphwwKAAeSDDsrJZqHjQPEO
9mRUTF0i0iKqu9B7Zh5LS6arJgcl0dW9dNGLJasqbWw4frxL0sEM+JvFikwMWLP/
6lna/jNr4ixG3cEhtBhLbrgBXvkET80SNARac16ZY7NbZFXHAm6f8BMtVg6X8A1W
JurYf6cuhJb/tLxBNqhZbd57VRSRDB5QnGpsd7QfazgBH8hwrImL72likGr8WuYH
iOIXI49XdFZGd/yGQBXYe35JzeNx92kyQM+rc0OefIORGBuzjVqtsvP1R2L238+X
0hP3Vxc5o9HF6MOaoML9OXXAOO6NhlbdClvEKCoANQJGGcEgS8uCNqaes7vixTQd
zjiXr1WR3sumq3eQcidTVqG67w3hpUPOz9KJMghCGUX5BlM6DZvj4fTLe9+hfhY6
5HzEqh8i3fthX+4EN4pY0kjuPFaPECfxgz053I4jYdUoRmg8M8YIAQqGkS+DMZHo
cZLztZaNAHw1m7nzeGphZC6ay24ROqoYcOC4SwiGKYO57RYLDYLhFQ8Aqbyxi0Mn
xWzV4tHfChn+gpDEJHvIqveWC85thNpYNPHUx967xUuVITV/tlXsCtp0K7trhEze
C0Qut/6ezEwT+9A1yVgIyh429UTLKIzi+XHPu94wiZqjymXEiaPFkasJJ4B3clAO
XJrsRWRUANDf67P5ilizzeAWzDF4K2PDUyganbNl1LukwPmv12f0LuToAcFH0Q3t
yJnfV0b7EahfC+lswMM6ScVPvJP89u7EtfLeII9o8F9lAUmGDj+Z7cHM2uhDE9AE
khHUTXNpchXz2wEJu2Ju8IHs444kQPTH1ZBYpkQkeM1PaXkHJvwaQvHExFeVUMBL
m8GUlOs/acIRY8L6B/H+vAl8IEb4R6fZnCfyO5pq1dpiLg6nC78kNjeJNu7bbgr5
+lNb9dVMt60Lc3NevK/mizFqIkrCPsMZ7z42Clq/Z1MjV1teJRES0aCJlE/S1ECZ
TJ+kqbkTpPSRqwQkEMUV3Tnh//kDfsX1yVrEfgd5ZmBFit3YY/MzqoyBsucMYAAx
/0QQc3T9fxYYhm2nDbc0crH8uhOWTe+bzbMF3Bz+nBzBZJ5/EV6cWMMVos9Im1wk
P5JI9OlP1TlCjoKfZkvBXoqtDCXcVnOXDCO1DBedWGpZG5RMGhOlDeKieuZiYJzA
3u9jzLqbF3nl43LH8BnZI02AqJh8V6ekKPBVCgWo9IcCMmF2nnG29i+45mJzKES5
wvkAyTR45jDxbndI1G9gXZFqeyitx+bmCaQ3aTaBz4jIdJcxsLXpezDqMjt6wvXF
S7QoeaLC4G7GjBEX/61RJzoyNh9cg50o2UDEX4WOe0oHT2LudzJJ6QC792srndxu
GSNMEyy7HGL+qF60f3l4ZRxLPaWbbSA/Fe3K9Kgttp/RCTYp7fEQ+/90hCC9oz5u
CRSxLzAAzmW8k9gznZRZYx0EnX5p4ulKkh6Zsod8+M6s0Y8Wk15xcosiCucn74OZ
pIF3Jpn46PKoaC5j3daXe2u4VGGsbvxkqUqnkyf6wd0zyTWZaHbtNQ3yykO8JS8W
BqdKEZ3yCoyw8qtQORL09zD2UMkMdj0PHrNGldvE08v07/JMUifSCG96AlzEYc6r
kh8QfaYyEN/qcueIz8xJfGNn3KUqFGuD5Lsm+gxgpmDuxtUOapYNYg0JCvIxQamy
tqz6tFVesshGvUNXE7mqqyvKtu6BPpjFRLTFJsJpyWQqVZDkmS0ukt9V+rfP4dIf
C+6yGPf7HgbEIlq4cEeMMrdKgkjRbQgUfIwQhPySRV9T/vHzdbp+77lfUTEeFuAc
xPNBLRO3sGyuyhFpCHNhevljzW38pORqaHByTRMWCw9QyZIrmHx9ppishxi3N8Vt
kRnazKyEDMaBaCYPawsNtLooERft0k9mDGaE31ckr2P2/Aj4hJRCx2LuyztyX2a6
rYhkSST8K3OxDdHEuNBvEWaGm8RF9+WvZ1E/IGcVyd2fUWAg3QyurTjgrD9tkSdZ
kxXQ5GtMj01GPwlXYyftc7ykFCWQy6gCH+3zI0ceSw0zpyKoSiXqTP5OZTLXjagh
D4JZ2gY4ennRjzUHe1TcJgWnM1uJ0tldFRnA4BQMJray1V4IXaA5lh+b3zugi7Se
QN2Swg/qUQbbbSSFmZ+Il9ibjzJsnMizQWXHPJESj1ioP8mbxWtaAS2mVciW+iph
ZvrMof+DO4LCcd0l87M3Fz55HL1RVEw94XU/PUBPGeYaV2zuoEHNDc0VyywPjzj3
kEV3/f2Np86bvyf/hTWs+GxK+1FJHO0QSvW39+ay+pzGH0PAYcO08eqIyBkkomdB
/f2A5YPB90yBz9hk15U40rm2VPOLYB6PtKAeKxZct9N2aTHtHCH3MXsUnJLfS9PH
UErin7/BqCTA8vrThTMVS+IjJ69WERZk7zUySpa9LVoA9+h2kQnvnJRkMe9VYTJb
ZSKjTVFDgWj4GmVhVmS0bxbvVYjW6IErwTOg/87k/rfNceODan12pslmRyG1u75z
4qZFRU5hDMDpnBs3x3DfYr0ZpAA6u0EocdWL3+u/YL8xiNkig2iUPM9Hbc/Zm3UQ
kSbSdVuybayFr7b8DNSyq/wHYk5UHLsPviARheZRkiJmzmHwQdOnH0T1Muam/6Dv
Zxlo3mj6Q/zDIBLxYX0b+BvraYElgHghP9p1cF4byLDWefVud0J7hi79SNe0NNsZ
NK7k378RMweyVgaxPUDs9zQnDwKYVuG/PiopjMR+tMfi3fwOVL08NnLg3G7Q1U6i
C7U8bv8vVHHE5nvB7GASqoFJdTxVvtc1hp16UFH2IPhniVZPojTX+GSNNbDea/xP
js1sFHbwucRRX2s6tBotHolvS/R/vtOr2Iykz7rIBcPc1EIy2+kCxJFwALCq4lrN
E2qn+DIMxYYwBCNe5gAb72mK0MKvEe9l57bPyE0jPwuN3CL8hGz7ORTRGA4Sx9ho
0yP/n0zRWGqHw826c0oJmDk91Q9PzgV0PXHoIMfAY7tpGdPRv7Zr42kUktiKb2pS
n3Xj7lir0N44117MWTOq9zk/r5TiMBHSQpagHrJGDb0GQ0vn2qRFLVgfnlKxJpoO
QmYxI5gK5wsWbe416C+vdzSqWnp8QMiMPF+L8IzMxd7fj66ri87tvpivcwp3rl6V
9pmiQhThp3h8q7n06SDjAn0YsLR8zR1CWNv1NGB/Z9Wpyl/HgUZX+QF4ZkOaeJab
a0rsYIGyJqRw7y5cpl5HUAycfZBEP3PLk/TcIB1LFP0ZIPcNyhSebNKzWai07Ebr
8WqJzayTsKEVnY1LVLDrVLfjmCZIVFYvDMlTsXr0khRXnnOX8DlPwBoIpxXs02FI
biNxL3BT9+4KvMhuMmbVTWSwI7DisfCg52MCZd8Yp3vSM1HPnIU8pXWx8qVUwXUJ
kG/2bHyXvhsjQ3SNC3A+oh2tqr1Z2ghmsX7//hA5NY9qPtz8DEZ4ewnzejbAgZNn
hiUQmpVefon1xwXaxukC8qyT7geNRr6xagugsR/FGsm0qR7fChYN60UzPFmlapaf
KfJ1q8DcRLxodhudz18h1cZ/T6VooeMUzY4R1eN0NoiKDXNgAQ9siLHoI48pR5Ki
qmkIAIIgq/ZS8Lc0D0fx7VIbjlJPsXpba57Ka4eVcXPPVw1dWl5QwaSAHFQkws2r
4v5bOqN5ySNo2Qjj7vjcuQn4Rmmwz03mcUP6+Y/AiVH39DPJtjJqEGo/YtQEfBGi
WNMGw66ikkDtqlQnNNZSOTkmZS27JaZfISBD6hFGyFa1jaeGOfFbhCHftTCHKJHR
7yBP3F/IE6l4h+lqwHoSJuTOyLV7IW1DrUsFopBB5bS09neChk5V+MWeDdRPgrwh
bdlccz7jQXTCRS1BCmHjhhcH/U7oawvXDJ9akBwJZ1dqDYNFSlK7yhRz6xVN1y3D
5zZXJATHC4WvMtJtWs0OJVKRSOwCld19Ra0xBMDr37gXDdtflT1SNEWRTLK2BdL7
AS53UyUP57uCPFFZPweCnvSQcz15wKabYjExAG+HO1mcIMYxX1tm6Y0gb41cjN+d
4KfdJMozdqHugEaD+5iL3gWjCxSF5WRFPvp+SYSJ9cbaeBnBWRSVcB7r9LvZ1Z0r
MHoqG+YxOShiE6MI6Dc2oCMlhh1zghGCT3a2ozKIoq3Qur+xBSr+Rf8NuawRKN5y
nHzWM08Xu2LfSD5LtWeTTEYlkjipU0Cbq8lexf0OCOiz+59FVXN7WHueiBtJUuMB
12N1gl9soVX2wM0GSQ7QB0HrHrHhsO3q66PI64Bn/asL5yBzGKG4jZXivA7YkSXt
r+ciK9akL7kYAIXJHj0SsbKeBw3ElmMDg6f/SUYZuXMDwHeAxUJREc1NgKGaf3uM
pe1BhUMzuyv042LuoG9tIZba0CDbHQ01rv3PUdguWQ7NwkVILXaJ/lYh8+vYa1z1
P0hfRquttga8VTTWxc9B56ilsmKTOMHGsTfMmJx7McRuz1/wSK/44femdm7X9Ywe
6+u1O7O+qEc29YXwAPM356UgG3B0+lBJ3BrkYME+NGUeJOiCTl5/bSN/SEZndxyD
tdFDTyYZzxX1ozk/ys/yve+nXaXulzmHryX+hwzGtVZ2jUk/i8Epxvv65WQstGUB
fftlM9An/keJI1VZ32s3rkmMMe73sBgpNeL22eUkq5Whcg3RcFXzw1AtvtSsLuDV
7alFO6lJB4BCygYtfbz/16rnodT1F8Qg7VU2z55BMN6CvUs+CDKa39QRKwGFncK2
qlx8zITxslzy7jq082UsJo+gVEjd5qM6LB0BEBvR1ob4Opmx0yyxe0nIXmXBa1t8
k8yiQCoY27TLBTAW+wth0IGqgh9hrdVvVxV3SB9YK80xpXt3xZEnbZbxZi6BQDQ5
j56qp2BtYYR+0nPoU30H4Rwu1b7i5U5NT8RGdLlLyvThRvs1E1x+n5OS0D4aSgMA
39BeViWEcD7YxKlhl4GYVPYy50DdbPPmf6SeAoDGbCUN09efKuy53yykmrpyfxR4
ZJLFGBV+XMBJ9NMpzp8kkN2jeS+jLyMSJkaK/JvSNFuhHNApxHB5nL+Hjiq01wNm
5Ub9uPwL6N/xGH8IL4IkCEF9S0A7jy6Oae7ThFo8hVWV4lqRu6guWwYHZIn2W+uR
QPPPnPuVsOA5gYuHcJUpjYNsL5wqnGTN85lmaoozE8EMhtjfxNkKy3afF+tY38fn
hTI6Cp1uJi0UioQWLdRQTHk2nmjxXgmQ37IbdMPJ97dLfBsJIvgvyHMdR/DsQOBG
7j0Rbb6AT1iqikW7cI83o09ua81/u5fSTFlwAUnp54FYUmaxVdMTKFAmQDBCjqse
9UXHbRGRrJPGOVSL10Mnomt8xQo8lRuPzXq16aN60KgXc07o31+ypSgTvfV6fIIF
yf07nBHCzlYv3kXnsK1Yl8QFpE4ePNYr1BsByD5kEgzCs6CNgRmyh2qzMMTxhPbf
soUNLjKtYSgix9misVYwohRpzloMNZGOAtR29IJ7fuR4peYSlg2mf9wF7PB2/oNx
bpQpG0nTN/61ec33aee5UKPIL6LyCJSB4aj9YZgvOEC+mddzVkf92ufWMUuQuxe0
q1EFmUQNGYngd6pGTPfZLT05GH4l8/A2u8U4EzNZ0lHR2wjo5F+8GqttapILdbpU
hm0uUkRONlyZaf5AWVKUDOBH0OYmAy2amWEkaSrGQHAHIuhjsYNgoVdHVaRVH2vh
q7TgathNpaqzySF9Xtf0lF6cha42JOrZ0V2g2b6lLjIn1EVTxOberLjlxrp8bwzB
SsWOtQ8RruLLIZ7GS6wnx7szpQL4NI8hAdZ+zk+dWBIt3X8wqYzDJPLpo46pl24U
/xaCmlsFJEPm3gmwN4hS8EA3LCzlFuT5TFP0sA8eU+MJTrrti0P09dGLq7+9atvo
2xVhn5KdvSgFUkC+/zU36wR4JR9Nl4zy4JUdV0gALDSk1Cyw8wkG0urOqAQT+CeT
efAZcIXK4ekZaW7/dZETzDFsp9382JA1tpULWlDSp4HhmMK4kUXjXc/Y6GHM7+FX
OF/6jwlZr2DgBfz53uT+/q6Yr7WyUSkrgltI1TV2Gj0/WkZpQNiNaaMCDTKB2dnT
jcju/stnRQnCLnMcMjkV0THXCKtqCn/3ZaVbkS/MwzZbLLwFsQZxsNvG8RNlW7Vd
8TBrNRLRPUUGFDX4ZsGWQr6/MQL9cvV4TieM+2DbbKjSsc+bqo4CYbZwi7SYtmSg
RuHUKx1RhZs1bJXa3Mlq6icz0GAjE1XaH/k2Fd6iToprTBeMC1D1Y7QnMbTK6sri
us7+bkhCo5wdJEN+bq2D9vGhjYsYLShcnN1uNy+XLwnISu4+zZREdAIAtc4YLGky
pUKY3ghpqUAshX/tOnnoDwqu2RatsXSCHs1S3cUositkO1leb7n9EA28bN6CdFCv
vVyJq9lmJSDkwMh9RT5DHOhcD2nVOk5xHe/6F1C/cPP1uumU1b9FNmLTGgaucKf3
xoLXTEgLZ0SvMQqgqNpL8c69xaf535zOnptfKfIKSRgiNtLK8SQqquDNmAfXUtEe
CEeW1EhGamtUsyCyW+nEtz34CrSvIYc0braJ6PJyh15Ceg0rI8EKJBRYqaNHKXVQ
WlOma0C7PFOlSyHZuLwjxVySCo1bDdYjkdT2/mPY+30T10v95Xk92K7GC+5OKYOu
98y4eXK3GgCRIBaIkwQckGg/Se4cFlbrgpbQ/dtThdoSUqbrMelyr7w/e8eaFuaG
UMYV0XN8EZNfGqo9QSVVFAoFMYPxWZ0Phixrh5MXP7XRiqLQOzU4v4Y+mzMu6z9w
OU2MwXEtN+M7iZqf4oHSS048PENA7/OEirAKeh/HfWVGtzqDQx1PlRqVVcZCqjne
2cZ3VV1NlCnW9c+5I/hTVPqNb/SuH7Yxx1wp7sLFOW40v0nLUv3F4oHJ/H5umeFd
D/pajLHdGwe9x+SaZZXzy2PgBWNPUgS0EorLPXta0QmAOOLSPF7gm0g0IjBcP2ZQ
xrO0yVviet7QZ8Q3ZJvGgL3y/PLMHQek+DlPAxgK9qNdhohIgLEhjcr6jFFdeDaE
3K76dnnROlg2SYrGQcULL5Wsh8sL2bS9kvYcxde8irMZQyJ28nXAmk3XFm/1l8dE
Va2NTgYH+NLO6lJjift9T4zBR82AO2zbEFmKuQOId0GgAGM03CZyGQ9K8Yq2ekVv
/SkSly5p4s1wZ17bfplIOx/qxxmJQlVKxxcxRHlY28xVX3XtP872t7jjUDO1YRIZ
Bf0BJhOJ08bnM6ucQw81ygO2RsHR9atPY+ZI41rNmaH6R46/bSb0TdhwhpvdQWRy
c4WljkAHo2wh8PEG4KECVnVxWSxN7pVqQP9Apci0Z2btV65RDmhzjy4bpLxUDbtL
CNRhw7EXBK0X/cnZT3MzTz1f6MWZlEgVmtcST3izoRIlEy4MQkqbS2nv89VeDezQ
W5YbW3UZyKlR5bMJ9E88flPbRLV+p9Yo4EFbZooZHypD7MlTVy3QguZQdeNUpOxN
DxJkdJIR0r2+TsU25Rcm6hSs/Ys3qym6MiYJHLJOPUXhQrfNBCN2VIERnNVqCdXb
N5wxAZHqdXN+oURzkti8WVl9YJU6LUb0S3n1wOmH8KdzTZRTvX1YPE1+G3UvWBvE
giGrNwGeGAyf5THrs2uuN53ErTiCED6Ez09pl2a/buLCJMwnpCs7Lw7zqeOgljuS
42T1K2DFxazQhinZ+zkZKmYNTPpin6wpgd6Ik88U/0dZdvl7EAm5oa1iMacSnyKN
k3TqdqoY/fWNqN4ONbRV6/b7let9DALWLoYTMVNSyco4UXuaF+TjAnwK/mWbls2p
XmzalfLDuLwqWCFW8iQFxVJr5b8R6ceLwfGedqVEus/N8fHA46Z59NWPKbIKGbrf
vwHdFH1e6efqsLei/eIsNfVMcYCFJ4EGq4Rg+tsLn7ttgloFbcsL8fLPqC1saxKh
zXW9cFPfRgIws7ufp1aGMHFJspMCG3KYWtBEmkO/oC8nNASIzW3MELUHJ0YvxZE+
TZo5CsfRee78RwFXvpEL0uVPQQ7AWG0tBu/zeKGq8Ow/gBLeFjmWe3S+9s5ihD0Z
dsTD/OFCmBmMkzLBLPXhqD3ZuGg7LVxSTdosUalxos2zLYFmnhkKZNrCa6L0xknD
bcD2PNXjp5N7IKTfPdjf+/ccWuXwBit6OsdJBp6N/6qDUktyrdohVj7ht3OcRXME
b1Ki1KGzOklOxFpDgrYS4tV6ASxzQzuAV39vdXfK47xoUV1q50sym8ufpFqOTBMC
uSlOS630WLTNudlzHabY+H/FancuBCzQAeietYUjgoMvIPVaHsxV/+0wOC5AaLPt
BZw1cagNIFrc1UFPlhw61Pywt9sEKSPKHB5wdR2hAcYjrqkU5WAL6f2MqkmJSWja
5QmhgqnqdKGbzE3HC/lVLFo5DPxJ6iuZg23uU4ApVjKpXO5WpBzs6a6Jk3TAKpKh
nHJswyTDNGrFxDnzWJQCkj4Nt78aFz9IFZzRyyZuW4bHUNFdbFjVyiB20JNhqD+l
VUeAikKITXfdFdpy0WRWGDSsw7HHJDidF/1brKY1lyff9oebeNLS6/YCIqHvyQpH
mXn3TA7T/I9Zh9U1n4STI7u/RUusYxOScGs8/s/dOoaNVZ+MxtXBD1v8xPp3e/lY
ypoD/o5zlUEtTd+rbyuLGBVrT1hYRWdjrWxPy6qc222K31qe/Kob0H1c/JaTxXeg
+DD/L20rNy3ZvRog9woHskXhiHUVBd6Q9IjZXD4ExskrmsmHxcdkhUE1hlpKOA2O
5FBBEqF9uxQoD9fZFbGlQB67nmgkewbD4r7EIPkYNMPQJN3GmpBATnn4fQlajBwp
yLK1klnKcIZfwzthB2muOa1P/K8Q9EMIFjB6MzyN1yuUPnFnZN5f7MWG4DklYRLS
ObGQXgPT2zjW6aXZk06qm4AFNhnF2yVLGpEBTQe+hUbIm0iIMtIE9x8fje+JA/AS
khrvkjA4mxZ8upQl8R+1+3l6jw7KqDmwt/R712eiGuBgLEA0YuFG78jzQk7APu5O
9AzA9g1HT77D5C69OP6IrCXpbMfWTYtli58WYITIt3CBt8cOPQaXAU8FK2xZVRFm
+yZ/mWJQQ1e5BRdCUV+D8KWUIibQsznorI1puOoouA8x9buqcsGfPgvj18UN5PfF
Zt1N1P4obgDu4/yazxpvUfjDN+VaPIFV0yPvIFNNVrG/pPZqAqxeEIrWAeZv88tC
3Jc6GVbdyx5X1g6MyrwBHXKYAInKWH07QuS+cqQFkkQuarEcp0yhGsooPsXzSQzK
HTYx9BQx4uIWXfxfaIqKwOq8xKjPY6NzLRbAb/ZxciZ52XA/gi371uchUAwGIUir
K4519N2JmfbtrkVFgWAZlE8A2mF8djYuRS2lBGLuLpHL5no+88fXVnMD/lyLznCN
Vk0JYTuL50SZQohBYDzpsoDzi5KYdlYMkjbWTVdNQNTq1865hJlvihQJRoX62NOC
foR2+uoBBMbE8MsiCa+VwZNORe/0+E91h817mQ2FdYPF5esBkdouh8zTxwN36eP4
TJWL5LB2pd9uK1oLyz0o05kCqAVQmzUyhr7W3IMp1rxyNTPTemFNq6j4QPhVcHfJ
qWywjYMfd/OpeOVbW2SyIuUByMA0fBu27olEeagzS/pv8h4lzoynAaAWKX/iwQ8t
v+gxnz1ZhPup+ZK3z4FcpeKWWzYyltCweOJX8j5+C9YfzVGRPfBeBaSU6HfKZOo4
zdCuAC+eRMlb8HNeW0I3QGKpiiwwOp32+dIBIhuPHIkY45PLN3z8vgnvkjXm2zCh
NJgP3clA9E0/sb3oUILedUn8mcSQ3BiDXJFL2JMGxXJwSn/JAP/JZN1P//yiyrtP
wBTDSuvC3TS7a5OW196BECrRJXZy+qtC0Yhzd16UZqm9Z9LWgCuVyPjA8C8/ySsD
5bJ7KQElXT1mbHBHs40gl056SQKDZbOA6jWljDjjTgxhre8cLUDCBDolmTK49Ecq
gkSbgQXo6dLQrLCd+7zCdUZQtuowgVP1wQ1rgbX8c//xVVrYajkpFHDtzUESjpT+
lbVmBfLcp5f9lN1/GEWrM5gnQsKmKG10Q31cteJmeuwZl2cezS5HlFgi6T9lQoqw
5m/gTQaThVJxt3ycjt26pW0nSWUiuOUHGZ9rxbLenLcHuK2BliRxuKzt579hlJj2
8XVEAGSv2KH38ytWY93oNWPABZh+/aJeK2zhLZPxGFhDea5ImI85uwSXK7NtRxLE
7cDlwps0/XIv74VC64MYgmy4zAp0S1OmW7kRNx8axpAU9cf2RWp4qMDtHK9CM+ax
FfLCBEVGqXr2fKbV23ivxoGYmkx+QTrTIjJhltJijEWOARh5T7embudYwetxlMNj
MfAIkvxwi1g1gWBFonShKa6Um7Ia/x2F9OwagjzX2m1ROmax9q6i4xRYrH/4Uigw
TlkHTF1SwyDjFZS5Rxqtv8ny68+CDKv7IXUi880jPfaZbC4SkWLVTplKKX56wX5y
HVZP7a4ud4WttsZnqtEX3wH9A369T1Z85jyr/wxNEpC8rtAsFFbzeHflo4aLnGiW
3Lw4XmtIdGyhk4TPaPFGuCc80hl8/PHlmzkCJ/h90K4En3EwmUFFZ0Al8dUYWBha
m5MK77jTAXwOg2oB+8cJU6Uh/CADG7vUJmxkrsAfEdjJc+1eM3T1J2LLGtJIHnTP
Ruk95m0z9HpNvGoBMw6MLKNWFF9tAh8WRsg7AF5HDvhFHepHZ3A8DURn5Ujf859P
tcEnMwkACJnihzhGlgc7VXcQBTZqbOToq1C4vtUILppdVqHGs4QjY3k8oe2bjQee
eUPX9k65PHzM3x+bVUgvIygJNWAyumcwl/bkSCF98eGePN2+0N9jSz44qpSZAi22
z7Ca9yPjrO80A+InRdBb8iF+zwpDR00lt6q3/CO7mshewyfq+6L78UAQ//E1Rcn6
KjJUpY6t+rWeIPhGU9oH06r4wpOHeUiXLLtRORIQoHWySi8l3XHtI63OyXSrSMBK
XWiNpQix2itre9jzJQgjHhkzHDZ+izrCp+G1O4c9bbmgjlsUUIgGXYw6pt7/C+Ud
z95MWtCUUY0I7JI7wlTC42Na7lzMgmeKR3MFmwbdV1VyCN+pR8jfFCoc336z5u5R
gL0BFsEs7mL7Kq7v3uSpmWIPb8qjW7S1gNt9o0fO19rE3y1IUy2SCfXeVBC7RQfM
3tcZxXE6MaIKCi0+Dq+dhuVcyOhPHj0Ghw/FSPE67d4LeWSPbu3XQcjQIr/eujf9
DcS8fNzRBimsIgC+z3PEQO4XQk+CIjg6uzzarpRVcxLy+iCPr7ThRu/ebQdF1rHj
SnthyapZuszbzb/CIlET0PIuxJiRSnlh093u16hwdWNNovnA7/+B0Ijk1JHnO32a
a81d7QTmeV5z/UwZOxQm9/N5EXGNKJqqRrLklEcay13ylLd1CiCrYjtHDHX5zePT
XqXD+6HrEZIc/RtXEXMC+e6uxDdKJDAg9jdOo0qT/nGXc0gkG4PEZ0bAmmOnEeQ6
Z2hwv+Qt5W1POkNhvIu9ITMvktNOpCwSyNZdOIyTP6geaf9ApqRwusnwrNgC1CSe
FK0h+l7I62AYUr5gejOwxVzxRG8Cdn3pi2R0uhSU4YeVUmlCa4r2xUJmtwHcGFQF
0EBgPQnnAEyBkh9OFagf5f6R6xIkJMO7FlEZxpPfXmVl+snA+ksKlzNpwh6mtssE
lgv3xDyzXGGJFE0pt/7bgSazj6GaMA9PR6vNAYxkqRCl8Md/uV446LTYm22gMVC5
jKP2c9num9dIy3dj4TMoJd/J21PmdDo8oKsg+NhA/M7IUNhMhFkraGBqvOXEMxlZ
Ew+azD7VhCHO4Y80cMRczR+fJ08ZxEVWmcpG9f1ZMH6GRKAM/ls3IiP4//ByWwnf
aZn02wMpKu1hNv0BinfV6pC1Oa6obqFoVxGoN8mEsErvlT96esGahq2keMnSfKmv
I0IBWsTonUGq+Kvnr3411LT4+XPmMIqL29dRZ1PImsGEEF9eqs29RWn6vvu2tUwy
oMs3O26O2Q/RSuzLq0Oe4bzNkX19b7P0csdyfTWpHhMOu9SzsPZa/qnfEFbrjDqC
awdMRWoEzM7FdCrCQZWLv4hQ0aMB8TQw+Jd6daBj3HupO/vY5ttmyCsED2Pa6oBc
CxMBeZdg6Vnatof7OcjRZbk2F2eGiaotXhrgRP7RCV6HpKPNK68V2pGPQUySEhxU
4H68gsqRglHh/iGlM81mBTREZ/tf2CTo2SdvQbu89NC4/5TbXB07T0A1V1Dbrwer
gEcx+f1YmIsu7bXHwBe8GZaVvwPb+WZH0HIsdI5CS8R0a1jUojy9M+1sF3wK2rJ8
DcUPi7eITB6QGU4s5WPdkgZhTZbA4bqHP1uBMTVCBVORYkin34Z0EnYy6h/GeplO
5xEwT0M00ST5rwEDeL8jZ5cngjLPkcuYZmqJhGK1X+hROOiB3uHInPUjkJ69SUIu
84gbvSdvz9BZA3WIB+u+H9C3nHGkHYxN/kprU/1QrP2OFKN+77cm3gEp95e5I4xf
uUAiVVJlRNi8wICbpBPZWQSpEnyS/ILjyVh6SaY+bVo8GmbS9z8iFEW2dDN44Q/7
sUcsp6DJvOWs0i2y0vozcDCzsln9rPA0Q1oMIeDAbCcf4Z1dBqI+2Fn0RP+qIpBM
THL3pmpJN8jP/WeDVrwq9W4aDPenQjCYmmMegnZwURhb9VWE48FlHo//Wc3F/6GH
Z7v92blIPmWw6L4TYMKNtjdB7ehwkNIR56h1OR2Q3hUJTFWYiWUpxZ2iGRbQVooz
gXcA+mVB5k26rw65lWik4Q98mEUC1xZ6bXwuTNDXV4Qia5YhHzuuirMqYsYseoNL
LdgtRZTwI4UWoCFg3HspHLBxDzIbuM0ATl+XvcIUz1kjBC+r0Wl3RJ8SnDDt5pvK
h1qGKH45CmJSKuIXUqNNHCIQXDOeEGyjL0loZdg31Ej42cqh0u7K3IrLO5xqRwML
sRYu1xOFmXlrt0r3zY80zPdYhlQ8Wi0wINd9cNh3+Do1c/221HYxC8Vh51vXSshP
nKP76U1Sk/fGrxFhKcQDMhIMqMXNw3f2V0nlof4h9bEsZS03lGQir4BjCRTVy5Sq
wpmhcCfNlYNRiTvXAtgZadOV63KAo1bA2zYJMZlb66BvtgtU7oo5airpIf74b71H
e0JCPtkSJ/moK7OulP2jeeeR7D+4JyB2LsjBaW+thQgaDBezwo0+SvzGQIPQpsVK
0dLjON+ZPFSR3Z2Wn5GAYvcuKFJrZlrhXN/2xfSM/OpW5PoznNX9DVfESSBr/gQu
M174gOkYKzx+avfKzd0k4TzFNHyN3dCR3kVe2LuLmYVQT9CU4ZC3bWqwePMV0GTL
y5NuO4xdX5aHIEwcg+sS9shFW1pGr2XDmYmPfm8t+f8ncoCMO9MerCxKEN/7a5d/
siTbSt1qzteGJ0C4CjjMOErwh/y/3aXyuoZP6e2NUUjvHRPSbOXJZFlomFYbr+Ze
522YW9h2MEk51IPTxKbBDWsngZbEUJFJ79e3t4Bja1TU/htzvs5ttMn6fovQCs9G
`protect END_PROTECTED
