`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/pflemyhA2Wm3Nkth6DGkAn6GBlTt9N4Ip68M2xLQp6U+NXTBEjKei66jji7NbU
WQ1ksJiSTd3m0DAbKNWt7Y//+eA96YBdzscX21ySelic/o1aD6BEEVWkmEQUiKlQ
rXhYlF/kHsUh1wchpYI/fDLq1ymoVsjSCQgCy14RFD70Z8/CJJe0DzqOj3p3C5fD
PqSamgXJeljzWIKsB/vIyMu4CXud+YLtranx9KZuuw9g218BoyxrF167kZ0CVgat
xr70IttfZLbf7fHS82l8SetINsTxWM16GwepXqFEcjl6uAanyZYN9fjr/MP9FR31
mt4DOP4CXIZZjy8QqLg8VUD57p1w7upT1RazBNmUUaD/cwJh9vON6BoHaNcRrytx
e6pXAvO8XpK8mDeXcZpbDx4tXBIar/DqfOi2IHysz8vnw0g7qwLi5YpQVJX3+LHc
j7gXNcQMnE7G/2sqYycd5Gmf9ExDe+EFoP/YDdFWRCc=
`protect END_PROTECTED
