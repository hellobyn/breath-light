`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NapaMOeHWRtGx+yGH4jg2S9y49FrjUsvrGZ6nu63XaZCFLXEBQEnv1E9rmqMHpiZ
ssUvNmof7pNxXErQ3mS7PwbSRlDMFExwIYWA+kROogmClqO0mNaKITsCB4QRUEXi
KYMW1aKvg3+Yr+SoEWB2VrKhIbTQcp5pvqwHiX2TIH+j7JDZ5pbeL/ZlP7kY6IKK
WkBdjyjaouEGoL592YoxN1A7P5puyr6/jC2i4llOuKc88U23f0Ar3uWIkPOG3uGe
aVfM4jOFaO3tn1ddPM0TuZqLyEs069gwbt/RQYEfYjaJCdX6zp5twRfq9qpT/BJz
Yao4qxNpFhcjWD5Q7p9jdB9a6U+T6sh9nXY+5K7ddjGKvxZ/U3QCYyxJH81Fw1v6
mS58I/VZG65vkKi6zGtapFVgUkIXi4P2fOB/vKz6OYE38vnVEo6qs5tAyUV5q0wf
ynjESGwNVEe0vJzFTIa5nqYuaHPhNXrLnRv/1sSLiN3pyGYlfU/dGZ1o2Ob5IPwL
Q3hEsU2GskwhlVBRh+Y7qEx9fp9gdrfo5OMlJWLa43UxnGq1HE11My81DGEnawCh
aPE7Y4Q/subH2FxwYnKQLHWgSIPMbQbMd8ecsLLoXVlqR7yjuT0KCZtP6W3p0GPb
gimDcaLv2cv4rltJdtBsvoB8kKbAw8023R2q1lBiQLTzZtiRTAAt+JnIK+ww+pvm
WpWbkdO+fjI5Ba2zXDjD/TQSYU6fp/zj5E8ruXwbeJJE9UbUvUHo2H+gz4n9ZKhk
NQL3YD/1qj/up67GPdkIcJiheq+zZDizecXKYyONtj8SWQTkZHqJTEvL0mNAEr3Y
qUdKs4RkgE0GlreAfVtKu529q4S6j7tXeRDGM7VQ+y7Y2HQhjfSr0fdru71q0d1H
7rZGKjY415f2e/BAZcY5C46XZCWKmN+KelkoSGfz035xLQg2EjL3L9nAvBhkevEj
VEqeVajBhlXizBig38V7aftwFqRcxtIwgdMJZXA/Rpbq7uvebFQJ6nCOqi0UfLPZ
oSztKP1+7CmGFemyzrOLENVUKr04EZVq66XTEQaUe6KcHAJrLh889D2QHJ/gruRQ
GkCcUIWtUIlJNQvXOferb5q7TK9AY1SdHv7FumsRm4Kge/eI0F3JQYGV8Ei41JP9
snwxwdw8+E8TCea9s/LafK+l8v9BfeqzRC+qwSstIJMunn9kvJkfy7ZuWRK2JbSg
DSivYvNtQ1VmtMzMTREb1DYoajS9AqrBjt9FHmPmEmk9iFQ0tZVi73D771UFKax5
6lB51zdWNWuWUYAsr5BNEk/R5x5QodcidIipYIXkUd6XUs4LWyOcgoObj13Jmhnr
jT9YHt1Bnc6oz4HvFAC8p+pHvMKic1GBWj+xF7wBZ655xqA4bsnjbAGMA4a7lx//
NQ6LMvGdtmUSaA/YQNQJ50D3wRH/Wa+QoAAiK6YFsWuK1YRElPen+sfuSysTdESX
Nm21hPuq6dhXxD6xCFd4qn0q1YhUeZqhPjuKg9Sy8U8HN5yTne7BcfCNihVKbomc
apHmFeDvNNB4XeFB7s3KGT1jgjEZa77uJHklqE+R1WSKoulla8yiblbKyPNO18Gs
Q9eqoXyBZspsQtyWf01xHzX+dr/BRTahGAqmSTvXts6myQ4CiYpPrs5tSlxPsAl3
O+QGAbEYzPXnVU+Ix6Ff/fmp4XfswbDkWrX9pEfl5OhTu5T9GOlv6JTA7bh3M9RS
g3iqXhGPIxDrZbcSvD0t3moUu3Ib46cp71OQnfi/e4iVEHTSUaWO7LSsNXfoKq+p
f3czZqKhOHU54uKky0e4F75ye8uUdcSCbcCn75HTNUWVeolpmsnxRyPqubXK35zE
Tp6T6Ev/YMP5wm0aCgiLtXXZWjxB1pogOhmDBUYf7ZMtH9LZTDMlJmxP8bENAwWf
jlG2EWBozzKKd4a1yBz8bUzGJmF2TM52CsnfBUKKTUFt8T3hAbwrtHUSOUZ6f/Y0
c2PYMinFDd8Ol06301EAfjZErCRTXsovO2fCvR2ildZefEvRYSt470J7fNS6YUXc
AEm8Vyi0GS7BVK5+rprML1VRsw2/oWFWhSpvJDwHhR43YzfF0fUqCHt+mtcm/HoH
tyIB8UmwVLLyT7Jyhu2p8Or6lrpapqspvLBVDdro5zZJbY50quovoR/yJyF8vQtT
Tqc6IBmQXuIyip4EfgjGPb9UseypN1UEkizzkSbwqdJ5grTclIgUkk0w/q9QQJ84
nt8cThPfFBMJjG93FBggLVqLmpQ2hEHVHtK/8+3UCA5pmOzr8ppn1Y7nJxr08YXF
gFKqwKbWgGc+XT8qqaunn7Vx/4EN1w5n9zEpPDs7v2scU1itgTWHCqmyTu0wWtBF
g+aujikEm0iIrTphDxXXtoETUWuLJC8ZSJxU7QurXMrdOeTmC96Ppj7mMtBFJGxH
YUolQMNIsXS9fhfcpO/BcysNgESOzV1Fnch3RzrNMpXySn0WDtCLT2dmlLCtyF8h
zSw3S6iWyq7xeWklXg11xA==
`protect END_PROTECTED
