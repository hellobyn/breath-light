`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vf4xFstD/6+qgaBFFOyEMrr+hLgu1oJzjg5IBxQ1A9KGiz9ePFUyI5Sfd+QPCi9k
94Iitz2JL4tzaD87S/hP8RzCAVtX6/PpjX+Rv89Ol3q9SNbURNF0732q8khatSYJ
Mal6lDL0+FxfVPmAv1skU9ylfBG5EKgCv+jqLEnXPbu2seAkoxopfFstdKjIKdQ9
UYsvOYglKjxWDpwlCRP/IHfTzfwTyy/+KwuOpcc8w/P2OljykMzvoHF5lLmcIYYD
2aC/W7PlZ8H2F9WU+L+UsiinNYSut/+Z9cmTRlzzJac/EW4oib0wkDqNq+bA8xV5
4U6QW+WNrVBU7Ud+gObC30QX0KJoK27l7xZy3SJ/Y3onvsLVhr2ei2bw9W3vZIGd
VlHakmQ6Z7Il3/17UAy2od4HIMhkBH69Wb1tvrS/WBhKbaxR1dTbQmnxetQ2L+q6
NtZaWbqWRFJ/ik0Yk/4fzwEzc0O4HaOsdP4NmysgS0RbZA9JZ1X5iIvATdrW0wMH
vN1XjBwVW6agjFLxqOrCMFYsLpQBCwSfv2iRD781v3zMNOhEr8bCiHEfBm6Kyqcw
`protect END_PROTECTED
