`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YESmegaXTjr1VtdVCduxDHJMDi9sdZim6Au+r63kadhvaB1Jj7A0Ap56g3qGU6Ql
AoTPPJk7cqOFXALOewG/WCBclb7B7Ew8wvI2FOa9dW5+kC2BPgY97X7Bp0tCyCjc
kAr1fsI4YsVKGNQHtl3sFjxjoLFK1Bsx6Wy7noo/WzB5nF9GAhPWWN9W5sQtTMg7
USyclDTBZKNB8pmNCXtNQRIK+tme+4kQb75egbXtTu7GmbYPv5qTaVss2TUIHHFu
aysGD/yRJ+iiPDYD81ZXLKoQCowvgRpJKKHZsWrbMsa/vB88lI9Do0oPoNDlTGvd
j/ILDZJPXptzSLr6cpTdeg8MSjQx74+eQBRtNz/Fh3CLJl2IdPg8jJq1VVhJqBn6
86hgrekbx4pFNjZO8R05uBQ64ekZ8HaW/ANJMrpOUQjCUqN/p5fmHxxAMfGzqG35
ICBxpIJsW5ysQyI4F2Gx2pVzyxQP9+9b5WacUbGupGQ22dPDmRPY3DR2NNN//qAV
CnbI350e5uKmmhsQWv+dCIHuV2t/ZEu9+JS78QFSj990jkgIAFMw69H+Wz8h4UyM
hU/b5eaWv39yWgMre92w5nprvwbup6utfjhCd1XnEdvxvpuux2osrbYv9Rz/r4G5
XBWxQDOdL9F8sp/kOnl7RENqRhAGmjh3KWauzi5hAAUHLw8Tb9Ig4o0vOulQdGQb
XhtzsrcWltxRGeK43iFjpOhx5a0rbKNocUD36zXU37jd7VEUvBO123+bahRMoeHB
v8u43oY8344dZlFxx/ZTMINE4U0kvahw2OcAA4Y6TcLr+DWia7LmIpEQNJxrXAC+
JZCk9aEmBMA1OdzbuWKcLiCzFYjUwhraLGDAhlkL/TV7GKt/QuMGQ+Pbzh21iTVG
QiHa6t3xoq8AtDuTqGRho4Jy1Tx0TSCIp5xjlcwANNGiW6Vra75NBATWmpGFGGzD
4oNNktv3PDOOydx7gjrH9eFv2Xl6mIHUqYnlHcdJui8f0mE5VAQnaCRoBAbWIuzf
ZiEqghJROJPeDSmOQsjyvUdfxD5JbG4bheLXBKl6aLakhoOfNA/8Mf2qFCqR/nEm
i0bOmgv+fj8+KyMygMIW7vkG9db+LcflB1/db1QGLjdzfJMQ19Gu0k+BfrmhlyVh
9DDdK5YifwYRdpnkXn9XTFhEe22rw/r/N6QGdL3kkKln3Xo0WsoF4Uf260vMC6fJ
UXaRFOBNeBhIP8WgC0qA+Otbv38fOGRqtwKIoVZukMzTh18v3417LdqBbsQG6Dns
8q+YOwqQfc5vzAaS0EPPMribBIBiaSaMSKkOZ77V1H7NcYGVgmH4OQEgODrXyCZa
pX60epB3zVEamLtv6d1DmKeDiaX+566dOt48kAzXPHc5fiPiZdiH71fDlxxHAFVU
retB3V+LpKaFB1OPVTgLu/mfUT8M0+6UVvLmxDA9AaeqvQJ4SLNMTHmwe4pAvdiB
YfejYqE97RJwJQi+TFu4j2TYy4ZjsQok2z+MJ4ReB4vOEa1J+yaQYjw+a611wFQe
/4aGoqbIJqCNDxarDKhiPXHK0fCE5oVkz7T6Mh2KAdCyP4E292lioNdnBznVHNSO
85nyxQvdkFVrCOuTOFogSaDXFIQDI/7buFvsIiv8kQk87QO1vlMYPFMuBP/7D8M+
OeHQwjrbo8VvbMpl6++sbtl9PIPkXpb8i3PON7NAD2gk3utqiXr8DtY8pxb13V+T
1FvwSxDbq1l+dS/igrDgRYlQFrLE2dzDXDCM5ukqNElBNc1hamirGyKN7f54r+Kb
+3otwAw3z/RtxKmUflUh8bPQEjiScBrx6ms5sDGlV4a4SaRBV5IHDf6w19AQrQlY
FQMrxtzvyd7Hu2v+v1gdRSbmVFyJ49bs+dfHDODPDqAhkMZx5tPuJsyD23GbY6aW
rCpbA2AGSOgAgsU53bQ+PVaeGWhKTjwv0mwE50X85Fx+jJ6h4nWRsFQm9qA653xo
I7NwaoTnPbMQHK0sTQoL8PpHwI8Y3XcsFEuvWuira53YULCmFiVoPRsDOHG+xuDt
v6cdlPtU25Pok+aukMXy/HkuhCCtDJEZFik0PCPzQnTqMt0t6/rtkF3i9qlZ3LSt
+Rtry4Ld0Xdc65/n8yQGfsdQZCZ8Hg9BLRoMZHCIUi2yifHn83IfxsGm0ZWiPR75
iQ2yQ1eNq57taTruJtDhs6K/swI5QBrmyU9knbQUcWNU0pXPlA6CHaaP43iOPoJ8
XJDepj2z4ATReQfMNBTUPIoi+Asj5hV9oINLdkPAMBi3HGqInwN9+WxrNyRx/8Le
wsQbln5uV4xcTAXMFbVMS3hnjQEbuA5mNODSFBv3WGIxjg3O6yVunbnoG3sVYOIW
vTit0iuhmQKaUVQlgjH849mdPkkoTTGxYzG6JOBosf8bFm1rv5GAlKBvvSUUjwJI
oV2IoILkMkmgY5h/jxtj3D6Adu9poZiMQGiRw7W8Idv5hfV/bQVagFErs7/C7OWL
2VPPIUiGDhIp6CkO5YbatP0Vntax2T8CQKTMOnrNr729ah/fN3qtldABLRMVH2MS
gqxd/nBpVVwMSbrmWcl8g321XX6gb0RFbou0zC6mUwQhpWrbaeXd90gljQdhB867
oxnMtE7E/86oqy6MISsZJMCx7PBM7RM/yfXHJYoo5sv8nbRF7HCEWh8EnSqvZuwr
8BNTi3rly/Lwz1My8lKSZmB5RRwzHKvSynVGIO8JdS1CImL8GajksfUMTmCXWuJ1
o7YlIDTCg+CVvCvNGKy8Je8xliUfCTU9AUx1+STS4jDDoaeKEgj7MVKkuNf++Za5
L/pK5BYXi7bd8rq9uxjoMHBNAkfnrhHdtl9JUuVEZx+JHzehNBVCbhDdtCPg9wAk
86Cfq2vc+G4Fyr5yKUQnYSe2a6FBv46cvnEnZc6LtXYBUjzkVFwi61Xn2Z2+Qi3Y
WDm0tPM6cYowd5DzmzQYbxWSxleItWjCe1Xs+3j/IkBjaAB6wZQ39D70H4VG12s9
oDEdgL0j/BIE9SpZsWBBi1ag+LYadgoieXA0UICosYHjERkdQF061H4Sx9ZPuesw
qEgjoc2mAAUzthTB9+1M1KdumLFkymOAvwNO27z4xGttRa+W3j8qpFHT3IHCMMOG
dhsad7uNCkgzzHprh5KhSceSquXR1gdC4DiYxd81f4H9I7oAmHXyVilrg+J056de
tJ1Xe+1UsXw9CUfMxV2Cm5q2kPMmE3XSJWEFvMjl1Bnf8OD1nEeXX25bmVWV6bHB
s+T5Qtgoj0zANc+s4I6m6sOlsSnt18vpepAoqJRu8sbnMaEnD2/7uD7F9mCrJPTL
uOXdulafjTXDr++yJ3anPGYqAk0HFopUa09o7pzksN1HX62emzneR6KXn0PcSjed
e0+itvn5INu6Dm85tjikyjBfG7cBbC/fU0xYaRiRE3PotfW/S2uPvipla9yJoH4m
3+sYESe4PTKZkH5OQ/T4U8aaqEU7Sl+AOsNy0bZMkN3zoj4lwZornFZqfez2iZHj
XxunW+AP1tDZXXF5CllenQNQOgVqy4EKwc92sV4zQxPTKNnFygeFWBYkiHTh1c/P
ZxKu3ZaSEOI5W90JKi6xUeJfVjqC7jytGIgAW+U1hXgHr7OANKDKQkZ2cTk/QNyo
HGAZbECP9YUXJ5EoUIv4zsAgUFroFbjyoPgNK4eiKpn0IveletAERkn+Eb6kOzSD
4MmH+br0MwJmvtsnw6rRAwtV/2MZ/3bwVNg6squW0jYVesYQ13EuxhXVtS0M46rj
78OU83Nz1i9XScSveN6M7BIjsD94++oGdr4RmgQKuBbD+NIcMXbTgCg66hnhJtJO
qgYhBiY4nyw7ElGqjLtVTLbbsFD/tWOfwxAfQgvV64h+7K/IXObmIrJBSflHDu68
bN55G6STm6jExSLl+TbXrlPo6arirulfna0sB/Lj3QipY3b1NFS76mtaXCqTxLop
ctjSNRMMCABnTeO6Fw8FpnUi4EVsN9OJZCXSjg1GY26V52sIfjt1oC92MhmSAOQR
MiqtnteuaFLp3TCp0cVNdbaRX0WJ+fJDkrD0PQdY6Aa6vNRV++1t+wcYze0No/KO
1VfJ3H0W1MhDL6/ZP4sn4wGUKm5zoBWnXJDETrC/OE6MAFL7lOhkTgkCF8UxYoFp
wTIie10AIiX59BbJ1DJGVo2mVrhqllNbwzOkrn+rYVErZW3EPvgTVs8zKFc+P646
44ftl5Asyk2cBj4bt6sK3ZbC1Pc8TUrXTA5cLMENYq70IsP2cpjdw812pooHYE3Q
lRBO3/CVR3VgQek+oVrqA9PNq387uXIskmXl97ltleQYJpf7mT25Rq2DsqkR19qe
0szvt40EY8MTVNWixItC4oTqHnht0J12zv6V4EyorZKsJNVf43SsiIPREt4O6khq
aBMh9DYXMCnt8u3n7i8ydFq/hEbEkjIfyd6KKL0Zgla8nSHU3FT89qPJBneaVBb3
9AzapKPniu5Zubl6ManueemAauFXIChgAmB5U6iX27hTnIYAqJQed2BtK6oHVXWs
qGKMTgbBLD0nZ0RqdiPEHpSdT4U2GHQhhBkgPQcy/VZXgdqFoUugzo0MUXpT4wav
1Dj80epkRNQvNactmoVKaLOt/CkFxvRELUnnaomSRIdP7lyO37+wBJ0hKO+gV6ox
4EI7DoyFWsOBUruCxXKcH0kRpVEwIEHeVj7kSVoa3JLrsWoW+bJZB3lpo6nHCDOk
vBgfghw/jbS5FSoRUcraq0RJO3GfdoD2rDx00GZvO6gLI+TjT/Ou8nGI/yUXKG63
uQSEORraCx3oGYU0tarN7CLe7hziULMxWoGwkrfa6rAzqL8uwNc0Qj08dNST5iir
OBJEUHYnWhIup7IkjFiYMDCn9f1yVnkaCTrVXb7qcXHidPKPrqV4Ynt2FOfC6Hg5
TN1FmAlhF2qgLY7QXFQYRf/cQ2yb9Ay7h0G5+qhVHxvV3SDjJ01QYoheXa4ojGTp
p2fMO+ImDyGq7eCrT9uFXlVtq0oy/CcP3fFHqjiEgw488u4FDjCoxaBMQ7rvDk9O
`protect END_PROTECTED
