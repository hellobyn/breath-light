`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLwfUPVVVayqZD1mzAlT8/byL3TcMccqpZOcAJ4gogSdOhA7b5MuaLIB01BkpGGR
IcptDWoHfppnYdIZkN4HZtdqTzqpWwX71w8Kp1+OvSjhH74N7klyWXEPjf7OdoEO
A5aebhGiyEdBMtJ9FTIb9yd/WcdeW0/auOE+kvyLhL9132LbbGMEGOghCYhp5guj
jxkVzhev2jy5AntN/4lRXWQp2qtxbRYpuPTk3AzJu8bbQwTJvuZYudCoYU7RXg9A
ZO41ThGYbiIXKat9Y32J9NE5baw0Ce37bu5rpPEMiarvcMQGiOg9G2Ct178vn+Aj
rtotLFCkiQvbzCql+/MESgPwIbyegjtd4O8Qteo+nERLipvKzWaQMcXzKzTi7jYV
KQJDSdz7bvOgK5M/y+7270l7S+C2bxFmhT7GvBwnz6IjzG1G8sIvQEl/Z4+rbA44
tgvH8blbfD4ywJRSHn+aXwdRRA4++OQI7aAxQWIwEc3iL5o+LDuQ5Uf25XZlDFK7
3V7Zk6X7SQi8rIcGwtcHO07nZc0llH9jmYW3B0AvzajlXIObpSOQArSlMZQE7yim
WOonZNxyWLvLsYbbnYJxxgTNJ0x+3PSTcjq1JBgEG8E6QwoUAKMJJ6Bfs71FpNvV
FmSklRiYSRRK7GBkkH6kCD5HKrsg9zq0aC3SrCVL5b4pkw9+Zj07TChiM6HgQrHX
i+ExdXwa0llISshw0MS7kdKB72OykiZqni3WFc9K4tUxF0b8iSJg4Ew5yZNILr/p
4+nMNEB2e4myS6aYb6pZUyfhQrW2WsfDeZmNnWR6TXHI9ib8prsADbpiSoNFnVlc
2r22MPyG1Arh930XW9F7RNl+tMm5Zspv6U4kEyWHnTiiCFQWbK8NaE421raLx7Ss
OUe3yNRyORdiW7n4Z6cr0Q/ANE96W2ySpx6wCwV3qPXesmM0KWSU92PatAAeg6yB
k4CyCy21Zc1Kk6JfcwVjoZ+j9XmaSI30E8gyXzPPcBta8UCfDqcBttQBVPut3DY5
GoSJvkwELYNNrPx/OJBb+O3VLqkppvP2J0IK6Zs8MlsJqCbymNJ3FIv2e8aTA26h
2EJ1ukB8JerVfGzuNMUXpt9nCb51MeEMATraWmymr+C0GQXGQ9IX4GfDovXz6FC3
Df265TJSHsNmhOGrxxOOM5E9U3UgJlBUKnI7iXMynJaIKWWmPv1UAYvT8fwDdMqd
SOBGa/6jMR0RsyLfZkR7xlzQpjgjNiIbYrBb8SJILTXMZFNBahdEh2SHPYdSSsSQ
fGJhBR6W9t7rWlxaz9j9/DTkZ5mmvhSsLLgwlUoJSjjpen0cEAhCvqC39Xr4VyEe
yBGegShDSv7swk4pmzsTTxUwYpiZs/HUdvLPaJY/2HceLBbNx4EVkczSrWCYMh6w
EoMLSUJVWPIUBLT83ZrmWbgJ5Toiu9wq6GNPbGprGJuioQuLlcTCcsK/DUm5BMQo
A+G7DryXGkTAi9GieXYDYDaPfLpmOvHEyItkzS0SvKJe9tXZHRMS7iGjdXPxvG2H
lhclrxaEgQZSJbnLIbaxg16n/wT5gv2WFyaJ/1DojyDmKIZ3udE/OhuQGqwoauRk
3cbSyzy416jyJ+2mcL/eZ1E6xYIBqv18sz+gXu9Hzhgo53WV4hTq9WmGOvHHvA6l
p035BkKd2SS4TqOoLQT3eXD7gMuTYEiU/t0EXqAczHDRazyrxlfeIYD2uSA4ril5
ldTdykS9QIuUUyaiKmC3FkxRVCqdSkBZFicf6fvvCd5L64a7NOz27PqEG5hWJ+mC
URVKnfwLzEcVoF/6/zM/8vwmeTzK97ZAInTALoSDBrQrHN7JhlV4wqHFiRP8eivk
QCAngnRf1tmtVdqpyf43b+frm7gyo9ngPnL6AXnJud4LsaB+YtwMfaRShx11f5CA
DgE/oeNmCtfajmMEUut7KpGXFVKY/f0dfa4kGVkJGKXqGmY9mNRiY5ULTDr4FwBP
qCH3BUCvuXSXbbd90Me2cCz+JlZ+elEpeG1eaquKaw4QHIZe7ySIL5HjchlbBpMc
12W5q+c26qTLOZzENOPCZfz35QupDajXkPDLEkdOuAjZFmhC2jgc39oveBuPcsRS
AWxtIsCocd1hGvZ4fQbbgKZrUoViL8R7jXuF9fr05PE9enE4KLL4jfSVxB1B87B3
n8k1XmoZGDota0zzKETzKCNOHi3dXjtdlXpxMUPxBe6F2wEbITkhOHCzYz9jyuge
PWxCndbu3w6TteiC8utcC4fQW0u5095MB9E88i6xpdphlGXNX2aZqDi2lBgj6cZp
CtPu+r+Hev0X7wz7DLx2Bp8jVleokHaZww6DJUq3K7flOXs08XGNnONui+ThRezR
aJsXjrqRSMbrWgLBVH10lHGc3tc0blJRkx+cALYPBOKFVzBtvzYU/JWHpt05g7j3
j8cKDBdco6SiCiK9kYuGjYQvkGmhXkwI7HTS6DVWDWqBIxjfIH3GB/SfxHUtntyn
dLdv1eHWa4ekX8IM9r93QMvWoJ4KQClQnUhZMHGoSiG9Ww1ctre5jslXovJUMYba
hbfc2LR3e6/f5gNGEBv1vHVzaVRTGMy8cQy5q05UbOnjSyqvHI0hCrcM3A+tOmi7
A/EG8AIfXn7ppH+hVOBDhoJJiNJ5sG6h+LEY6Wt6slhIfwhZsGp4+Tn3Rkr7wiC7
21flt0MWNGahTpT9h4tMAKGaM9eeBLt+0n9sz0GaVOWYO8IHhoRJxPqZ1mFDvdjl
pJJKn8DO2dCarFKF1zljpFA53rMM7FUeDkpSC6qhaWqnX5s0UXTTzZLzEJlkEVe8
rgbBtNThoVZKYy1YiHruPzKeIndilliGg/5ROs3p7olMtwkHWUjPDWBUcKd4CC5/
tN44462MMTth3Vh1nOP7FSJ+zX9GTxJEnOe6OIv35MLhe5jF4y2w8xrOd05oBFaU
F/x+ZbAYrLmBpj9wHCCqPVcTlFC1jbk6h4LBGmB0BMUr5STge2KwBcC1MRAUXtOi
EGIKaKc75USN215r9SskZTlDqtLp+qMRnNw0jqxqFRvQboz0NmE/NT5gvHfiAtrJ
vYGMNrO9yxNbZPKkGXnxlBhCMV4qjAsjFedtkvyRE1xy+j2m4YPKn4fAcHBYtUlJ
Rwezd+QWRRjigVe9ea5sQ8lNqNb11VDPTyMHRvPvdqNS7ECY4ie1mEHt6tUErJiE
MXBO+TIsEnLrKsQDn2cQqmvh7Nx1320sAg7KVA4rbt27LyxS/GpNP47GnBIBznX2
igRyO/OJ7CQ7bPk84pblTRRngiBg3WtLr2XHicBmmmp/5BexGnqZ8EO3LJbCLoCi
6umpxWrplVmkL3yyAoFRu9C/N/fDII7c05EB4iH4vegNfdZnPLNMhipXZmPbvNBo
1Rrj0x1qCR3Qk8gASdt1MjcvnB+tCJwDUD16T5Xxt3T24uOOfsU3ud+xq5O2Lqax
rIovRpynfeXhYEa5w0QOaK5ByBTWcUTIwXnso2d5tBTBHiL+TJSNc7npabkdH8x/
y5lPLx5XfifsO0sPZ353+bRcOIJqu1wXl3tGzVurrk96CFcdjuOXZNmU+93Hxwwg
4gAAKLBuqmkGufFf9fIRehHdfUC1cEf2HAJ4NEmjKanBdY5+NtyZiKK8CrS+GvNe
hh+TWHD0kLxVSvIOSJ8hUzXYRp97BPVL0gplLtqG7aT+mWITTfd6ppUJ9VDqmYkK
atwi4IVhc4RZ02UUTxF8/KdEeKp9OvBcS1MCC4J9spKng5seGyxWpMrgm4EcJ8/u
3ztA7Z9jiSnjdV8JgTkKZx4cziAVRdviCzCOKXh/uecTgHoqZaI1IbFYHdNe57nX
E2gJmutsWrTKawZcxXOT22pm6Sgoept9xwZ1OKmLKcAJt0nYzJKzzEISz0htBQsY
zptHDIqK4LsJ5Acc/iCc/Jzomk6LQbkM0dOjQU35PsJmO7rUsXVjV35/VIiu41Ud
itm9/DBKfqemeXGei+EEcDFU5pbowZ90x7xkqsk/pMlSrHdPydVk+TSKFqadSbNh
iwffgKe8hBS8iuq2tAExumxGuWvdue7D3zrsVC09K144LJ2VNU9z4XFxMfEMclBt
MusFANWkVOvhGzX2fHuvVAL265bfJQLx5cDvs9pvoViukt7CnYU/jFDomUgamux0
sNJZMpkyvYFIVfnhQf2n+aoDFe4OZ7xjJV0TiZpENXW95jr2vgG++525UmkUBb22
wbgNhiSbKXs03nZ0Nx0KmkwWB1yAy/ZMlCW/aPmo5ll37eIPVD8kjoryW9Zxfcn7
ED0cncix1fR+UxluRIOymgAF2epyewyH5+xOY8ETzSxjIEL8adH/CEcwe3pj6xG2
9nXMxTfRPzRJUZyRdyjUDxafCq3lBCE2QbHJH5hUCTt+y0qYiGnqQehyluGFiIIE
DaEui27i2a4scdFBH50byh/cgltlzzv88NS4YmHBRpSmPe8LyhlpDbDGeJrUrCfG
+qvsvyw017+zzlnfbEW3ellzF09gYkM+IRpXBNNIvIZasuD58fbQtP2ablY7qAs3
MVjceJebVyqbP5eWem8LWREAn0QN+xSDHpuEoOMZjGUnq1RAKDJDQp8wabG0UvrE
666WEq1B0Q45FkLQmzqwkd19OUXun3B621E02MG6/JXI54q2CPooIiz6W3zBndbc
6m5LK2Z+iuRxl4u3EmVzV/s7Gr9BIzym28C0jrbbAGs6xMa8ajHfI/694Xivbl4W
934gs9ELpWTFQk6ccJxTWrrrr2juoM0eKJFIa5ldBbfkZFwsLY7wUsj+ozw1KvPF
T04mLNMkNdpms4CN2vuxzQ3hIpRnMK1BkevZUytIHfkaJZwFwI81uqcS6e9g7vMZ
RCpI01ShAyXLelsiMblVJN6qQqlHOpTxJIX7I7TGomiyWYfErXlhXL0aW7hyphb1
SMzAXpt+t4RDr5zDpGSWxUsZ+kLD/W5nK06fdHdOrJ/tStg/ta+IZkNtHGzj81rx
PXuJBdynkMUxszf7Wear6D+WHrOXV2NxbZJZpjfj9q8v4AvwjvLGGRUFwyn3QRf8
HH36q5xhWpd/CU3lQEUYVmRcgF5vijgX9p7/sNus/QZz6mWSaxm+RQFS6M6+32hi
jaYatX/apxnRD+XZABsLyfs32gujZry8wL/CX5AXGjc/lO/UGj0pCgTcDFgBH2nJ
EuGeLfiOO4Dtw915buUYpk9szfxe+E6PEUY58FGN23t2YSPW5OKZp4RT3RBs/nxH
myYhZ32lcKKLWOZgzSNdccEenDmSYSiFDm4b+pMzjH3Y4TdaRMnptHFGavd8Vndc
CE4yiv6JCM3vf3nSQvwI802GiiMvkcfJTBnYelD2AsK8sFWj+yTV4PibLV39CeEV
/Qe9NLTsGrzZUy2AqM6Gp5zxpKA+tEjjNlN78sf0SYiVGn9qOJiWz9tMpv9Ghzm7
p8Apa886i6twGz9Jk5+1AGo415U9LVEvx/pW5wGX07oZaHRI86xNuyKcfQBOakOw
grQ9uvpOOzP3+vqKBt5jievFSXjcRfqnkJndGQxy6cp9Rr6fpgYgwaO3hphDxU/J
f4TfZdKqraDvAcnSKF2DgIccmpqYe/hC7cqjsQkhYNLY3M11ZyU/py1hb3lJZidy
+zCGV0qOA9oM2oIEzQcqesgKomMTxoTJRr9Zt280yvibDjjT48yVq+OA1cwEb68a
26s8MekjrkxZ+dd2S0an7RKzrFiDAX45s54YM2pZ/VTXNdioF8r4OsVCW0yBL3dz
qXx73LkEzDdFEiVM2kN+RQSIxVVXMODbWG+ZsdqiYdMvb17NsX88AijSQzDNPHNO
GOdhtArg/vUJ721bI34nFibgKIbb6FVRZQIleGzJSIacob4RQAEAZ8rEvj+Btutz
cMa9lfWkHbpeZC9HZ0/8Ef7BWC5xetJDNMoq00LVFT7W4cerAVjwMRMiG/R1q/rr
FnTvI2f0Al+qP29EBsmWmIJvfTejdWrNWmBs8llX02YaT574hLNHV0JJChAKLZq7
jpVSH2qqj0lfsKkBEMNwYOTafvSUXaI5iZI01D71m9M+OBl/q8U1KN1pca01tu0d
fVmlWmB3q+nyDmrr9J+ymWU8ZjCEbV9xxFc5mhKdwW9RvixBr3zSVJpkpwkDz7v8
Rb/gzdwt4/lMGxq9yPGqGm3KhG6bbrQpYW8HFVkFkFmHzQe+Lzk+vmF+tSnaPqyA
cLabAzSui3UX8UCaD/XsOnyrHNW3lVjtEbMckxSW4KYVfyja2fu8Y+EWvaLsNiC/
iIFuneOTsTOVfGAEKuungmM7DmuuI8ZlqytBv03+1fNL0ANR+RJ8xUrC2kXErdmP
2rQdXWfSZk0xZqur07mxU8m8iG9MEMw49P0U08WOjfHVWiy74gZprxkeDM1lRt0W
BYZZplbcraPYmzvcT8zajwxXZ4JqfjDYTEVuS4/L9MUPt6tHRycDBH3hKAeYTxVQ
8jn5+v8THfhGZSTSLTYm3C+YrtYj/eFH1i8/EEP0IQdY/BFwyVwpQbUF7AGXG2U/
Z58RfAOcUdBXnAisgMgsjtY0GAb8yUBxE3cZfPrStAPlYyGTshJaaKRsG023zwXW
fiEoi4dTxmZVjGYAnXv9JPhqr7tD3XhykLXysfgv7ZB9x15YoTJEiy2f+O2E+VxH
78Lo5lPoNjg0uMcW7LfPqp3XJ/lS/IhXHXQikIDUMRyOF64+rR6qqerFhWpf9bFX
0oNS42qosxT7qhYvXX7fnGm20zGAtarF0TJs3jFRt8QCRrFaHJ9kOTkYY0gfANSb
rTtJc3VK3CXX1vzISwvm9KN3kMMLiZVY/AFa08dD4eP2+mKD91lOVjlHiUciqT34
f1Vp3aE83X8l2ouCJFh6TCYtennmtBCWFfdyYcZFV4XZHhEaqlS9xRdKRohHs2nt
F7Di10Aa4aXmohUGN9t5MSRMAiiKoPAgCswmzaDon8fG21Hra+fG64ojUOyw0onI
kPMtmrrxycupUnpNiR6THhOEgDh7vJaT1CL84dQgYMeUtJJ2m4icANDp1QCBfh1j
fcuuphxWWXj7e7p0q/XwWPK+F0W++Q5qLv6dUqzfdpsjbCmxzFhbGwNwqhC9+XrP
DuhgcYeFMkJCAdDye0TGDY3h4daikcIk+wFSmI2rOXW67rRqNcr3CJ3EAhjUrTjD
qPYvD1U+RYhTmN5ZIoAKxdFoi9jZpREh5WjcXkqDei+Y7HRgeTC7rZpGaHeh4iUi
UWDBxvNhWArFxrQsvcVnDOC25EjDkoavirZC1Kq8ppWS3eZFM/EW09TDbtaANiCM
RdlBWTyr5sDYTf8mHYBqxm1vC+sHMOtrhBuV9BmMMYU+3yzxayhox2F2Dc5nO5pT
15oxjLfjW0INRGRT2nevCmcNaqGNA6cWK9VF5lo+qXCmylwgX6953bGt9fMTWiwQ
wG3zELz7rDVmFvVXyGR6e7d9cZOCcUXdqW0Ym1pcWiPVcYIPIBos+93ZeIqaA7Nq
AgU9DoZYcq4lUm/XtuG1hQf73iLgZRjZmoy9jfthF0sNNzyxFDs9GREGjUcLRhxo
QQBwaGa91F9iLRMhX29Cjng+9AethqNTnR2i91qRafsj9eMnLUbVUStaQFKxLc5Z
HfbqvGAE4myB4pN+MnERw/oS477jYNpzNsOTlZ+QeqBcXYJtIyJs97Tgg7uTle0W
i/8PwUoI0uFDw6ffQtHS60M6hrhH6Vakhj91SVSnrkZzX+ZCkUq/Xd+9MKyRFfzQ
ZRSYxCzLpOtIqeSYaR0R7UR16GImNDEsbuO4TPxq9sguxhPrnGzFaZlaC/NybG+i
kz+c0ZoXQwDiavkBRbOCWwODz68FD66h4hpQPRki70oPSemTU5Chwck8RUnArrdd
mFZ1DScHIvniTsQSx/0FPjHhiqoY/HaUe4ZrpIzeXTf76uxpBZPp1EghDdWCOw5R
zs+EN54PVMoOrccR0+X/CkF3xbHoYqgI/DQ6Zgn+qKp4ri1Ct44OKfg9bC9OtmEG
YKvrQpH2bpebC4CBeywbFPM+oQQXR4Hs+6+MhQpbe18=
`protect END_PROTECTED
