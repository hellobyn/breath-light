`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4gQOjtL1xfWlACRn6DQBLBm1Bi2oeyW+DsIMe0I/xfV/YOZl4TTkUx+c65dmH24
jilAFVPtBNa1ua0Y7movKtoco264hJxZTKmLPsp2fxo1WDxYTWrUPZzpnCjZCI4y
8HOA4VfmyaZp1dmexyBmrKPebxk6Afx/abx6A7aocm/tfbHnnwHLSK+llxjcEXXz
16LFoj9yeVZYmrHXhLaESZbbRX7lSr1r45EOmpnUPKSaFm01QGYmxaWgEYLz4lt6
UeLd0o4dyRvERVZv4WN54/FCg/XBYHZZX4h0HmeiU64YQLAFG0x6cs0S0iQ7qefB
6mWg2YIcRMUrTzkt+Mnm8J2oKb3PBO9xKX4MY7asSOOe1fGIyA59OTWrxAJQJtis
RAoEMtT4r540pjz90yyrFug8djiEraoiMnrlBAqtiH6mTAXOrJelcev5UfNJQqHt
/AE3LI/WcfzNIb/l/onQIDb8aiUBTLs9cfVN3cyHYBcypMqB925BLH/TQbC60UM8
gm41B2FUeMuxCJiHLm6ofh7SZ2yK1BwMhMBBXfxrFirBp9ae2N9Je5xIIwGjqd74
ajtpkeuwc2OycRIMkS2G8/ZdQT2XOEqQ+eZgF8y3l9ARLVLsPkwrohKonaVWkloq
6FLQ04I7m3m7MjkOFn/LToirkIxeiwC41I0xC73iH7ei5OOy1w31gg6IkLSEyX7m
mQLU+hslX82QLhSX7jL+mJFuTHNEctnFMj0sKpAuQ5yIJa93DZQYFmyCZxyDvEFo
GwD52EQJlwgtZb7KjJRH41y5WPnwJB9NaQ84KhSMydN4BUc+RR7IkdofWIbLLke4
GSCnAS4sNhCHXOnkOz7vfKiEo6G+gWNu78YC9bh7zYyAEM/L5IubbxcyNwkvmgQS
m8qxUkd0lBQmNZB7N1JMm+G8XXmAqek66m6AvvVIL94Ry1aVW8CeugWq83wLcgTD
qaIRHRjhdt1h+ryaso0j5bLHEulBlgM4WaalYiNU/ZFL0TrrMscjZwaevV03wcZJ
F5zTnCRCC4Dzxd6Jh96ruw3AyyJdAE87T2PErm0TxztEBNGg6vLyj/eexSFw6h+R
p8rvtyw0CBCdi687roO7mUfDYWLUR1Hr2qQRpNRt+iAMjFe1YEEFlwDyiTDBeYJj
Oc3Dmr5sT7GdDP1EkQllO3urvEx6pDMKz1tGX9RX7yFufJ4Ebhtni7nrJFN4Z6/n
oo4IMGjbw9UQ4ViHAi7QkibHMPSxJw7xFAnGTQcPcjm+aC5NMmAnOrEyPgqxLIgr
mJqtscDBFhWAEV0g6Bp1eyg31jRmE+d/ccjIDp44K0rXd3/UdsQbh5dIEkCA7fBj
HHRLxpiEgpt9DeaUhDeamDmwA3bKMgUXBlS84l5q6T/6uswYrfb+GsfIfNa1PP5/
UO1rmIyVaIZfPs1v7tBs5XakbYUBpvVmZLAIUZDfEbqWJDIFNyFIOfRSwhWmkkR2
+QmifAPjhDOCrARoIwnVLe5voQH3xRNCyj/XG7cVjHTjRT0s5+OM9rApvnCts1kM
a4vBacST2HF1UhkkEu9WldZ2bbAnXt6Hm3M5sfobBa/XX+4nAOmZLpfLiKldkRSB
s/+KHc+dbJG3ORqJgtky6HevabVQwieelxpoQdvuuPoiQszp2jP/1Psvmys9mDNm
Ueu2tcMJN1TzWK9sFvXcueyuYkStR3RLz9pEsDTHcN1qLlTdKnYII5OQYdheBBSk
NBFje+y2PzW8XPaEqMfpqiTGVUBRwafquv1d+w1AQsjthI1+5uVMmG/cN4g+JQHd
qFyBYssRWU6V1/Ae+GOgeyFTWjkT+bvQLrrSwYMUFdz69f/6wqUkXHCoxDP2EJW1
mHut/G14cPM0FPVRBuDhaYUsCM0OpjUujPrxgD/sEUhwFBaaqVMSuVCCxmUrsBdf
SWRIlkZDrm9HfqPd16u9FP10VYlF9IHeYLrn1ZcwIX8zGbrA2u6+qSmy+Nn3cHWM
UcVb5RvsIjx6zszjfhNOtqopWXdGyzVwOp90N/uYoKEeozzBtKSOf4ZL+lbZW2U8
CyT0zAuSwt9REEIZe/soJQncvhVj+QxwtqAbbEOkiyGNVjZ5tTApKHd948UscSSk
X4D8vYiprsdkVy4x2D7Ww7E9rzU0TvQ+zmK3cTXcDu8=
`protect END_PROTECTED
