`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLeLc35cPaTNV/YZTRKFjxqFvE93luo8DgAGTb4DMqCFuOtPHfnohEXY1dGLVkgs
d4dTPn8fHdau4a/4pANYnSrGrCZKKUjk0843VjlUtxTbq/u2MdFrL63e6SVNAmb1
mVqVWt/uSSGMrj+4G944T0w2Z/m8Tvkp6xFeFWXW9lWXmEMj+kUvUElEhW8rW62w
tuKspJhfmmO4O+iHI7a3zrJBXBF1g6QtNpJeA/UjctL4jlyXcerwy3vLdnnIYn26
gLJP7TQOfMtB61hTQea+e4OMKBr3EuvvYV9MLK3H7jqQi+7ueoogL7QiDOnZ1VSZ
QR2b03NJEL57QpPSgaytk9b6vAKdmiFBI7tEP9++3KDOP6OLYy/wJfNDcRCdbkBr
9VxIgxTb8Zy2Yv12E+/1ha1h3LbdI6qsePSMBy/J3uoMUVoKtcld2nHJvQKcUdRn
jFsYtFnreGP2jnc9ptMFUM7G3xdG5Jydv7DeMNOd88i75Xetdp6qkZy3lIQjDRxp
DjHVthVqH7fU7DwTc2lOcpihl+CLW+FG0Zcp/ZtalQPycZ46txNi4nLW2OcvupBZ
xXAkixNu6+5hS+8UNCurg5sUYHXuFcQ5FBXYRsgyYVeqRAox07sas+fDWvvOuPnG
LFNzQm8g5vD9ULta2aGkuA5gCKz0CNDM/3RzNdwYA8c3GeuG0ttz2nfTSJ9QTOSY
fnSyuh+TCre+vVYGm5J5ulS4Hf+B8NrwQJArDlz3+kVb+h/YYqC+Dc4qmb+n1k7c
SCvTS0EOlVaBqeAZM7zjb1EpNliMYg/UF/Ih26RTLp9mZBB0b+31+6HaLGb7PIiB
l7iaJggsXF3jkPl2UblLgRrWTk/FmSpiLaUFRJDFqQ4UJ/KxwpY4wRz8PdZNbgve
rpimKvYRdm0dLohmaTL7Wvm2asipNaq2zsegaf3AkBJoKoy+RtFCZq+ZnGdcvvBh
YhY3YVZXlQ3VU419XVk79GDE94hgP52xHbNCVSoBze1MqaGmsX55xkvbL4p3ME0Z
BuLhDgXou43NKzNd9RTJlwR5KtHN/o1Q/X58IXIZGp9PHpuEFCX6+aH3KuLf5Tfo
o5ksrKsJJz2UoVtXxT+06ihA3zhxzpfbPqL712iwg//OwViHyyxUOyHCEl+A2Z8P
BPPPg5OM8qn7MmLUel+V7Ah4DiEkTMwWxeRsjyiPGy62QeXUxP2hg9ugIj384hsd
oaYgA+oJMclrQli9yQkavnWNDSTF4/i5JsG0DsEv19WMiCVcY2TnzDo2TVYhcp30
jzNJJVndOOVYYmqHXlW4TYCN9QlIkwNzP1XKII7wmZ3RweTWTSVLGKP98UufLCnY
cPKf0J16Lu9dSyyKhclklowyQkuKT4gXWL7lJhqdzm2xnR7OtPo1kTUqxzVp15Tw
moHF6idkYC3iH+gqPyxOMkIJ4lkACfUboeXFa7GqMe1TB//2UdTHGpDUCXbgmmE3
H65td3r0szkOCR+RFzbMQ4oL8u6geAniszXtqVJIpENSydz1Tll3iEqsCejgLIea
8frQ5MaKyg/l5tNfG82c17BdsgbYeBcF0hUnCrpt3GvoAyNuWI7bPBnaABepHu9w
J/4AlYqMlfJycR9FU6mIZxcDj0sCNi96r099844fyVJiGyEfrxXgpQD051KJlp9r
S2diJo7OaT3I/rFYDmcsiGJQfjlr90s0BgUJLagZJoO3woVOPuIQy/vb6fkcN+5z
33wYpeAJFxmZNqrCJE99V86o8BypdZo3x0gpaO+W4n18s7NpGG+1/+Qn5Dpo1juF
NT9ve77KoAdtgaygP/yvFviIcoOzz1AGNt+LHz685FmMr6XUfwsEVjXMO+BGsz2A
tukzlS7r2Mb6rXhSmiDNnL9xzkLP+KEMiEoKQwNsVJ6/mrdTroqBQJEqreNQDa1/
1rUicr0SMIgLj4STxSqSl7yp/DC3lbqb5vGH7Z8DpAqSUpdgxlH4PN+Getj0u0j1
o/p0cQ+gJXfOENh2ENhNQiSMCc6+0IqjgstADTKMnoEEeYj1OOi4UdFTsqMOV4LK
dq27fmII4HhWjSBu/BUQ/uwzyJ/MhRyrpwCbGHDKiWq4Jgj8XV0nob8LZNG7LqE6
VszYMgikMtZ4FLv4w6JjHIpkoIXHhfNnDH/tX4GhZOTi9qWW7Yzx+AvWeqOEYclb
eW/bxI2SwjUx/ZPeyumnOLdGd/Rvi1JbkoqQrRKwerJfcN8JecviPNzhBo2qaaj/
8tV3i5JOoswDa0iIAkVloQ2TO9CYPi3sIBw9QDq06iaRh8QWxpEOTO+uL9d7NUrM
76LqufATnsqTe28oVplcgnOhen28nkYu42icwHcOL/d8LuZayUCCNaiwAKi4yP+x
oh/z1qOQ8+Irg4sKMQLECaMYsNyRxLMhf4ZHYR+KsClueBs9Wxnu3q++VdoytUwG
KQ9iVwRCuM3s71/EZ/MWEPLvIrbVfpcmoxnAdDpdtSWI/fJilJ7wKalmOq2hnja7
waNfe4lB8EVJtEzxVWXbPobQghIpLPnmTJsuS+F8bmEilBnWxfMstVtE7QkGf5oW
7pDfbOLFJ2xJxhyXucLAojj60OUdYvHfIKKJxVkBEYRPafxIr81kZABorBq5EGoy
vuDcZAljcnNoIhuUkJUBOQ==
`protect END_PROTECTED
