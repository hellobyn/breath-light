`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXivA1MsB9Y3mhxd7HeeygdxwdGfn+ZdOF+nPBdQqCNhByaQeEXVH+W6UbQTJYbY
F116SV5am1Lgryuu/PBVjqoLRHezIg3hQFaMBFG1taQqFrg8aiuKY3dhsbalYB9P
mduWAasIWrYcPRKFL4spNOSSuUUG64LnVmY5e4yQXVERwzagZxvLa9Y69PdFqQSc
BJa1nahQgaO4SUv8c7yOm4f1hI7OZBjMfsv8nYfDbyrBSq3UIpinuQU38ty2X4TD
mEpvmYhUQBZw92EeDDHrgzVavA68LyZopHgpACqLedSpoxwYPOdX4q2noimYZRi0
7Azmx4uc7dxfCV+/fyFcBheYKxWYY4C78u4MTt0Qzopua9AuKkLqM2KZB8UYis/W
48WIJC/oSKpJ6OWAxmphDDYA++6qNzkEe77TWCsmRKVWEus6UT70JDfZo7uGR/bq
mi8XfIXZAnJzECctzugqcQ==
`protect END_PROTECTED
