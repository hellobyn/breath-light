`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf4PsPjkQmovlGG6lTD1+YCWO4ZGTZ4ODiCPD1tJaGha5RQ920QejKcPywitnFmo
0RdI38jrUratGS1OH/oPFznBXJLcBezlt5fmKB3kXS+ngp0lsHdABJrFZCe/5eSp
veJhQMAxTPkkzkFkRaCi7NL5k0N6yZ7ZvoSp9Ik4QBq5RK7uRu0uC6TgSC09zxth
pDXbZ/1ARrfIXRXHt/sMR8R91c06MCwp5eOU8X/DDuae2x71rqR4QS6L7X47Bk9L
H3lpTYKcOXadujh90zBV3XnS6MpBjQEu0pRXAhegfli4FWQoFBeh1eqwBktW0ppU
9ynuKK0FFcBzBKshvNmRdVtFJEmzhmkNSsIgNsx6TlPiijtO5NlOR9hwqWwWQd9b
KZsbgz9c+DTPBF1NbO6ZFhcmlj+feECKklfPxB/PAPUIgaXuSAI7Fk4rAECOKrE9
v4FVuyCVXG44FHbhN1YGaUMhZvMhD0Lp7RxoYaYvXHigwWaE7G3P+h9wozmT1B1m
CUc1F54JiSNYW+lpAOVo2tBaIgB2f1ZHz0l9KQtQ8BMZyKrpVk21LC3KFEZdhL4Z
RhvMzem8dQwVuNe5Mr0s+lhqHldnlHw9sVQy/hkXVjfSDuU0oJssjlqdEXWNvO6f
DsvTuWEG4c3dWXbtbtj6P6A7CUrat1tbHDU8kZIqYKUN0S0h8U4rdLQsQoAMSeuW
PDP7ITpja2tX6K6tn5n9aeScl8huTbW4Dr5qX65XJGU=
`protect END_PROTECTED
