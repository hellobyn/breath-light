`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jabFAWa3UMRAT78pYkTTTNaSVRu+Vj41+FkR1E4Z169xVLXWVTu8U2ZQ8GTmHcwa
rKAG/qTNEU9u7GAl4BhF0y5sWIFuJsjJn09iizp7BDRVircrrjmcwHDW82I1+7Bl
mnfkgFLqIjLvdqZWzd5TgTW6pQLX6+nxtfgkPaCDCjJSPRBRBnZC+rhlyKa2AI4S
bL7s3zjuB3Kd/4ZIA5Y8mvgskFpJYesZ6UYihswM3lIdD2ScMfDPvzt3t9WSeiUv
TzYkOughUyPXzNm/+rV0agFeRNgFsCHXNzFo9vnKjj8HSSZ1NnK37PB4uuKsYDhV
2RiMXfYj9vSpqMaogpfwZleMF34U/AJSJ7GgBNg8+9aSQzz8i1ZPSyp7n+CQlBYJ
A6M577SE8wdnEQ1TJUc6ruBa+JbyUd+pVJg1RXuQ4z8iFCtCc6v+tQ7ucm19NlsG
COkUkyM/nUbQuwGtiOerf90PNt2ReTUF5Ya0Pkb0JdI+yCMcmi9pEG3RZ25FwNm5
zHWFkWLtxuwjlTsUJQHo4g0ZASpNHErm/RsILR42Iuc/Sd3WTTsl8EE8o965oSkj
VuFZ3zii5c37vsyDDVmwAvTaD21ywIFuf5ar1mOHmlsYkwRHDFq9MvzMzDUksoCR
e6ZMXtTaw/xanS6SM+tQO5FuUbqVnCLR6dZ7XjaPAqB4kCmnaVbEYtLec1PbKEin
dHlKRsGUKyssbploDd3SiymT2bnGLaRqhbi8VwwGhkgSOkDKA4+y6F2uDInG/CvK
bZujl3ze8jQs7VHzSWYRX3WRW2JBAnb4n5W3DJKF2E0elzUet1jHiqOBETSdw0Zk
/UZStWcgvtlsTtn2dah26JiYitxXFc6TrvUDNgzVz8UsrULRmbHrk3wyCJTsmNvx
zulRVeXgVmFFpR6Lfd5gVtokAsHYOkkMzZxXaAwWDKLJoH7cr1PnhA2iBbLsXrUF
vlKX/gKvc7izw9/wJ5sISlR92Ul0Xp9Gocp+i5ZWtR1t1uauua6QUnoe8Od+t/Bu
NY3AlshKMtg5htb+TmTpC/uqGQhT9KFDi9Xjt69tDs+TGBFktcnwXifQWFw6/qS7
cAaFOeW4VNqmbvR+tim8HtWa+mWVkbmtRJRn2iTx7/k8zj/VyAvfddta7rO9Smka
ZlFuIj6QRl+LSGcGXmaaYc3fyz8P+eIJMLH7HOLl9ywTNL2MfAwZwp0SDOkoWeQA
Euy8K7i+dnqUCEqsV7CTJtYDInzMyx0b953cP/i1MFt8ppeK1uCQlvzetvsXd63B
Uz+CUpWTKQg0ygBAk+DqQC5VXHdBrombuSukLOJW1+zQ4tNp1J+ycDTEA7x3joLK
8HEar0UHjbp20uRBhOPVG9e7MQrI3kXphB0blrI7x+AY0CIBPwhEbnpxY52mK4QW
vbouFcNYUCcJX1ncrj6SvmjPqDNVcaO1YooxLBXfMNr4+MYLMXY4i3ORMpjEgsGI
22AFahwKjjOUUA+xZSAP9kHwPkaTMWr8PcMekbbP1wXqkxsMQ3p5qaTjT9YqNUbY
r7oIUBv4OGTzHDdIzoxiw+YMvGUIBZiPSA5960qUZ6IBRiZaY5j20Rpue/g5tzVN
Cw3y2C4Xs55Az52yWIaoytlSMDA02CjUY1yPpO9JIlu3eC1F4xwzgZocYy58kFjq
erzCFC+Xc4zUgMpPZytAE9oyksTMiEs5SxDHKDOImiMXYexBat2EcyvLLz/IYMKF
AwgMdyfC+VnnJQNi1uE6Zz108KWU/TgCRAv5PHfnxoxpmYPdctRfqUTSnD5AqsQU
ZuSlQAQ2Di19gwxAfHXNIeFbhagxsi7TRaYVNqYq+O5odO4aD5AHzRRTKbvneqx3
M9S30t81TuiXS0MvGVwJexbl+yrlUVzFVB8+seXgXTowFnVhyiePp4kB38B2rKuu
ZoFdSP7jMAkFIZf1nS0UU/Q5ExpkReMu7GxUeOyO0a3eR7dWJHA1J+gsVMsRPuNj
Lruu4XYWtlWMvWg9PM855hLovF1ZR/QPDx34hyPQOk6BC5PR75VmvuUjQ4gk2vbW
3DSXwI55fpZglnOu81YFrK2DkFptRrG9D5mJdbpTEgvXdeYxAk3MgHyX/OzfiMl3
I/hqB4Rcni85prOCah47EcrZG4zEJcHIQ9TIIYmpVQO4udzU0fHdHK6/Wj9WY0S1
iH2iPA2CtpMI1nLqMYwCeSO6VbVXE3kqEHkzjlspwya6WAk2ddBu8Qqc4SF8/7Pd
2TgjhL2lAYVte8002yiSJbhYH3xMLTL+A/ipneDMYcw=
`protect END_PROTECTED
