`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvYhvLKZ90nPI3IUZ2X5to4RWBsf1a2mzVEZsmoaK08IdS+yPHTOb++mrhIHiMRG
ZG0Ab0v/xg18CYw+sJJzAAoTEDVroY+gzB1l1FhxMCHcqHjXpejgj5oLIRnLthlh
5waFlVvOM6QltTe8NtS8KZ8mRc07TuXffnzewOjHQM49t4AWSBjHsCfAt2/iuapD
WMV/BEin7l0OQdfd+uLm+LQyKT6ILnwMChwKpzr6l5RxxOBN3Ehxa0li+WGE4V07
b22gS335nGOPTsVcTvI3DQzfHtFcqxPv6jFkmBZ0Sw2wp3JBSjb2fPBSLxfm/+//
IbPuSEhhHzHYrJUw96fZ6QrqBu8p3M7lxvhx6PpWjG3WgtBHGkXQuPNDfRv5jGQG
WhJxdzPkjnZlBAGJPbZ8up23MnuaTVMbJXl7d224aagO6VeU2PS0pevI+KtP79/h
qY5dwpOPND30iUHXaa5NObrYE1P6kWCwuAdkdtzhtd9xZO8LN+jeaHf4DKg52jtX
dozP1XxY4qabBTEz6cdF3fkDDGg4R/gIJZTFpIl7a9wW5vnhACSUMRPW0lpGOhIM
AEWpiIB5VBsq1a0TEnVySQc/gtCZZkh/UNCFfppY8hQtAFN3utkW1Fo4ViDurijP
gf81fHMBp2+wJYfPqNNrvcvif2yo9xbnYrQpUVlQfCFZfsdbTCme2nXPLoTvMf4k
313kEMiAKp/LmuJXlBgnEI9Ro818y7L1lX2/rkdjYS69IrCNxJ79zR3N0hoCvHb7
+7iQLnAg3SSBQJfOn23ngtqYL6bfCt1etQQHBMR1oBGMEh1jxTjkJzyi/bDcPke0
L/cN2VLJU8brnaVT0POtkW+KOGbDG4APmCcB9MqTWD4htjXBZCHmGC3i/LlkF3BY
nh/2UbQJRq+CTcQdzfSuNvGMUs+bBkBGF/eVFbcOMJl1jEWwi44r+GWREWkv/IZ/
8LVPTxOr3oBeyaTacBvNVx0o2/K7Mq1D0K3SLsGh4sdG/fYn3jFbCOpElvZZiT2l
h4f4FrhgnGEAHch6GF7i3rj06s1SN07VNanIo/rBhLcUApmr8xrnIw8JUlDSjek4
IxYIbhkJRvhARfk5JvtPWOHcgMG0ImZJ5nXsZjiWTtiqynOfOoEmA8Z3t72I3gZE
MldT4t8GE+Uj9RNKExAjNOKWChHTCrKJf1NKQhGtehZFM7eBby/3UEykihoTc/Ou
ZOs3VEiGERoE01opSs1iCWvDWe/lsCYi/RZW+iyD0oU1bBgeuJIgyf/CNeQToAau
60Ix8Q37lintlAN04WKt7UVsSZsCPWBYux7AWF1xxhPtwXBcMCWgMJEQxoQ4ZRK6
72eSgEcD11SaKSAT9s9diu4XKsaegyQMeo/Nf6sGly8HTZHlQzdhFGUSkdRWQxR7
jMWQGNRdWRdVud+rNRr/EgUOSTTrXzWLDwb1yL1zJsH3SEKD9Bswxh6rTLC3x+cP
L8y0u/wnczOgUsg+QKEcYW+krqrWMUJRY7crFwxwBAwB/eeP2cCegvCAxdYY5GAL
HBZolzZB4uH48c2azZnNr8e10Ci8o6i2UHGvp+CuTh4llcqVrWmsCzlhoWl2lpo0
5fs7apQAUXqjFBMbLe6Wxo5Lhugpg+tlNMeLTE1NwExQhZINKzGUKXLxeA2WgT1s
4p/keWOsNJv3oEXsjL31UzoAtoq304SiOxeBI3YcT2G8dH5bMJthBAmsVjPMcnYo
Chemx1EO9ji3Dll0fyN302sUh1wvv2m3cahBken0LzWD4UUBktc15W/VGY4Baj3k
vjkg4+qJg0hqmIqKmgxBfx9XiRlByElwaxQJ5xYOP3pDT5sh7nKgSm8OlyaQIeCY
Nw2J6qtFkB4K/ouvsZf8FDsUYGrqVWFNSpy/b4kbnridArGaxV14BEHVPxQ5vipt
0ky3NNDhiv2d/00Nl0a5WWvqxSNMTaOTpoIauFVCinmC5AQpbMfyB3pN9Odky0CV
lsas+yNibconsnZJ/zFryAuXfHMM+wdtbQ6fMcWnAlXMAJ1NvrAphCN2AqlT07Eo
uMYPAzsgEH7gkZhVzX3t+hTpA0SRlMaihfYkmApwLWIDYZpUNO0GrVpxOXzuemUP
CIuyO8ERCNTQntDf8f919BdaLl9qwV5V4XeF3sTl5qJHTrlvJqBtdha6/Ka4b8IN
rwKY0ppjs4SlgudGgWIyX1mcSjKh+Mj6RfLek0RF4Fr+KtODPwmetu1rUtOPj/J4
TQrLew9We+VIA3kqae7LiGJNP9iGoPOD+mIIz9JHTt9X9C1srL+kOnU5Av9hN4FD
pCfmAz/arPhnItnrTEoAL1pDoJQ7oeNTPzVRDVKxUUiBKiEY1JsrCke+LfgVv+os
d7mNAln+EXlEvPawIHT8Fd36Zv9xyfVOqMybWvukjtsNsh2yHOhAGikdFGTEqqxa
jjXqZoEMcPrAxOTukeQLI6zvzIiZPEOkaN9CpONY9OtObdBmeH/m5E5YELIJ50G7
/ev5rVHZfIvE6ExuSP+R+r/O+CjmP4gzIGnbWy8xMFDNaBg26zKFofAudCD12Ug5
wnnufv4WiokYSJzxC6vxNcth3IqY0+1QslsmYCkMK47JEQgUGMtDI9ETHuXq4hCo
sJF+Wl4WxSKPdSG2xBJLL89+hKKkYS0lyWIl75FcbXuEj2pYDD65GhyMNV5frZy3
GBM24XX+cdzLj1i7a1HeyOG0QezLL6ZkiBKSEi8eSYKpIlaUadQeto6lNCJ7wqn/
foWQeHJ9rXXMp1z644Vaj7bwcFmskMmmwna3ti8M0POBS9quOEQ+SLkP4wuWyAdX
Cc8Lk5xCV+/lwW3ks9vpRAcXSDylKqoLVKTgnWpFX0kxJRmB6alGGtrtVHqDdSQx
WeO43IfSH+E73arQrl+mDg==
`protect END_PROTECTED
