`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbEsjIpAJ0nURzhNRmAgNkHlCVMRnH3IQhUebPqiWwAQrJkZkVZCVI37GNMnDlTM
X5HnajlXruIg8KFWQqTPXq9crZw0x7sivh5gaQxTZwbOKwsuilcBGDtflcrWUtd/
QG6Y/UKAZpA+wpV+7HcuiEGFjr2hBEcoSwIyaxgM/7A+K8DE+fmqRdafZ98z6q+G
GePrIJovpRntzCBpVcl5NmQ6PjP8acP68L20/a8qRNPsFaBrpmeqwl2NV1TcikyX
sbvHC9AsJ8/6nAdpTboq0MUSVQrkNiWvsPaDfJJTbFTGnwx3LUVwsVDs1dm6ulVh
E+Uogjf0u2jlUVuDREqk8M2qx1DX37yiQzXHelER4OUNXjvER3329bh9pvOSQMxO
58ITSq4sweVbOHNTSWzl04CDUNWwDXn/YasljD9E3lrRk2PA1IhyJsiKb2+4jurv
8ZK36YwZuf0tuact2U9vjFMuYCFB5jn6yrb6YKtLmaV2PBTcTwbBVisIyoMHPclA
PyPMsHfHbCI1pn+2CjRKWtb6gB8AgH+GelcAhlZTNvFiODcEnuOn/Uqc5q84E85K
EAW7X1N6eSV4s1v4bc1dvVqMWA0Ln/kXWcu3gsrtJrYQ2aFAUE3NYE3HFFUQm5/f
e9P6iuUyjEqz5Usv/SOtJCb7DmBuP4Oo4D1ldw5D71CwdFPvW0c3DBiU7dd/cY0l
ut0miC36kCQvE2rvdDuVlrA4FjG/KCGUEC73A5w4siNmNrhzAT4yZfihXE3DTFtu
TcyL6PVenBGc9xPng/LLX9nlDAg1pD7T806SkahTisHzWLppo3mpbqbH5jAFPIOy
f/jNIKQWuGgDrVaOh5FvTNC13WxHGYQvGJebMs6j65HeSONAbjgq7P1vH8MSiKO0
sRvwTb/9kPQBfv7HhINwRv8u3/pAtY8rz8pi1uiRutesJX434pGEooPnvos6IPfy
FdKBCK5qCXrDsJSFeKPT/MFgPDIbl9LJ78XqO2GCeFLbk/IJ6BoeBukyQGNBkKdS
+46Br9CX7+HiXYVfLWf06rtpR46Z8LRelTFhUOfLJ4ABZE4R1MSpwG7sgqYz2mrU
AvcpDzqESa31C4boI1hnue+kx+DREUOD6gYB5enivZlPKg9wFEhX9VgFOjq3iFVs
vUeFxSD2KoPoE06Hpzl2EE7+gO2z179GU4UkAV1SKyFFnB2koCgHl0wHnXKVRV5/
kGD+nla4TD4q5BKmyuveFX/AWey5+hBzYc9qRio/wINbOHGIQcGImcOYFRDrBmq+
dGAL6HHUCL4IzVgJBn4SDaoXhjzz47oUd/dUmK6AN2kvsqFgKlcUvDsiVdMlcnc4
qPaHParVAiLKq448u8oHJk/OXLDg7qvxST1TSTazHQn73MDB1XmFToIZVogLwCmA
n+7nyRcev88T1X8BqhxMm///maHXp0vWiu9FodIEU7bteUdKiLz61h5zYcf7iovy
L8mwJVSQSIm9iht26fceWkpPY/DnLGVgTv/AnZ+DHy1NPIPlNpFv8fohZ1gskX78
BkDHAt+qgHMRf1OZEXzRmFYwVGiNlNqtffxc/1Lfg7fr4gd3upFFJdFCElhPeBxO
wYj8rZVOKrIQQEvUwm7MF3YxW+StWB1uNpRfN8dBBj/M0WtITrpqm2t0gtb4VLYx
RTG+aPsCKRYUvqzt83mHI1Ahy1qHXFLLtqSDSGmvaQrqpmhvKHPsFteYQbtghmDA
aG8PSM9wARREvwfa3FgyZIuxnsVzT2DoxF5RwcMQCnBxo4ijisgntzDVIf99E957
iALRYoIZqKs4OBoBWsAbKvE4v1Cc0Vk7GQ+c9Dhj/uMfyGjqERqS9XtWZNOCBtoH
rn697vuajCusCw5IRYfBtA837pj3J8QWEc90cBa9kt5nALCtWIDSGlrvMoELHoib
dBtLHG/hqI21QthmS9RW4H8zmt9uLab4GDx5PpyrsbfXrWQSMn5c7tZAnHBhwGus
Vytvuxivv58go8O5CMT3LLhLOygZ5+iphi5lndznRI0XOEPOk2nBfkOvLvo6eiuJ
G3HknXLhXMnKHNIFNRr0jtlQWQPRvRIxcbJOGF3WKyna5iWmL7BcBqXSaJT6wltN
hM3VpXJqKkRUg0pD+zDlCZdfntgmPCqACKkMF/pshDC91vVtKSeZFSRqA+e5Bz9d
73+HUBL+7z5g0ASN47qtMu5oyD9+XZ+Z9kyl4griiu5GVjTFHfpVpgCNsN3nv5lb
s5OTY71BXwJpTCAauVvkv5fMnl+SpmehkWCS9Yax1+zxbD+93jyBptgkb6VCjB/D
ICzBydJQgWWE6f6Z8dzR+y5QogVhLpczMDv9kJ7iXG1IQjPr0cNtcyJ3DEwGW10Y
1QBJAIiip3dLgbF6/vRoTS0Jx52C9iolvCIZO09IpOJ8a+IandZ4xaaNrueZOo7m
TZNU+wSLssbR3yHLgjZ94zfs7bESto03j7TMHVg+A2TYhV0PpEh6ronJRFMrK+5c
ozPtxAY6tvaZ5p2y00kjwEr6IJwiNEEJ56R+2JhGR+4bkcnYsZ5wxUwhFwMbI9Np
kXcF2Oyu4ucqUR2c/CRIM7pr7QEeeNEnonc1dU5hNZxALGQXLeGIdqnRuSyqtmhk
Groju4BQj7Ow7vQbkT2KI5YYKpgAYWmaFB8J58557zd7DygugFudg054towgwHh5
otwNAeRorcBEhvek5x7QErQ415QzSjM7/11zIqXrBBrGjyl/sQx2B/+tYrnJIjmE
fhDdi2sIqjJKLfTP+qvxUTa4RpBJGnMXwnZz8s4P5ZC3Ached2jN0SyLKNxVHLUl
hhvCzekRUvTUSr3J9FMM+CIEhsk0mG9I5l0UKE9tEcm5/ca1zuoMswr60gWFnf4R
Lz1WZ4CdshKGA3Y3fAV0soRqBq9uB6FEbL2assNuivc50y7HGI7oKDGYAm+Xs3VR
VhDZiP5JZ+g85WBLv2hx3Y4IFNx6CkdPsRNh1G9O6HG6gx5OXA4v/LapyPF5qVLM
sMLRE/9KbW4UsPtrjET2USWrYARfLG2fChhanjMQbInzVVAQZ0vAM5YLe49lDEs/
M/J93gDpfvSypeYaKa2U7HZzrJjwY39Cv8dL7GPyvkJdvyRYcpZszZBOT+QzFIny
m3igTOtME/znkDdpAAGwCCbvIeqz+ve7onNqUgjaJ7zsHAJXT7+N4vOC8oDbD3Ht
d/fvERRULlfuLz1cbYN4Yh9cBJFKoM1hSTyXxooqW+HXgh+yuSkCmkPZxhnDdi+H
Vb2Gz+mT0f6AMr+paL/8FuWlXTBm1KwLhjhl7WSKlxWB5acTr7Ev9RIr56JUIN8h
j2CXP0l12dCNT2nx0Zei2arFCkGkVvzS0Zcpa29twQnokkhyeh4D0zoLjPeGxC7b
WIhyXLZE0vBK43nPxmJgewZx+N/5yF/e+PWUliNcqQUfPsUoSW754BoKagDWBgq2
ZviqyQ/66rPdM+7sTpW+MF591mvKNyEiuAkqwHDoJtmOQ5YXJtbMUUWHBNQED/b8
/k+VRRCXFpS4QTBrPhYhstBhNNISIR03Of/pf22awNGF+Cd5wSkqBnD5pwRXN7ei
xS/8K7wOt0likQkL8Y5B3uPuz+ujJ3Dx+lYbLSZiXGVoWPLTZKksghVWIOYd1U9/
Q3AjwjBDjg13Sc5NyT0uwJ44BG/mlxGmf613zp1FVWVoFF2MQ8QkaE1K3nIun+QJ
7qI5k7v0r0OIPANjSdCidSVUccfqw5uPBdlXG+gAWTc/20wfAzRWfpabef9auwHm
xKYSMonWle0P8/Otp1sLB2dLxKiPxkVDru4m8tEJGZo427nWfSbG/qBs35IdEeQA
3tEzrTLFQJJQLcw8f/afp5hg7pbvDq657DQcUljAvK6lgonjQj3RskqDLIaasnVI
iVDWLqxS9YLuki5JDKPnEqkfpn8oo6QDRvNZfqzcNRFsP+ooaYUmtAZJUL5BiR1J
PTPq8+lw69rpr6EifJPvA/HX6NDG68Ylq0/nbMvLNiYHD5DNvWyuZudPLD+ZRu8i
2xAHhfR+qUTH+CDORzLWAD6njNshK9Dw4QhInU9PGgb+1LKEsnEU/m8A/Eg2PCtB
YlY9dtg9TllU8NK+eGhURBUJDIgGZvWlAWr8hZ39JDzI9kUXw3N2UfUZQbg2TvC+
nbA7xpyDueGhoEG5+yi0ux/CEwry4g/kfStIa7PDQQ5QUs9da1Mx6hYZA0LblXXq
UcelBbBkBX6sxxWOeHiD+Q1u95XC6Jls2vtXCCoO+XgCRu0cQx8lea0U6YUdk8wM
ee4c9H195BJ3aI8ajko13LgO5Lz1oSt9NxeoZuHA+0W6DZNVQjxNr5AmhPDrJ/Qq
wpGuJjDGhDVt2uxTdPH9sr3UEeUwXI2QHDZ8woZ7BbYS0Hp6GTpOVwp4zjt9M/In
3/8y4Pm/3LK7mHW1HScarkQuuIZNrzhgyVacHTbwommj0I5+tn1QAHB14hCEFcFf
f5cP1/Cuf72LurpzFZMg22qeuGL8e0BtCRTUJV6pWFKu4XezJ4UD5Z8OBmagDk4v
x4T4e6CgqgMO3GpL/8pPQkjkV44IWDuNSUrHv5pcoJk4Fjm9DR9QrX3+QLxDBdMG
nEP/w5ICgeXOFv836HkXclUSanfc3H5uij60/g+oC3of1y3eYq1cf06etSV7rGTV
wvfja4d8n34DQKevBUPLQXF9uTlZkJ55zm1b/K7oPQvrkjW2JskWOhg6H7K9BK3I
GucWIbPn0gNmU9hXXZIXyBTzPC6maL4mRLHCJEMSzujPkWw65SjSmDVGipWMFMTp
c1tnOvPt5IjHL6Ut3OsWLHUPbgZbgI5zhHsYxliJmU2TQ8u3F5ReU3XqGI2dTu+3
vJnWUOMSB3m55LUyl24XZxCfb4BOBwdVFf05M042jRJ9wJp5D90HEFAxmAggXQUF
AAP/o5RU8kQdI8lbYu/CKWxArVFEyvPeaE13pZn7ebZiqMCVmQbfJjR19N68Ggqs
evrsNxELOR8NJ1vEsCHEi5VwdFU6WomuLuDc26ztV8AHsHTfnQulhd1+LAnaDvhT
go5ye1FMVpvaDTEGy5djTegXS6/NObA4a7zXGPueLEqZ1oFOZaDTgcWsCRjmdnbN
vd+ZKWPJWSeE08cEZOtwolPhODkVKtvSZj5LklSvbVbw6lDMjtlJwFTCg+mouKpP
30aA0vk+Ph72fwCLrh6O0CPfjGQds7D4DYttHgmcpnZKYj1HsZkyne8rSzng/eY/
jeaosEQOmly3wmZT4ymATrtfcoa1R3+Xb2TwjS6y6+nkOy+3bG/N0adu6ld2weJm
`protect END_PROTECTED
