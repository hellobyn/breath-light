`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJ1xn5VYAsJEnSdxR8Qyq0TGHl/Ukq9OyUj/Oa5lcO6sxCEwPYxOAcSRoMbM/mFj
q+TXkmkOSz4QdsM73AofquDThmQom8sIIkJoSn6npvp7ICD7hDbThk4TOLso3iva
ibUheNMjKcXkvOqwlSSpju0drwn/yvlOocJOpWzsSjBtA87uYcnqAOHqXBL2/+N8
I2S8EjfQOEG48ouDIwHPdztTCUsmTUYg2ZC9bL9n4EzOiRLafL1Wy+TA+435GHwt
2+5pJbAUD0Kn7qFvJzBSvedYYf2UwcUburpgCN2gDxgy4/uPmub7fT7O/033DmIS
Gv3mCDc279rZh6KiVelAxSjWzuboL3apkZ3pzql0iUROEufSK51asq6as0MmYe6R
bW6mJyExLUghfZM+21+FnIQ6GZeb9l3q6JscFmdmAC2uDL6P9ilD5IIRvUMcl14n
gaFssylJMp9vHxXqXaLsGSFmZYToivFCguDNdO/1uz+bnE5FPuz9NPPl31YoH0p2
Du7gB+TxlmYVJ8sXrZSNbrWOdzYDJau38tY1sw3vNgC/atrqlaozM63t5vCrU1wf
Ks3IZzR9JRCR0Jmd6DzzGWV0mPct8vkFL+ceiDpzwvQbOjpwCe7zZphlXL/vzRCl
1BvLFnz++ZlKx3WsynKBGJhtyb85x126C0P9q4UvzOBp5fohhLsOZiFwmDH0nLlg
znpaC/sc8Lxak4HXW6HOVDY6YbQ9wf26m434eHPCXQabelhQXT1XbjWRyfjIob0x
1D8X71OLEfDQH5JfPHkkGpmvyc8oTOG6mLgndgFP9hVj/3715MTQc71m7MMeGjZj
TpAGFGdwPN1tX/HxJuQsCM2zGaD29e5z6NxpqhNFrGZa8rqs3vGANXF5lzITl5vr
XRF+ZUvKVRtfM903TqSvsbRSIKJNVMzHB7fyIWfajOE=
`protect END_PROTECTED
