`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l3gv7XvRBxytT5KHkGFXUqWhLZi8AuIIAWuNus1qJocOHYoNH1uGFJTnAemeIWyu
iz4TBPMlCGNru3NkxSULfd9knzwQrU3Q01+ggHgvgYmjDzhrLBBktTjap/kL20VV
in3FU7sLJRjSFsF9zwfpGYNNenla0FvWKskg7jQQFaBAMhw2t6zxmoMpZxwLFT4x
kFBN52vmecjXCShqNAmFQJpOGXmlZE52viw0/dE7YRnqGIc8/GRENs3n1dYZDGqb
dJSopcp9yenb/XjGluwnpj7NqMxRneVJzxIWRyx7QBWMBPYyl1025U3LwTxuYDsH
Dqk8Uq5c3CjHLfa4TPLlmikKj0rB+I/KbW0D9b9nxHgrE6gOBFaKed2AAy6tD3ln
QYa1/K/nWqp8xNxHLgvXVDyYucN4yLOL3GD7X8a508aaqTqM4GcsKF+SqhFOBIRb
HcgmIkzr/llifo/f+fG8obdeh7rp0Bwe5I6rwmnxX3ZtqCoGDhRJL2loXSL/OSVR
2NK+ctGg3c3a23MQ/0XOfG7UjS3TgMK1eo/LZUbsgkPLu7ARGcpct2CnwCtduJDh
iDK8DiNiRfck24xUEHqsQP8qFdH1HnUP4D2+AObAi7pKmKRMq0WJ6zCHI7WM3gaT
9RkkyRMkzBFU+v6FUyVkrBHk6hmKwZ87qhBSM2nRLi5Wdy3mbWsTBn4eF6K8LsYy
17wzGb4CyIXpo+z20ipwWizUhbHUsci2X4cpoH77wzteXiBeLjrMnjZ8id+wZtln
00huew/yJd6THLy0+ngFtVxx6SoyvT5m8joGZQP7C+ad9YZWOP2fYwfk6sTDs+dr
7+tYdodXMnbUmxtd2RvQxTRd3HZcYZVg51wdcyLQ07CdETbzeMUA3EojeMiQXxcW
yQI4VZhKJTZJC+gO4Udv1xt9nOrZi3Ob7X5VsSSCOhRDSPbkBhOeRFjgTeIQlEMD
90EWmhXJHb3PwzSNeUglmWjYEOK5LaPTzTx3imgPQDKS05ZDvb9COK2svpWluL3i
KOO/N8HvvdNJyQM+H3/NQEHVFMEBSzK0T8pBoFFIH7Up5nUq1ZLXGRs/5Q3QASYG
/uz+6T4gz0pCtVMg48guat7S/081hbyxonRGLwVS2b5lqsBu6nsH1B5npz55qTxJ
lFbibYvPpy4dromRMHpTE+NWUjcXkGO8hgNKvlUxIiAKY4Zz05IWC60eawhphgQ0
u3DgWdQY1eCXGCWgBw8azOTrOsYaS8yQozWO4CcV9qMRhrZpJJgs6P/o5G4hXCLK
+rEDMPw5baesexg3sFfnQoZGlCSeBqHwp1ciw4+11thvTNrEituz2wEyoE57med1
eM1QtuNWEYZy+2Hz9tFM+ySCTu9MDOwv8P5WYZUx5AsJbP/0TVbN7pKB4oTt270w
wPV8w0l1fsb+vI3rjS6kraXaMLfYb+QIyF8pAkoEG5KhABoHYSWpY9cDSkK04HFA
5Gt37fKxAZD06ZMYUYkeiFgzv32Wx54DLVIQko0SXyNheEIOr5CpbGc6zS3VTtGb
wq8jcN2va1WVpFDTUOpRbbA/wSvOg6fyuRHyJmZJobXIFebPaA2ukU1LAgtRKjGn
Qv1mCK1/BUc16Ax4UVmLP/nNl8u5mtdBv10/9S/7rQg5AwmhAYJ3urT3HSdE+bXJ
R9THYUhPLozYEHIghwThUrgDshsL/v0w+py+lmUNx7cT+KRZm9YF2CwSHGAec+7w
M2AMGoJdPatG2gJGWxbNrkGVaaDYbYi1dr033xtYXKAm70//DcCf8xE7QQdJsJMD
WaOPdWA/DQvc8XVPPHf+9yojFi3o1qP3MG1nAN8bcJtoFil9wU/dGqgvxV1DpReG
pzbUBmg6CMiXgs8X7bemMP3JMzCaktOo1gSrwREkV6LEQr8ekEirKUiF/48FhZRT
TO/Oz3JgpTRpHx+eogu5yRr546JcA4VQz0UqYyoVTpPUCJvG/shgh7FnE6Oyqaep
W8E3wOp4JKSL64226P7EGqj4gNC1zXyu8YUTDbS+t9T//8IuqD7VW2SprABSF1ZA
9qxFX6ZCUiAxjYGaERfqSLB1JV8d/dhY5INcVFllulL74a7gRKFJs7AK1VlP/YBO
TXDkQz3aVZ1CUwQfFM7dDTtruyi6neT4d/u3BOSlRD0IyNFCw+nmN1EnlKOqFe0S
eViwOlSpCzVj/ZP2mfNWG1tputnJDq07uaho7T9KrvsfZ+gyRMhn5QH2yDdfzIGT
fp7hxWKF4ZRGDfqHvqt0Q57nvUrBsfERcdaPjwLato8KBREeXeoqRp1GuOtgclLd
hmxkEZCfdIn7v4bMWKjSYBkNwJr3WKQIjPdp51X6LphJKweSUvdL8agnPrArPw6p
gKzxA4mFJId407GkaTmzFFzcIKw9Eb0j5Mn25k/qcuRb0Hch3t23QkMJMXbdd+Jk
Upl0SiSGhyPAFAZvCgWFP+jHRenTcJMvQBmW1PA028URtFyyKTWIISL/V9YcG0n/
gYpCaEIirqNNYXXasjW4xdSWK/hoNNoHwGw/ACdYVzgkRxyKTj7qn+QlWZi7gIBE
+WJLzQAEdPbhmcPRkr5a36yESd2Wo+pVDn5LxOZk+tEOGsQTTNbDKi4tl0szwZhy
3OAlYjnmZklWWvvHHPyeji5NH11la3EhHMcS70IDaWxDsgi4TbExAbR0+wQWeiR5
AflUawNlzpJ4Qs9hhSNOeQj8TfkVvuxGV0aibceYZnQp3NtGWSAXiA7/lbLOMhDN
Qk/Kn4I75B6nvp6oGGSOL5zIOOP8d3VRLSZawumS3C4yZ5cqMsq9JeoF6C75b2vc
sd8gGu5/t4kk1nTiZvnL+y186V3DsdHyJ5xaFhOXnPtA7cGfId/oIr+xy3PAwGv2
MRWLamL1cM785+JT1fmV4kF0aKNYUxh51KIhIvco2VATWOKE1rh9mOFydOTRTdJT
/lQBKP5AUgZOuctF5MmNMLrln9pr1NpwGdcmppBGGX/4Ida0hqRJjfeysApsXaF7
JUc5Yg2EJn4yWLRlmTK/5hDzwxHbeXfbjCk8wB37upV9jWOZWiFsbEPSOVFWrN+D
4+zGGOiptr3EAxP7XP/hpOB1IEBsgTdL48Ux5SGdTljV2j5gfjtAaOBg0lxPYjtR
+cgl8fuKOH+lw26dL1KyttJLxQoH5fvdA4IXvD7B53nhb93MGvO/JCA5kEtdWWQx
N3ABVzBQQUerxJd1yEfdcZ5VPu42Crjk0C06f75+XgctLnNZ2O6lNjB4p52QBwGD
YBt8M4KcY8ur1KTjBdr8E2ILnB5D7DjctqBz3uAOo3vSx9QtzFFYxmwiZeuJpcq4
+bbXAHRjbKzEzoUROK8cmxFU2bHU3DCFyStHga2YcQfQGm5h9oQEsBx/M5Omzu/+
DKGyu+ClKx+nKaKAcmdTv1B+iUqzW2myzdj8TqvY782DQCw0l3cAnWaNJaiBS6j1
ZS6vkQTJIup2hX45ltPSe0oibnR49kKFvymdGedWRBvLrAVPLMTwkyQxH5yDZlJz
CupsNEXmVYtOvnXFmc1ftI+0eXXofLaLv4PDr3XnrSnNiKpL33SiFSiCmEVol5Pa
mY76iCYyMZe1CeI8OAZkapnlDCZfBP39H0I8tM04hWk7PXF5FwVZLO9Do87JussW
mBQMKOw2+Aw3+aYdt5VvsAajHtwHCTe209qdclUZINR+RE7b5dWLi4TH0nqBXZzr
Zel8kRnWw7MzzDEAqaToPm2PG2+jDvNEtAfFpOMFXYoAimQtPLZ3bsboxRTCmnt6
0DOZHbDrQePc9gbn8XiREx5ic1hJuE7cm59/CDfmi26OR72pQvwlvWS9IALK6Kiz
tKDCfxAeH7P4muifJp31Jbh+c9bnapZ5fl19RkeaMJ0jk+djz+41pSictuYOLmKo
Zia4OK/LO05lWAtf3zSVas2nBs1fhEH2rdJZs8+Rcnj7LF06uLinYEYiddRnUJwk
pvnbDpc6LRLrJY4m5rs6F8yAnLkMz3glVxGhFRr1x5yTZyxetGJiEEm6bZzCcWmg
41qKqlk4nbWCm+ccmoeFIIwGN9ZD3PU3Q+k48XYw3uYRWrRrbhyOYuYFgp8JqPaN
4/blaHcQ0CxsvCr58/bx3uqiwz4gFCVB4dIyWPs5Kg1FbsD/F0R6h6IeMfI9PZ4Z
pIdEn6OTG4r7OMXgNVC9A2nnA3oULzZlEyfnM77zvmYi0tEJ6s4IxE1D/j8rWo+b
B0zmNa7Ho/lgAw1lgjoO+vg0sJ1ltLgtPO05/cEAr2hJ3o2Nvku1B8SPAiujhKHx
sGy+RORRg7gjsdy5g4uHB8LCNfbQ2/xzk0yg65dvHIUgNYGm4f5EY/pLEVPLbZoK
tNuAWGs8AA5BAPxWzRaFVDvDCWMbMxrKFr1p9KuhOn0lEJFW/8NbNdmAZaaARUAy
rLpeSXGKeawTlsED+UKSn6BuHlHZemgnF9PWUe9AxWGBzn4nQgBydf8+EZG0VLUS
2cA+1wHZ3HSJdFcqXxbuu1HqxYvm1JszN6w4YqdU8qMZYtxFp88bVQHdldmzktUk
LO16bT0WRoNRtb5udVIpcTiBSG6sH2tbB0PkXCxDjfx13p1QALlF6QaNmUR0Z8na
nSrW2sL5ANUdtaLKTSI4vyhm2tLBdXiHPkSED81JnFqAqXeIGPULNGZljdrTMzra
cyZJGRGBSSeNF6p3pKmBE4YGuk4tbZj3cfNDXwVl1NLQvve/vOoBm+BizVGg8AzV
gjr4+xYW29Jg89DcDqzE/v6ko17Y+4rCLpLwEVcX2I1idaahNvSpvRe8BQLyRImC
hp/n3kh0ciVayrOpVDwq9G3vL/nOXkwqUTAWAGXfqKeiV42+MYEQOpUx6ED98LIv
6UKK4y9c3ar5UcHb1rwa7L2stE1dVwf4JlYPlE305jo49zuTPDbM//mmPmWYacAi
ocOYpKKPqSwdy22oUwuVXxX5Fx5nlVQdzcUscYfUc0qFho26+btLbmdtTSgRn30C
olSAu4SM3D3zpETU/nvIVIoYffIbpsKYsW1ryLkYiGzwOexNELZy/w9f6X7rYZ0L
9lnWxxoAcHNVN4fLjJb0nYAya8fZdsrUmNKRP4Bx241k1hUnc1HoVPEr8bYDY2hH
HHZsQazjqSVcrshdT7ClOfTGjABCmX+RvMBEaW/YOoDsDZo6+LWZovad3PdfIVNm
i0TXM5akjv8TjLrL1De1DoFU1ls5tKUqnNcK2Q2UnY1su8tzmzZzPSUwZ9RGZe5R
gU5xJB0gPHwUqDE96E2d7u6NP2HbWf8KTqzHwiwn0+33aST2dwWwfVbnNFBYvhGA
1lLvVHOz2sPMZXMCs2x3HfEP5yMQ+gaFkAVMvmFzc5N+Af4/qAnucBII5r9Tw3co
74t9oW7o3JSFY3CGhz5R9MLMpBeCOAFnXlsn+vlQhm5UF3yJJvhod9e/bEHiHLzy
0i9XzwAEin8Epsj10CFvI76q2oN4ClVpaDij/GLi9hImlhn5VfgHcAd47V3RFCGT
Mc1LgDbE2E2UkfNIjPAbCI0DTw1kbOWkA7pYnqRxBP39C+3u+sXALcL3RnBgSOop
GBJu92saCwITIeuqo0K5U3hc6adLxRNNgp4/fKhVKFk//a6rEbuCajROTsklBV53
1by+u5gLelTf6mKYAHTIxJMie+3qIJCc9I9LJIi3XcRBr7D5RXleJ+40jQUxXpHP
MG1XDz5MYkQXSio0t0FCXMl4GfkJrbLGGeTzN+IzrBIMaNu2sgqkSGmiJTq9unlV
itwMFpAtjwfWdhNkaKPM3iqx7LzMVTE7nTx9Z8F7ej8AyxKhTGNr0aJTnY6iyo1q
TTp4I+2YXXKvYr7HYyU0K8Mrf8O+4XKnRXjR+EXcb1b8BlbWf5BwavaoEhCK7VpT
VgwacHS0U7bYUwXieXWveIFMPFFIFTxaRQfj3AG2Hx0Zp2avYTTb3zAUeYmwqUTN
IYAYMnwP/vs1tmAi0Bo7C3b7zIdVAA2IV+2Fc1ljjtfe8sZrRDuDOcZhilYvuNxV
A2nIbXoguqm17C/zCfCsj+FARcTzi0wS5ke61Xg60Ivf+02I7BJED3mgwes1Xj9A
Ss8rp6hAqX+9caGXEEdpNiTGwexXVs/tKchOOsPeugKzKQkBImUIcpQoTvBfi+cX
W5t0kz1G4OY2YJ3d2bknrne/P0gvgk7IdAnwxcuPahKixLOY5UTlwE8Av0V4e0OG
LsHj7rrhv81e1S9lEbN0wznnx6zsaBo0Wp3On7TKe4OnaqC+nOAq+L5sA8js2Rwt
GMNJVpP23O4LKCRzkjD5CgECVkxEeKY6837MbCJWF6/qkTnDR7QQOEmfmKoNBdrs
5TiMHvpVHf/i+eISwrhOzbhoPKefXzWgXLxCuAm3DiKopRAoui5A/3QD4dQfvGJ6
bgCXSMewPg+/sJAJ069HzrJWsOyjBzdGMq9FOPZFH9jmSAy5w/1VZx7q320sVvHZ
HJdbmwpJ1LMeZDqVO9km0BrnL8mv70aFU7Ds9AUYGb5H8vle9KP5S0fxLPsz8ojo
Q52dHQ/iQNb3SGuNWSfvsLAim0S3WRny2a0rWkTcB4eyhXhIdiRRDKNYMVH3H1N5
whbvZXQ2od6dA2zIlCNEozL8PUaayjiaiavao40Gkd7InVsdJQ6C0VCZKSZ8MqUq
93Rx5/rdLmSq2FvO37KEBwjvhJ/ZHAss8oO0TeZEr7X8UNQtd4wOjxTFNju+CHpa
m/Z/L49EVqEANwf/Wi9B2epkOH1MePy/d25CzH22LFaC+kuiYZQSeFhvb6YVUYr5
eyTiVONh3csakj+yif8U57QQaYvhqtWbJMjzYBv/Rk9s5dJ77BRRynEg01IPJxs5
xkoxhaZnB1NV+jq+1XH3PV+cqX1orhXMVwZaKCK8pqfNJt1q6VAE/BQqyWJXABkw
LLlci59W033aoahYdG8ZlRZc2ThBeUt8jWAL7qt6ZWOER1JOdKEqcP63/OxvIytz
hqL5As3beiQuQ3QGslfyYLVwsDdgQ4/tUdWJsCHyT14Pi9InamcKZr0GmjiPeYuy
EOxnxmQD5PFLWUoF7oWcBMaaFr7MkzodYjMH3KYkO4iRorl7rAWeeqQPt3Fj3xiE
XggVs50PpVal4vicOptVHeKwlcJXqzsqB9I+59jZYFCho3WyBfn53mJHKQhOgfva
pQ8R5ypDzLCbIIr+AiEpYwt3nXpMHcqxXatQmpcCORq282sIOJkoCSt9IS1xPvSf
hPlAeOBEXGzntPv9Ff6KdiR3WF4Z2ydBnidI2Jh5U8ZpD9iNgV60vxBJYGLOn3ls
EfqT7Qafw4u4KaoXy4UrWDNcD3innlYW09gpJAJX8PF/Oo3ut5zCEdD7+MExSI1k
QH1bnUl7KQB5cJwMCQsRxdO7h+vftZOZRETqd4EGzu6YcaYwCvdFydUJlyLEOFNv
2v4i6KiC+6P5KbrZo3ffscaQ8xcdiepPVV8CyCvPYEErIUYOti6ZIDT0lqdcEbQi
IKUvWvsysl9Bryv9KdWwqPlpLsmquB/W7RUUsPWtji7ZhxRbWknJglzyb1YHGViV
FBOoDjqkSQvf9v9Fc6VRaWWBBMFejOUEw1GD6c01V8utlvU+r+GweuZKIVsj4zvV
mXVESQFi9TBAbVkSnzlAnmTwxT2d53yHkgQ3C13UOz8CSFvIJXsfkyoRqN26kame
exTm9CGifBX3MRXnMAz9UGAXyE71kURTNQFYGYcfrMYl8yAppr1oI0SEptdYxBfg
/2uT5A8X+e6uxv7UMBa6+bj1rwIR+TD4JdENjXKqbPZB2GnqXrscnWIu5RAedXMl
y/BroG69AqcjDSzF/qCalalYJ1/aRzAJdkIn1z254REGfkupN2XRjm+IhjWUzqsg
O0ZXbqV7bol+NbBp+6nDSjNP9bxrM94M/9sNBT06LpjvamqYcO4kbDtKg+VFfQOC
NnEjqNuU55Tah1ZiHGujtZ9UIeQH1HjrdDsPxLlVwaOZKc5wgpw2EsO0aGuqx5w5
eqoi6gv+hlcmv1sodiZTQXDLnWrDxTNfIcAaKT+CHx1/2guW73LMg7OIAdJK9ns6
kc0UWyPTNGN1igzZLrbCwmQxwaZRMBB/HHyqEIu0wRpmu0qZGWh0qdbNWeN5yX8k
Ro8hhd/5qfs88FI74bpIVpC0pLWuW7TBylD4TT6QXogBJtRpjZ5jofH3cAv1ILcs
83oo45qdT8x8cUmZT26GpWIwIKwyn4nEdmbXrcZsM9tJqaFDwEEbz+nUsAoAuoNn
R9M24dY17oV6DwFbob1CTuC6fAmMif9CNSyblD0L05B8wghxFIs2ucC1GNankful
Y4sIBMZKor2wNZd6V7r3cvdLx0pFQoFvkZx6YZUuWYOKT/v3HzLVo9qN8SDa90np
nn3jVON3PKUrW38BfD2yPIJ5vLB5MFvdF+AaMvakCEOmXwR+7yWRIqTcqT7fWCx7
7bRAofSSYMIBqMZyNZ68GEvnGMyRFUVbfPraLtRtKsyUnhFIkGKMPhegKMIXQvkX
cWzv4IAxrc8zevrsR7oKMD8AkdIZHYjXc7Rm0nCXtOAg3MLTXm1OE6Ha4JaJy2cH
BV/cf44JW+6dRNwMgCB66QE4jWeDvf3wx6N1YUFK9bhxP52TKBVriObYr9HCbvur
g859hyJMoE3cF+64ls1qRLXghkC1pMlonafRwJM0MeOcFb+u6LDispVdLlfIF3qy
AOLTb9KTPHPEYpn9KxFVvj71/9jeLth+brXaOY4AIWrXcQWN0VPAkbGh4sW/46Up
3CR1RSulR65zAO8WTFWrTbAQFi1UArAtXIt+dJYf/rvj5lgvo+Xr3A3gBwbT4kik
BK0XE0Vd6KA5pVl35udeezQX7OzBEUj3epv9M5SYYz8M4Uupf9FOpdsojz5WJJ4p
abk/f0uaMY5UP81IgKn7tZlMSRlG+FTAf+ZAoDV/6b8jYgkVIfUtEk94QAeLnFtL
du8cj9QyfOJ1hdMoqijFKuWEJBEIKmNf8RV7Pg2q7UmrKxXY03jXnzoVNVYrfT0I
jHgI7OcFyhgqklNarGgtK15t7g08zOVLtgiQoWgPB8l5HUsmJCCkG9ruDSP0gw2p
GKmgn3DTh/89ovpTCHcFMo+Q73e+QpCcf/vm9+OsyumyAqxn7lBlwjJfX1n/wO8v
iXNW+INAWBQaGEFKtvXn0JrvCw9Juo1zOC8GhXmIMlx/4e4uSqnCa2I5F7yyZ+zs
Ltvwa5PwOgNlyrwMph+h3BcWvmySIWfCf48xi9/7rhBAcO9ISCXtwFmoB+K/4AbR
rwNyS5bKTAmqmnyBxM+8TdLGUIMIIcdVes7nDnMYxYZPqxGje07Ad7F2mC3wyes2
Qgtlfml8P3exC2HgqSA+WA065+LExHZ4a9hJdiIjTBTBrbdM8x8Md0B3uzIZx0sG
JgwVy1gm8hYyYboFNfRvwMs492G7TSOVcYgdcWwpUoCYJdOiXYbAstjM21SBjuCw
MEKyYPoWCk1srql+IaTYW2ZLTvqTmoxCyhy+Nk302c7W/JK4uc5z0HwCrftzgNQd
NdlPEfDZOpqUmilPKSMNENMat2qsNrjKUkylACFWYgbGIrnRUumKgOimDPkKObzk
bnqQmSnY1jaK5Ds6bWnp6B20OexN6NK4jQSjrGOMIPCYHT/7DNBZT2SLTgGaP0Zr
iTpPOx5ym47j5/v9/sROgw6OIKCPOHNAqte5BpQgtnWdEBEtww8GFxB/5/Fon7LK
joDXQd1peuHBVOtXSZPPn71MDQkJlCSwAgJO1eLTTEEZT6LkU+g3HAlgTDmgP6/Q
6rEPw43+U/uYIFE6aVgfefbhgiR9+uN4vBvRejDz+5hLdblwrHfuhiiRNPI9A2Ii
zAyTNXjJhWwbQIxDNFFf350BhGwN2N0d0NdiP+ReGjMst75N8+w2tv53MMpCWwRK
UUKnLYvAWaI1IrfhS9qE/Xu7AuwcxEshEe8t69hkVmPJzeSZNQ5LYI69ytphaReI
mHh6dYb4WM77ToxU6hh0BathUEyZ4R4j08WCF7TG7p0lg5eoUFiNEhG89+Vp9nBB
FVlUy4DDlI3IRQXABMm5+wlu+DiDPuRLM1nFDGp42MPojwLPePJJ1SKxpXwj8DIn
e9UDGtgUnlhz/NHmGlGzHRaj0XMu3fruxkGwSrJqmbzgxf5qiEPKH3ia/4T05efG
uvzOeeYn5odUD6gOCTKcOaTuK5SkpQJ3k0iwohuVOtokZZF/Lyji0CjclrAqVR9W
wCbTHvtu996f1oPDU6Hy8uo83+5glcJSYmHJAGcCaGx7ro9bNpRw00sTR5FRS0G/
Z3IXvpxcPs9mXSooDyM3XqBVjVsttGgG1iJa/xe1wsBtBTUeIbs1s+H971ERYFpG
wVgC0lB0Z6kONTkjS35ClNNDmKx8Qe43aUlCADm9PsYWGnRQVaqCPz2eDiGwoL7U
1hSts3EjFa/bKkFM+d0UEaq0f1dYMhaJH+LXaH/GgRm+LAjdIjMPN6avquT7553S
Sff7Sqe1siKHayjX9ijKmyTaLxGHKminugiGo0rFWYuaaPIgVR9zThdptnwLUh2I
+/liZtvlHFLu8PnAAtPaPEYVQk91FiwjBJiqB2iuYCyjar2Htwe9x81hB2vrqANQ
szo0xHIaeKn8vFGTKB0tVkWFiGCLMiwcUsN3FxeICNrapRNxaWAZybgVFFRbszOn
uepFflPv9PbNwL86pLEa9HffDh09Y891Vu/NEQ6eqKFFW55DaKq94GLzX2aC5u/3
h0vfjkHRpYXppNO+rQCgrLMtf1P5YWRqDUMVnyljl6bzm8Z5oFN5qGBqEdj6LiIQ
LrN/6jgZ9LFifpIKhoQmwy6EjXFzyJuhr8DNX2m9U8JSfApHL87lakHNPiuMWZ0S
eHBLVcR4ultWJ+l3jjj5pOb/bH/PiWuLP8IEsvldBRt5hwi4lYpGsTUVcrdFgFsf
jBwYwh+3O39cif/3ki19Gcm6SVOiWGNoCLaVqSwCd2RepRG87fjSUBRu2ggHWhHH
ASsy9kHX744WL0xuYaLAfqo+NErYmPM8h6ujrMv+qBlxy3l0zjXwQBkTpnBna9sB
qUaFxBvxqNtRqTORJlJdYcRqFcA1xxr+8vsQSauvA4IDVNTqc+z8kyifhL8tsF7t
2uDG9eML6iNE0JWXWvJ/gfe/NC7fTb7VpZacPsbWOf4RibVpuTBxxNcfcZmMhPwC
Km42n/BroAmdUrjjy1+VNr6A5XGjmYKHZphaJ7pe8NCs3yK22SD+0AlyZFiv8WaC
NR+zQJzxKqiOG2MFbYoNgBnSdeA2Lb3L126cqlGw0tnycFirR3tdTH3mQmtsqDzB
mqpqMw8cd7pn/TLCuNKfbaySxN1HdK68XIBHOEtZi1vaUdyj67MMjHSkJpTAXCGX
W5mxz3kad92HRieXa+cvWknBTQn4IGl3yxWYQAqAh0Yt7VJMmz8lZ9S553TsyBr1
PHMvRhTDvMgk5kRz48pnnF5vyxWxnpfdcKF1/E9UrozOpqFL8PjXLOI8gFC1deyl
uQPbTnTbgLNdeXEaSzUNYsLg5jwg/qAtWkcpC6lBRkgw3ZF1vbdYBRj2WOMdDBKk
9tvXcbrGEFES9YMB/JVuSVnCEayG1uKIqLum6j8Rk62/+XlZv8x8MZX564rfWtqy
/uWZTF96nsHvjfk7AUU0U7q9+ZE73q/91KwdaGexu/vIar12OUv/tkaH5gDDBLF5
NrqrCGr+C+8EKvKzu8anvCqtrLWKzCjvmVY/KAGPUvQBSJXKGgocipsT6cnJwD4y
CP1l+AcgwgObDvE7JH4goa0oHA25Dxgamgfw+y9RcxEnaqp+TY5bGqdtPyIe61td
kkHP+70XVdxAUHsqfpFRnLVzl3nANDnVya85Cz9TGMeldxqsU1M8MjAE1uQM36V2
DJO5Z0YjOkg6Ai7PYbch0G2Pp51wDcVDTyMLY+s6tWrk10i/wZps6HbhjaTd4QOX
OTqboROMr9wNb5uuYquNlNiWe3tmmut+LFQVEL0ZHIJcn5CQFeI4OFbexIvUUOTa
kXYHAKVxqQTbZcoc0NpmqmXYPIBAgtHXnC1ThK5BowpSEwxIyaXauky8uhHmN3cW
n4XT9xbbYzrVa/FemIwp77TeGUxM4DtFgMOwfJbWioYffQOqEaAElpj/XLwyxZVJ
WrYyer7F3pORZ+qcJ/M3V3yVs+1gk72E7pTDo4BOTQL5UUemY3Km5g0j23v1UcB8
28bCcHq2vNPNZ/DM7bEfOS/7pIrCYPo714Qr1PIHVzJqxwSxeGs5HwKIX5lPU+t+
6irXFyT0OZVUW8d+lRR50KH5n2ZCuJJsWMIRqASfMNAiAOr0vqoyZKK+mSAMlLxK
8G1wIyH6Qif+ayVCr3l8MoT4rItmf4qjhbNAAh0LLveyCteIZezXuX9FFPCoV0Xr
pVX65aczRTSUYKCoy4DkT3hb9GFv1xkO270123bW7cNx09H/iDtEQRmWmbYBYOPD
eyAxGkYMMqqu1vrYfQ5n5O5IgUCv9FCYcJ8FDmdJ37dC63E1w3y5XJ8oTpZTDKjT
5+9rcZ7hrfRwc38PuGGl6XVvn7eWuYnTzY4SE73Dl70wJZB/3jlx2bGXPr5FAoqW
GO2/pE/SLut2HduJImpH8SOZbZXdMMigaZstoogaVIW2xdqb/1Kd37DFMRStzTMk
jeuogGGazlTL0g0gFhEpvPzSRfNlji9oNvEkpK2umEm8/UjXJm8ra701EgAsf7BE
3Onm0Hgcu4ut02q2mTvMmOMf7UbVzzWcd3Ghz5QZiRjDrFi6rAT7YnBWduHz33W9
Cz7JroMtZ0TjtOKGZJcFiDLSW035f0bABBwxi+PLOpBHMUh631r9YeVLTMP61CKe
1POyc06ZRPZDQeMBE74Ory7WuLR6cAyAW4kN0Hbf9T7QQESiEHvtd4vLBCQQtd9I
jVOWaN/nCV6z8r5xyhtvdj4lB61JPGRjYtLZ+Fd+TZAIYcf8Yq3i8pJJdPIF6d0z
oBz3KF/WKXV4XwpLJ0vzTpUvm7oW+kr21BRPvenxCZYttVDv7qgsK04vRhtljbkH
2WfAlifgInh8Aw2IqoJbl4Dht60nslRC/Xs5FtXoDslBBtYjgAy4HW9Hq3XMD0Jz
mp+vGr8NDYoy+cY9VY3xz5UV5Yw6hBH8EI0XHAoe1CIlXYkaLfqf5EI2w8rv49Su
EcyQUjJj7U/igJ7OW5xsTese3gsJmMROuKkLCImq7mx7An2Tjn84rw7hw7Of1pl6
2wnqhl8NanQOUb2Toy0Xpyf5l8EW1bbG7b/IntK1X1lGjkP/GpWlWKbxdPXgn+Uo
zUnTkTqp+i2+n0bhuFqa2FHvQ4I795V/uQtKMMYrtG3ePMDULtDHJ44cFLQdTnph
S23zSR5qUpQtNNaCzmBkX389n3pQcQ6oiHtxICP27MdhlvBE3jdXVdMjTCqOq8Xn
89VjUPER1jWgAs8JCUNjVSF1hAUmw7N0PSCM76y68heSG+lKPCGEhvFB2GmOwObL
7tkcE7xmEBMwCi6jHSJpgo3RpQPscOQlyifdWSH/6ik1SsuIUZ7SR/aqtiv2lfFQ
O6LTIsVVk/KhC8zT1hnU34+EGV2qv9SdfEqXwnS1Rej6qOfXQE04+rc6jBCuPw0m
5xUipCzSOUYwyMFnnA4dKwJ2bR3GBdUubml9sUcLg5dZEtdirnqBwGeiEWAtGrst
ue61SsAiqF7jFNqFwenSvp44yPEEoL1tj+uG1NhAtO4wz6Ew7DD/hO6TJmczP8Hu
yJN6iFQM3ULqdjLYG1p9IgWZoG/5lZg6uXLriCG4iCOQ9CSfGxlDo2aaIFRj7/vy
k45qRhJcCer1SqettyiXo708TNJ0zq6fjIaMeXiDSWQbFAb3Do7MDaSWmlUsKeQv
nRUiCFKgMQlvy9i1k8T5S1ZGC5CijYfd0dNLJuptHCjshos5WfnWYfIXqpuAhW6V
FYRwWmYpfubGvCOHIwWquT2M1YA6QWOED/nd2P6PV2zfBdBc7fXzYNXuvSdfhiU7
gu/65js/k+MVH5DmoNyx/fkWPDVgaSMp4sjqp9fNUGYfoumMm7GqNEXB5TyNzITj
/+VMrsJDhkWtP/Cigitxtznc2ucT6wwO+eK1B9ROLuKhbylTLhkq1xUDQvItSpgX
a6HQ+Ziur/Ff3W2nMvOODYKwDo1MpJh/xX1tiHhoX2lu2sbFQI8uOZdEzCR6h5r+
o1RHBAQFYUCLgLAeXgwnZaHf7We+NTYMEs6vZBP/pUmpTU/vftq/NrajJiRAJGXb
QpDUlEq5kBMS/DBD4Fyf4TYJHxQb94Dwf8XXiepfJTdAjy8dBsspE/cAwaJKDrhh
iaQcezpxHzz0JPGFn4x2TBBU5Sy0+FoY5LkBNqh2BMWZs8fbJMRfH9EmcHHejpxR
vR/9GwwA/GE2xuEIe4lvBuQa/UyRd++lnPcrVQyaCqWVS2bGHySEtxWbM0ewZRFS
LD5oxJG0p24CNfoJMaZD6fA/rT2USkyg4E/lI5506cXCGUt0vyNKTcH+kBH1Yypv
p6bYm4FNub0UynU2e7AFxaQsdKmd3fL6L48FkWV1KYmCpA9F62OEWLBnSBOC01tJ
dcRcmoF18J8MHMrGp7Orw2OqCDgUIlstDZgbMA1LGu9jLZhj+/YwlD09Jr9SJiWT
rZAjqXN/+H8naDa+RfdOfn9KrRX42oydcMbgrjfKh3ZAq0iacYzxuaqjADL7tiZ8
B5Tuqe5xgHsMKlsw+SzfRtw/F6TPADSYX+PoEYWRM4suIDZ/LOHH8a0hd/8050wy
Z2jaDWDFizVuAu6Ibf1K59Y+nmlT5LwnWfwBQMwq2Fhs+q2cYvCg4Hihh/aj7czA
AYW/OfUOWDYO0ArmMIrI1t2O2ojyMHOlIOV5aaRDPlAxjpqIGzicncQIXG1oC+Gt
gHOjOULdpTO5OskPXunBEo7AO46yMBhFvwcrA8lQB38+7lKHgnaloJuvGNO1OVbj
u9lt6LuTdGpee0hpBB2q/vQtNPtF5smFLJPJ/pmvql/sz6QSuPSTLjk7c0FN4k3L
FwPCNWIel49Tdt2XqNIFZdrbQW41iOQf0NAex4zRfI8pPl1H9ZO50O9HzTRrEhkZ
mA6caysyCUiwJNagkABUpYT6oqJPI2quuWzN0UM7T/HfkHPRRLJCRFGb2Tun+Wg/
wdk/2TL6/XCOwZl1UJN5cFOyJG8WOE8KE0xf8qru508CU8WY9zp2yWqM1PXdpOyC
Lqtrac30bTuq0QXY+lWIAvZreYksVKKOJ+tihEg0ZO9u9blm/AsWTQRH8AzqrL7V
ddbA57IIGje8UEwmn3XzHechUZDt3hBzLe8JfN22uwHld2gJonn1YgCeBRZjpjDt
1yYJ7XYpfWZK+qywIQoFTBq1+qJAsxneD44lwCbYg3Yj9MRqE8sb0F3sCPpoQLNV
RcqGM0f3NPbUiTo6lCH0MJlVMOUkO97/AQN/f4Dvvv+f186mKoJfC57JiI52QXKs
DX9/m4R8Kbub5OHiEkntX8urdS6ET6IYhpk+vhJH8tsaoStJrlWIcDCHpRwWWm40
MZDF8tPx/i53ADX/YcCujYJzyTPamoYdhRfaMOBEf7U1azLq1MMl5FsBOgp0sFPM
RUgfv04kxTDC+LecxcEHAaLIL1Jqrb/3mTDRzNpv6UhODP2xxh6a2FemKRLg3IZL
Fck/MXxY9CGQqwUCNLShBkZV3bA9cjt9Q2QTWl06AZj9ZPavpMvafMmFzprM07BN
jIVHHwgND7CWp8k7WZl7JxMKxZTly56YlDyjWwD2QTdSQNeGjBs56FNsddYTSqNT
JibqX8WugX0U6djYmjdkCf1taOPiNxKPIcM5XHXHI4DDyzhCumQjPOFmy1svUyK7
VbsTHieV5+OwZ9ZIsgH6HkOi6vPA2uZ6lo5Q2FEsTEzvl3cyux5GGfPlWBTyV8vz
u7V4DcKKKLwtD0RaLp/2+t+2MW1cD6tqRoP0vabVFtYq0k376kL4FCMCfw0aiQoB
7DdfenTfBhoJRdL54D/kTVWaMby8VOl6wpeAL56dTK6v2iI//ESEobh5GgwKZuAb
EMgdOw2GwhLdApOFOOA024oQcJ1xtFONiVDOXzD86VhU3ANfXollAALja5jfGUeq
1NQZZdmkopCNuRlGK0fucmig6FOvhMPm5CJqJMBJXgreTQPslp9tTuf7YnhnZQ95
pup2dqNP1l8hGRVw9UH00hHokhZ5s2fQPJytReFdiAlycAe6xI/NF7UhES+0fxx/
s6TchjW5FWeDjqK0ZbuG/GJuqQ9M6Eh0tor7f4qcGoSmD7VtYjFThtSkUjVzNkdj
+joZtTJtwfiFAHoUECUN+V7FxZIJgXNSVRNwFULKCnKPsQ4ZuuYkx4IAHjtcW5cK
uj89Tw7tPQ2xb6wa6SnRNONFp8M+XB24QRQdr9AZAnh9JOX464FuuxGka08ec135
2F6Bre6oSvEPEjEO8mBMGpfwLd0tTNemmPVt7Fmwr/GNNem/Xsuy6M9FLnpCkfhJ
NJA5l1mvDCx4HIxwkOhscI0pmwa5Wgf2Hxtrf284e22hYlBE8x3gKIeZn2RIwfu3
lxcgdp963GFhUsgy/o0tl9Gg54jxuzoAWBoJ6v/PE+0agKzNNUuyVW9Pjz92hmj1
IcayJCTxnmGpCZKHu4Vklz9dSgKiDQFfkQVpOXHl3iEhYduDDFMQd51Si+Rv2EnL
lCWSxdEdXvffe+wti/zBYeFBtfC0bcTWGaSaSayf0SJTQ/HD+6LYjeI1nSiKtLxL
yWTjgi4RIBDHSsy8tpy47LfeBFu4WpBy17qJ5as1Leg4vm/gS+g0wZLaIyZc3f3n
YAPdEd5capTV2ZQUhFZVfzEJe9nUE/a5dhAS/jPw8p4I/59rNPqFKZDEIO8nSWGx
9rwBx4jQLzkKwBdTFY95Y7vPtSRT4CpelyHvlX3bZzTMXVipxWp7NhycQIZH3aWK
xvVM7LWdQi3cWhOtodRJvI3MO8sLgzEuc5qypwoMSLyzf8DuikpmjHDOEmRBV0Zr
rMTZBIKWC99Hg8TOdDDRAEWshsqlxQ8zj41JGth2rMR1l02L2RIGFGAenbfw6jGE
2SEvtSNrk4eGGiIpEnOpKsGoG+bN5Jfp8XZqV+0HD5igrf0eyoow1R1TbHcZdQiW
qGGWAv2HBkIRVZDyPwnEUwB6VaC3Vwg9PGbbI6aksGNPQ3DH5f3Atdq66uv98gLX
BUKaLBinVvcTqF0MDtTxycZf8fmeexXUZYXYzfxlACXcEUXoVndmQjlmewRfagWM
Qb8xZ3Ce+2ssy7aVPgGbN3fKsefEyyoDPXOTdorz4JgtHT+Q/38suNY4TAVw/j7C
01Ah3uX+jBD3b+slFnmrBxUWz1pQilauGZEVBxX0E9/L0vUJY35OVXLVBtBSKURs
PrB9r9fJG0V77qstcf0WVIvo9gG4DvfFFhd9UOuX9JXfbslvvEBZ3IkaMPGBhPiX
+8KU2X2LIn2Y0YNksK4U5XTZLN7ainnesKzgJ/fjbVdq0c1jwtE1XgGHDVCrZMXK
bLeC5UpBWZgbCB5IYJZSxvrn1xSfwcW4Ez+P0DISOwXnB5lDYkdLUFq1hOFseH+p
QIecnHYvE/Qvqhb4mVMgV+xYk0ZqHHWgAR2bQc0xk9+U3IfXhsPvdr7Xb2QGkMS9
mOqCVY3Yz9acRrhhmz/uZGiqYTOCyWsD2aUV0EnQjPIM3N8yegkj97sEaUz3vh1V
0LJAVGtLErJIOPZzh5WAUwuvqWh5hJ180wv2zotOPghG1ESJnYRbcNXIVzllKW/+
lPUrmwMBBZI2Jr4ivmkzByk7WAfJm3t4JF0Rd3Z4LJ5tyRbJ8aHIQdPJNjKjqmfQ
IiCrmdMsGwqZmxqVEoacIvcPEPLTw3ptqcc62aRk98KNO3/lmYYkuRZ8gy8DOFa2
q3xWJorfq7QyDVpZunNV1MwGu7FyigzXDQfj7EKUfTQMmI8w+QGB78V03+goRk8/
YLDUJlk6z2yLOn+ejZIHUpGzJJGM3Nj2FpRfXSWJEF9PHHkW8cZZxwXVU8BHeJf+
Lce9wMOb6U6bo3t32guox5iEjDMq7VItF+pY0LTiiZqixPElrKwSSkJAjx8lagzS
Bw509Mb18y7yjKMaqb+fqEncNdn4xqWryfyc4/iBag9TukL0V2WE/z233IHk/Loh
ymiTAfe3YNicV8T8kSGKXAlpBMzmWEA/9cE2ng9hzvVx8L5AnZdHwxgIaQ1axxk2
CpizQtkI7wEqmakPGtOnPVhr69SBtqFX0f/8MotSMPc/EJtGS4YXx0KfzG28v5pp
dm6VcPlyEUhiIoQEEjqtuS+rLYQdvVVHd7J8VR4ViavQf4VIam/ggyqu3/Asu61l
TQeUQms6sOZMBaLqyAO1Z+WmCD5gexKntU81ScA55zwDBYpSU4BRyv6T52LdMe3r
0X1ejcLiGtAGgHVAsc47mtsRWDYvr4H6gPLbO1mmFQ7A/FkPoWMhy30c4CoFu+M3
2JLNZuQ3wYckObGqcKK5XzkghuAY5TwLEtJ5m4JgmIzdlMt77Mto4WGvklfn1WtG
BlTIkCxEKESWHRT6iXaoeD8Nyo5Nwu5Rw6CeP2oxeTdg/5opNY8ffDmuIXQ+o/4W
TePPz5ChSZjtfLaaxvGWzq+zkA3tYyRTvzacYYOQXpM3VGj6SQ/li3sP1V3MgFay
2JR9mndnKJSTEqfqh1Y1zB82cYzwnfd/S2022YnO+Oe0pqrn9LaerXYMyzzxdPWv
gtDO0Kd6i/j3wRGZkCdBv2lBMDjQeLORO/h+xdeW494q1SoYTf91kRkXAt+Ke3BS
cj5l9S3lwSH3EvtaZTiDSpnkcWhGBv+RN82eMm+IHx71p0TD2AxRs/6n8MV0amsU
7JngBPA0IPkxD/jLasUEjwW7oqMgXjbpZIgXpFwPKPYpOOhFQX/Q3QyhTiDygM+G
MIV3CS+x0X94GtmgHMIEuMTGFS0Ag1JqtXEw/rfK3wh4hy9jmk3iuLmMpiw3dG1d
ulj4geegH73Df0fRuLGIoWP0/TDILpdeUl/TpVnc/nGIHMpuhGRbWtQVoL5Qb5Tq
dWDptELbLkFeTe5NhUW/LRFmwl3znOtwfszgN4kxB9jDM+lUZuiydXfiTPX4zhEQ
noP6O6abUadvLClZlGJUGe62TVNdXLv210kh3IEnWni6XLndfn9iSkyIDaTK8TEv
eY/K7i04Wtlg2yEePoTSIJIVBMkt6+skTkd6O2yA7BZfcd8uDXHZSkUT48Dmm2H1
CAmUsNtfc3wn70InSDUzZJ5X4xUqToV4ZG61rkY1+LVwvmYOs7MgbkU9yFxZk739
WUQuHkEpimwWwmBopjuzJX9qgxf5AefYg+VSwgoNKUTc/rgfp/gGCYkc/dt5KPWs
Fh9SvHJbFhyxGHdG7h5hoZCEBpOlbxyF7Clc1e9S3XQNEPwHbCj+hQIPywv+xOxC
buvFyWXEbUVonU53ol3Edbdl2OVo08HdU1qYGxFo2LozWpIf2nao3pmz8L/EyyL1
sFpGo4cf7H3Smxz94RNl6gEG544JarKTSZZOTsRVcPHEEhk+6iReGTCaYewXo/h3
lFpeaS/3TtOZtl8s040rUO46Ze1U2OfCUBj8X/YtTM/Jyw2B7iIZFqFcIZaixi2p
Q9Y7EuRmCHDNK/5o9lsry6WvZ67z7gl6C8k8KFcs1XLje1dOzTnTjiS8iLuC0jGv
2K+umGLrCxuogYuI8fXdsTsCcdtr0zDx/pAH0UGI3T9L+2Pkgc7AhYUHdilRLmbD
OdeaT5CSR3a2LuY9LncWGN4o0BBVQHSzNVmDnge3tc+ppPnUdO9a0WnuNpSIpMTX
QhB98XpchTUKTTqk4Dvv4w==
`protect END_PROTECTED
