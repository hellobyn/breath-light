`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFYw5bsCSXpbNNveOiDviPV4rQYfARAGmuiMOmFAWUKhJZtP5DEiN+8s9PAOB+HO
H3zZam4xsJllOCOH2Jgw5aTOlXg1GGmCIL7Xr5euzmqGjqmiJesDA9MbqJQWBBaF
Wpn9ag3WJG/yZ3lb9D19YraBZnT/YnVsUTKOkeXOcsf7of1sZaP7pxYEzUD5Ah5u
kwbyGcpoZE4zovbyhx5PPZU7Se6ya4s391kIsjMmdzY3d5/WpPKvcZsbJYsjd2+k
9IDrBXLPHNwpca3PpRXjCHvLPrgaDiXjfVUeiqknvGKeG2oxc7DaiMF9A7ySq3DA
UFVeEnr6CIpkLkBH0xcHpFnmc63K+fu9X4LrZWAscfQu+nXtGzdj0VLQXlu7L6HN
eIu9OtrvJ7Kk6LRXxhSZLyBaTtNLGCGdeHNXmTHsopRP7M4Ezk/LEU5I4KrCAe3A
/GJdXZvzmJkw35jo4D13UTR/kRZO8UWQA6J+3sO5qMr5mTOAx/EtysCf3lDajIvL
7vNMVKdinqk3kbQ0gx2ER8sqOrfOgOH7Jf469nx1GQ53hBRN4YkJ3em91SDFBnu0
pA+ow+FiMC38BMsKLe6CLvl6GcBggnfCPUuxs71Lt+E0wCK0aJbc2ZnUCr1iTqBg
PeR6KiMMh6zcqkga+MoakoOzP+ZUAwJ55TNW8sxDiwSSGtF+aOEJ2rpNlx/6L3aU
uUtQQMGSyU7+sG+fac0dpv05tNVnJ6XoA5p7CuZqHQPr+bnQ4i2Y8K2yv2AdycvN
mIaY9Y5dhGKZDNnn1tDYIS2lHu20FzV/xQ/zehXs859x/ha6+NM3jbSIav0UDMv4
d5AWl6iwKADBh9+9rzd8bqErQOPcg/snwySeu7KE8bEcGz3/ZhU2SI8UFPGPcQRx
69UvzjjinGFcXOVU81A8bZf8/8pHuWfgHK3Qc6jahcP0sIsKLLY6h+DpJLZ0gL8+
SAQNi94XW9Iop6GymBYG1+HJcZbQhWZVBFkk8jcWyCLJJz+bRPfy40r0jlv4U7rx
Wao7KMkUEZ+2+TQFEgLVS29AL7vkh0Lyz4C5+Jzhk80v9tkEnWX/iIZJB2hvnmx+
knWAGSVt7QWwJCPntCsueHs1Hb5I7kDsHaKxIA4xX6MvMaRk1bcMbvmAeiLyOX0s
hB4Shgq//XF4tNEU3NQXhT5jR5lUq3NfoMkwX5VwILT1XsekNGDETPLFjCAZZBBz
Pg7T+FmgIKtSxap2+fXyOhwqFkCkO19MJyGqAhN/K9k=
`protect END_PROTECTED
