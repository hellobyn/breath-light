`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KJbemFdRwWTZX1QxS1evbRqyzuXE00ViyBYb2U3417I/hEdd+kUmMAatYmBVrRt
sAvSOKYFndxldvBmbU0M6rYCw/CIkmAvCclUQZ6v0P9zF0DVcLgQYfx1NXVqtV4n
xexCpSe4AGy1BtylyFoxMefSG6MaqmX9j+6pQwcU5qFux48BPRREekU7VhdanlMO
O0rF3ve8PgJ3ha37NqV11gRhRg+ksdOGPCndf6R3vBCIsOCQN2T2+EgsURiZ1tr3
1J3mlLeBAzG0kMEMoBpbQtL7USn0eynOCigL8YvQ1NKkuTZwiHp0qTsfhnJ8PyUr
9LUSp/KbhNmv1yFl35itA2/ZJm8e/MbcrsBvFHu/+mXl9r3WfcROs/r7AqJtviMU
QRHfJ/zMQY3kxiIuOV3m7Gnh4aE9ODP+lSC1GXKBkH9+EhKnDsC0ETa5UfvuMGn3
vemJLhqsuPtiumrycvxbpfZ5giObkr2IG0iaEtI53eHdSzvDtYQKTHgSChi+HCPV
sjLylIIy6faxws1rFrP5NMdC/DMfLzDw8RCAVfmGRoEBy1t+WxIgAqQTLxgtDkwe
vEDAG3Zbxs6pCxt0EjtNY+STBlWFpFt7otw5k6IOfXIQm8EamhPlvtowXjEie2E3
DeQO3T2bZzU+6reqSoEI8ua2WRgs8flzSDLyxQbOlD8GKgD17OqcS3Xyuo64GF57
o9uGumxgrgxqRjyanx8PC/kYPclFBkqNwcGRU1RycfZo5dGVldZAkARK/boEMfXq
XaOGONRcVuSudDSGKgCslR/n8iRl+AHU8CMC1/OfV2fNlPOaaP6k0ASQh2v20e0k
FZPkqFMVd/iyDYpKvr3CCFZlIvphwuMaGEAXLkLELQOGengQpgCBF997QLAve48U
VuhucGyY7TjYP+CpQ1ZP0DWlO+aloS02YE53LwIoyf6RNPjeN0fs1RFP7owSlCDh
ykhNOgNr/OgtMnAW+oN0XGMuzkGLWSAwqyP5M8MhHuULCIl97ig+HY6Vm5M/SF8T
AF6qZHG93UW/xnRllHnNAHOlh8co6FEwupwkJmZKy2gcmzcz1YEuqEVcVDJsPQoE
NszQECwroBujKiMwNNhjoHZLF4oTf6qEzMbcN30oS7CC32/H2ng9LXGClkA6cOau
S2CKxDj66+O01GWuJGThpd2SZ6oRq3M1kpxhfoDNiqX/L7GtUk4zUtRnkq4v88tQ
As7yXYv5tqr93E14cWcjOXkpHVhK4LzngdksZzf9Uzw3benz2pm6tmZSMHNaaEka
yxgBinoQiS73FbYfYysXVipz4NdE/Y4xpzegNv0TCS2VQIPw/ZDenkliNFA+Y2N3
rIZrL3OaEe6jn2NGL5Aol/vgjvO/1ggc794df1sh17bksxPC+CUOokMYSVGj22Zx
1gCgJevRj6GoRVyxGZBOqjnb9Mgqo1AZ+zs8NdOMw/QtAk9d9FIcVVOU9AlQvUKr
j0PFp7VdLV+XFjdCQvxrQfzWZEovCRVKy2U6zxtx1aft7oKDOYFg58tWYy9f8taa
TKzWv6fqD3IinpXwYiTL279u+hsF8uhmlz+ziJqYG2nLFO6IEY34gVqBF58kWM6f
8oe/7FtR1kD2ThtQ/ZdZui/E9kznC9yAAw8WRmAuIzn1oPntg1+1AzQkit722Ajp
87k+cWFZa4ipnbTIapplc1TOnaIPcxHkuzZRxL81XcQ7KsoR7DsC+xekgNvtv+yf
zIo6UpkXfNlKN+wCwa0guQclFH+K6eDJPMxVAsOJ8lNj/bx4N1686QbTl+UOoMY7
q3xjVrU23YFdkj7jKH6+vE+tmhkWEc4uBX55lNVgvs6TFuOh2fjEaO9peP7oASSJ
5JhC7o0EtII+VT5BgKuUQL7vgTAtgrQh2MjdKWrgUigeoHE0mMns8B38W3z2gW7M
B1lv4DwWtKSY9QtjwHiOfenkvpIkgZVE00wsv881sxhhFgizolgnE2pRsWeXP/V7
iPyY5TUAzCFHmWkxFlQh2mwa86pAUtYRysz6wZVGYPJNQX+oFJZ5icTcVCce0JgE
+tlQoV1Qg34gnUP6afNya5O4BQkfo3nSZB735EU1sbkSZQ17Cp9I/kzH01KM7Chj
k5O7ae+HA5wH1N4XmPJv/8G6W70lCZJlfLtvSUbps56OIsBFI7sz+UaOBMKQhTdB
fuPKJ4rTCB/al4htoLYNTLDkUUkoFILuMtb2WmaHxdLLbGFq/5JI/nM18pBHdbs5
u2JStdO27w3aSBm6swI3P8oXGYx/tLU1B/UE1fVO5/KKQzs+zj7wSUlQMJ5wSl9d
F8Kzruvd/ZgazQLaJbG+QqiS0L57mJA/7mb9Wz7MXcvxVDdm9vSfw5TRzyZOS7CV
K6D+SsjlFKUf4Ve+H5/tn9b4PDICmvxOYE4kgXyXCJYRajfwKdQ+jUPx4jGVAR1L
6Iy8wVhNFOzMhEXFR25x1n6GiV0zuCwV+ZsI0uvlCGn6x8FzFNFb0xSVUKvwp7GA
27sedtZ21dk1yb+1vCl6sULa0Ug+myzFLwUkioSKVMNG9RaT8gDJu7AZKwb+j9Ek
Zk9U63mXL3xL7SDqgIjnEngwZOLMajAl1N5Ck68MEfjYDexZkjcquGMbxiM1j7Mj
cE8lWDRs54plZZRr5IAo8TMhF1mxaYkKz0oD1qfinowWScrRqoCTbfUXDOzbBS+y
GMgPnq8NnDU0auoBa7yveEpmew23uxMex5rZFbNYnpB4ylH4YmGlURwf773aZDFr
dNXqKuja1jI03AysDylRTBBa6ehmTedIGhdwGmGZ+oon/pCLFPgnFbA9M5G8/kj5
nvG0g17WICmc+jNYbHU5sLdWTE8O8cCQZ8Xs6HgSaCvHotjCT59U5x4VboQZOElg
Pr6Wgxnos5f5i+UIrjLtvumLfo17tahesQ14UAuBI2KjZlVgFIqZIw3ritRLnVUT
2PJG5ouW6cHGuOMGy0CABTqL0QrQ1owiWfgVUvlHG9JqP59D39JSsJ5HxkiBMjLd
+v2pCZ8tvy5Z2leRK2f5JkX0jxE7H52HVhttB254W9r65REIqiXazzR2cHZofqrv
IjXzIe5ZB7gGKU7ID3i54b1vobd7QkLZGF5JK6B0Tyh1AMtq5wh8ejDo8Zwp7sHa
Ceo7t/7MMhlVAZpzOHrWO0u6/vOAOZL6kTDAFGEJPH+H9spWTEsyGKuVPMzW0QeX
QLVjj8zNLml4LEqV/AtPZi3cKBDNxFBtU30ZlCdlmCsSWtGk37dmfqGXTnYiV65C
uVNuSDJpxn7jUTGSD0KgtWClzXOcbWnhSs4RKo4CYhXUih0KBt/GcilILxNDAljs
IfZvnhUMpNjdn6V0fDNAWUCfY+RHfl6/vhu1kkjoHzU9clvArKXLQ7ysFYUkWtpY
yW4csCOZmr2W55T/ztTr5ejTQG6TnxKjWvAOGmOQucWyRf3X3hUv6OTea6RvK7CZ
rdY/tSWds6J8aSyOLyLGWt7xPwE+xR1j90bYOVl7+TXAJRNG2XudX8ayVX6r95hx
JHzP8bMlXiKjdmemoLlaj8u/slNqmzogm8jc6dcsrDlaCkcYImaadkDqFXMM9wDE
EAk6WUggGbdNqVckzLjHIzg/QCNzGVV5xVBFRGDQivP/wEuAqOAu5DwO95UoWxB7
q9ANjFTokkCEqSr1eenVimpm7ewLdBwJaoYqsvj5BsEbxWabEsrGxRs8avd46pWW
/hhKsTBm6k6xUCqbDcpa57t+8yvvGVaaOSAxzYSCn2bey5RQLBpeYOKcbRxxf69l
uNE5IVh9as1iHGt3eqwFccv6HiCE9izMaX0bK0FEqAEjqFshGW2RjOMr5id4+1yM
WzOlIRTMjqPhWPS2LLq22ajHsqwr34AyRZNGBO4ND1G85KyhelsIoYr/kyNZGKVg
vTYf2wYHOSS6xFfEkJOgJsIg2lPQ+1TP1aBtb4si2rBnQYQkUsYHQpJC9arhyPWU
mZ3UWfopQBqOAoxry9R2OWuAhZgSNmaldhCmsyCy6DO5i8IkEluaweVGCWiuylPe
FEU9NyPhUAT2Jo1m2kKQo8JbYUSJnYhkYUg9qkakX5kySjHnmGiO/r5NyDIN7dtH
kP89tfIysfWeGXTIwb8MkvFM0aXayOi/nhub+0fvvl+jutgDyXLoUvgmZ/frrItn
`protect END_PROTECTED
