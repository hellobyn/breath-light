`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWnBvKMMdWeOasx5GJWlz+84B2KOiUcvSH/kBE0Z3GiCiZQxljk1cr9wJaDen6e9
+AYXIum18yNKWqjTyGARxyTj5iCOM0l5sVH7ARW2OpVvwD88/Wn0/p7whXEX6+9E
HuTmzVDWpRq3teJDtIv2Uq3Kp0U05NxIuX1m92naAFMht6YQ4Dk3Fe0RFnK12I5v
pN6p5uwqMbKg4OGtg59KKUqhCyL6yR0LMu3uy3qJlk7jHSKZ41YwnPKY7/YhDga+
aFSHKhzgDfEFc7eSouv31552bPY0pHa2Sk1ZHe6htI/5Mar2VP1hzZ/5IGkJGxWh
2SiBhf04sjfDVThExAw9jCc9D57d5TBMlTMDE/eUDwksd7HL/N7Z14TLOT+R5+pG
K+xlRAV6gSLrGGiKtmyvwfA5NEw2MVj/xUkCDNYYUcIDSpLzT092znEAipC1VN8u
T++HV1oQZLSJnqDjVvL5EbGAiQ0wZsqYdDL0QReovR1IORdpwb/EP+jlrVA4i81d
0r4oiyFIPL7smnZ/sejw9ukrWaEvEYdXDwTbbeCB7K8QNqynGcLyET1ANUqDqGLk
bmMUaWZ+F1i5ZwVHLwrXngrsgXV390cREVVoiOKaKs8Fzc8lJ1WMzZG3VnJZI7xP
0atVGVFfE6CLHEGVv3/BfLu12nOOl5ezRdm6mMshs1lKLMZse1K1rvxzh3QomRXd
wpJ8fmW/wCtATOj9FlWqADRIsYK6RVXjScWqF9wh4VVScMieVNS8H/QU3vhnSJPQ
7ccsApt/X2daVRgjhRvDjg==
`protect END_PROTECTED
