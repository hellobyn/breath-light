`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0JR7l4cBQMDBDqrlVI9GkcLmLY18PHEut17/xlOQUSSSJ66r2fbJU108Arujn1y
3YOc10zfAbv3ATzQ968pw6d5WDWyqfMHKS/J3eIM7FimOEJzL2m6/8Gg7j3RuPu1
I8Ne4ETX3vCeJRqSsLuXJeXeEaK+Fh63lesV86Hvd4Q+3oyZYTtOu5X0IHxFb34O
auGzcXAsRxzNpakJPX3wJNlhu+KwdGbRhipz+FgX2w6y+ZsQ4FI6QMlFUBv0DVlf
kaE2OyBgjeJoD/0ZkD3804mEnfpOHSZv5NLfTn36ZBwDCg8Q5F/KwSmrre7w8R3F
0zQDGQkmd2splUG9qXb1zRVcHSUJZmL6t4Nd63XuDEKr86GUO/dipUIogiVGvSHx
YBp+XMSY9TH1r5uOg0qyKGimK/Y0aDBUK0Z2pcn5o5vOIr113ohoxoCUhNYAcvSw
/6fECA2cOrsxHPPJ3AK/dQz7T7VGZAovStpPjnGa943kC0/eYQiLrTDcFZFianmE
1389fSXRog+fxMHVwjHBxY98KEtC47ecn0PQ1FOo9Ji0CQeXFow6hLhzssN4o1Mr
K5SEiCCUTiMzWqj8mQxJCCjJDjOae0fAomBWSXkU0+ky8sE4IcMm2Yg9qSGVRfUq
7DUtjHBjdziyz9I0TxApg7mcoTy0Ti0hHJsFsml00HHJWfKkNk65Qug3jF9BXJ+C
frzYP+kE6DebLBmPuhSHSPC6NiswTTikWUm8xy8b461BiMAoZVzK9p9xgHhGC49B
`protect END_PROTECTED
