`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsgdN26+/R4K80v2fe9MLXbaTdIh9ghGToG0hCgKUJve2z/ooDQrxW8+B/MOEe0p
O6n3Sk4W2kOpolBWIKkLMSSG/3OJvW5PeqGaHmLlQOTWHO4Err9nDfZA43loVnqb
uykZ4uSmfm6b2Fb4B25aqeoJm/aFa3RDdjhewou4kc0oS2af5MX/frj3w/evcRGH
MWWd4EIu/rCj2159JXoq5r1BaMT0JWZ+ZgPjSjIRA4sYBMwgt2/EPMZirPKCCchZ
s1CIwsZHkOEWV2K9oNPZB58qXXLfAZ7gsQ9xJje0h+NbPIjxR43Ma3bHXJECWL5c
lhNcXv6fq98n4Ct5kyuqrd9+oaaaWNAht/5JH9hkecrCDbDpfCicWkymtNqd2YPP
sPLpogj32OpUFBPqeDs7roXOydD7HlOAyLkDBSvjX5sY4EV0BN3MOPi9uIZw9W/v
sCoSHiKzuraSpQkBI30H6FM56BxVjJM4IIO3b5iOZNbxYYG0ZjuqeRXVvWXZkNyE
q9o8/jyCpu6cIrq5bDlhQZYIoCzaKxfUvvZzgtlJbfmYuHV5sDITAv42ZRuhF17s
l5inJRR7oZQoNTgjFI3ogeGMPl8By7gFfQSOOznaydq0kdHcvxG8PNQ83szuWXQl
NlKkoUP816Kvcg/8olpjws9X/zSNd4agkWpvQaffo9sUiPpZPzz2JjKU/ikSjjZq
Bv0NLKqP0MVQVz28kfIAU8qXzdRAOhJU8vzkh0yB2qNfJDmCHyQ8XPzCYbQIMGno
to6UloRS1XxQePFhmQ1YQ9X11u/OJVmQwVReIagmbQ6QWv+l0D14OJ4rm/jMVCHr
9kuGqNeokuMBQkAB/rNQzoovrbLhuvUB76g0uOgnU5hXDEsVQE6gjIEQgNzr5SBw
ZBJA9HsdjtIHLtCuC/5VyjSEVES+fXRIzdnCDDv7HtaL/klpasQ8emPEKjezNPRa
AN/bU1xbIEqynoe/jD6+xhFTEi0c+x01Chq3lha5uUhFEMxZvD/wR6d3RsCswbWD
z146okq1l9I2ArLTK/Lp6aDLeI15LSKG0moSB/01TAkUqxUNnJpu9EMe2fdMsZuF
gADN9BIgcuuEmhOHW6ZfEZ1M2Uw1FGPEKaq1i5VKPHZVmckjhcSp5hzvWuU64xij
jlYGlnevo9MmCDPTzTpyBl+ao2WQq4aTUP9w6hoUl9HKnKZLbqMeCPY6s9OWyaXs
VbXf2acQmK2J64Sa2YTErtsmGd9P89dXP5KI9nN4ZB9o1ufppgidWpCCJyUsPjIZ
MfXw08hEJu0N61RTOiFkyUflOXrECaYuVN/fkv7kJQr0FGpD4A7gFrUssmam2NoV
u6YMBfegj3K+sfI7UdNxex+XLvRHv6GHH5Y4OKkI0bLnPz98+nt/qo0+MY2xiFJ/
WjLJhXE+E9zLvUMmYfKtxbZcnFbnhxnuAvG524Tkvqv3AYMoTp2i8mj/nCbaL0tP
kY8kEooRmKgEAOVr5Ag//vEdimzrjsE7su6dsCIE1wJHhCKvimRddUTA9TwjMd/F
onYeZDOHCgtZ5CEoESsyvTVJ1aPP5NAGYiqBwj15u8tLxiLc5zp5hetj+SxdMM7U
j44TahFX69loEspzSeAi/78YiiVBNRSIY1Cc0afpHh0=
`protect END_PROTECTED
