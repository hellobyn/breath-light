`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGksoLxV5LFuui9DwUgOsArsg3lXO6jSTNPV+Pm2FdPvFVVlJswuNyRrtarkQ0FZ
OPk9XfFnAExUJG3qojmb9U9Kc3NvaCFcDQrPp2FyKtFdr+0OcPJrssfiCubXdvfG
D9ou0Tn+lIkV4kwTQ0dAy6zFMBOLSisgtMqJW+md/jpUc6N3pNV8c5DztUoc/aLC
A+PbTPZzSN6cnccmr9MXEcJ5OtjAqLnmsEKi7nKFyGU6mD0k5iv+zIYfZmOhrERG
5jOGLuaRco1/UqAuCNYoHfuubK/ZEym/uxV1TgTPZQWRxgO2JXeJpwVk+KNxcuxx
wudpsqk5ynsThOvsMXqFnLb6sSisThy3oZXBlfNeVpwDO+X9PlOwnNjQBcK1Kh6G
dPEwXKjiUY4ueBWMGJtaRhmMDcjYj7f29izd8NYdfFDI6q+/ptHEDWtXrY3ccyga
jzQ6aZUooTDejNggA30MDI7htnBZN/Evul2rvRm64IYBr2lp2DuUp4jsPr2NAG/2
gfc1mKmFKVa9ka02UaSiKnvRQehlAqb0VYCfQfKNISRlqlq97Cj3o8KtQGzwTKSW
n/oHTDbRDBJXCyrHmEofAfwIEUhVdgL4uVpgKXW6JPsmPDkTPBsZPsZWq8jdybzP
6Y8WQt8HtxXlWS/GhF/c/kVuVSBKyzlPFWZkHfRPQ4GaVZVKVKbMew7wj5RPN3hL
Ew5fwJG7RaLU+vJOSM1lbhk5+iNknAb2MsrpvnS4Z0lX+Lup2wdRM2WaZpkUTyVg
bw/clfd/tIx6IenaO3XdNLcR9XgorHZ8dd7ttRkpWcDNVBKQuiXEXmFAwZseBUA7
WD6EGeLQ0sNea7fJdVuQkoz0bxaOtCIKa91HZBVjNohfD3wqpRMXAYgs3FD9gysL
JU7rLzI+0ohmcPAuXm9TrSCPKgBzKSql9RKUXzhJNwU4uPPSlR52HfP43xqWviD+
tlr6O01NEUnWzuM2+nm3NYcaN6WpAs9pZ0EPCRQOchbDz9BFjB9pFmvNZn1EeExY
kTupid0Un+WoG9dCnEICf3nJQHYpHOzCoO2C3Vya+UEkhZsYIqtPM58XMFrzsHSn
DFigpGd4HLGmeE1MBNVZ5NjTi8wt+IfHlHvXo556JfwlKzSQJt1ChKqM0ID63Wrl
ibOkqGypYmqvIIGv5G3CYAPnGa+P03tht9vboCuMceEOIrRA/MxYSZBg4WTo8nHf
zMVbdtHbFOXA614wr9VRgxUlxR5IUfHLBmrV1y+2/UH1K1uX1ot2kDulXPHONI+Q
qe1q8SbdhGkn2BgkouKKTuokWlh2cvd6jwgFo7lcEa48UM9hAQum5e5UoLbxhxck
axVKf0AGkW7thamAdkeiFnlB4+bkQHKGg93bKZfAIOrTLbTXFSxjxW+ky7G0ezWu
6so0fKz7H6dMXsUFb5xUCthnf9tryrUlY0El7GWoFiI58mrpC//bfDJZJX+2xYcO
UnkyAvwsmAuHRofHvX6yMNItyoI+ILRPDqZya/GNunBaU3OIy7qIUXZqvfFNQV/Z
plN3iDsDGC7WH5dqqSvdyZYK85WHXW2+jsuLS6IH/pgQhd2vLW73I6vew2edtg7W
sUk4CEwF069Jgb8A4mCS2bwYr9MK+BVBvij90qBFEIVznpuXCA9lyha5A7+vQHV3
XR00AV0QoHg69Gp0vzSFtgPS2LSZ+bqzBq2KX5hGaKnLOyVRGSjuW6E8keDnbZF1
IkYSOgswycdHtqHf5gHucDBFQLVQBiDKmKEnWl9YfC/wTwsR9PiOjeK1u3VRqZQv
Y4fjf2LjrPWzHDJfk/SdibmrVGPRIzdB2Ub1N8J5KzvfZXN5lQw0SoybCePkCq6L
xH4EC6smbYTHt/9eLU0W+w2vhj3MDyBAG+PYyHv4wBx0AWylqypksFLL1ZhVbU2F
+0wzhwH9pP4PZTQEaIlnuLfstEJmspqc/ONRgfQlaMWfPp3QDVLxXujiqC2FOF6A
v663nIJl8VvFoyD8jdz0Eb3QYK1F0y46wjytlh2qYtmWYILuC2irj1bUrRRy6+Vd
mmb65MDlt99etq23UHzgb+X/7jGLi9+I2Ex1Nsqql9vzM3L3TotwpM1DBYJZSQmf
w9RGJss13JI24at9JCnSaZcIQv/HA5yDQ5soNn66QLk10uLa/V8rjR6NRWZ7n7ML
GqtYV8RstVsel5fKpqWepUByDpLE5lCB7TGzLBFz9aGCoJjgy4/iNN/ejiBC+2/S
za5MA2QINQsU9NuoVS6I+7r4rd1ZIoEsAJ7MSQy4QMYzZEyi1H5rwWqf6azDdPxa
zeRNFC8c8FtSAs01/G2jlXtI+gL3ISiDvRtZg/HUgDYatrksad0HSH3nwcfRx8+Q
akt8p5H4f2s8jMOQ6vckyKc1qInmBzTgw3kCRpYq0gW88pe60NHGNEN0BGaJjkQV
oNn9pJSdM+/SSJUAc9i/RHh4WOoTME6ypGqVRTcRw+EMpQ5D8KGBMM84otJxBEom
W+BAKLOlkDi1oKSmYFK/qtJ6183tmgFtgXpkg70TwjGAUCKwBJUizWH+Ih3e7f0i
LNUbXsCDdzUCQSExvG5zvPdPLY4L37Vhd7qGhkt6/qV+jjggLVzxidCbnK3N0IoM
kNz3PunyNhNTYVl0GXQMn2C2wPiCXSWAWSorW2zdUEXPgXvtIjG6tSrMrT7EzYmE
wwBlKXa8493SGrST9r47AlvgNiNRXgHtJJyE5hps+C0cHGueEPRbTVsdPHZCC5ZO
7/qJZrnQsN+/nJtZGs0nILlbYTzsdxH02RWIMU80SDerNlyBWpQPaYorB05iC8m6
/7ufmZdR6jqD8z/AZxp7qd6mVAO4irUFbM3wzgUWRIQ4C1oF//7Qlf1jEsUet8Zt
5nRxg1Fe4AVQL4mZ2Qa+vDQBsYwVgwJ37C5b/Zoid9NAafBtc1O1SpiggKWtm1bm
Agip5AvcJBQ8/ywCwjYSA+BoODFYicdawggiWsQl0aZushA2y0Cfwte8lT1R04qw
rXwbGf7/fYz/+o6U/KSETJVFfhYwRUUCVNllpPBuYG812CBsBQCas8GziZpbHis0
TyST3oQAty4cPOS99QhQ5AES/9tVBgIBI55WL6HhKlaQf66xOUhkXDiQLGWoNfLA
qHqn5xrUM3kr3AoZSFiW5LBVA6fXVRHhVG/96JDuNvPZkfLmTmegpPboGbk+rSze
dLvmv5Zr//qORm7MGpBySofbBz1lgIMW7qqFGq3ZGD+GCdAAHefa9XY2sKA74Ht6
+KGR0qzVh4iiPMyKvXEdlyVDZp3ABmLzWKJdlUYFM+uOQJLaLNeknPmQfH20crxJ
UPGi+nC9Gn7k4TMhFWTWjATzU8eJOaTfl4tx7ahD2dGK9aAa4fp2i6YzJbkrmadZ
a2tp29Sgv+mC+OjBRX6hjvx+NGdtKF+SyidQKaC0+woZ2jycUe0X64ZXiY8bou0j
pzdAenhNIymjk+fAKS53WsQ1P62sbx6kLPSExIhSrY0ebel83/v5l4ijJHWVxhcc
OIqwwEijhzVE5HIF6+SSNlTzQwTETtM8mzwYUBQ0OSG5ioJfuW1gOOk7RtjWoy0m
2CLUDQ8r7JefH/11b/CapfnCf+tLUaQN4mtYEKxQ41aDzzH3C4EjA3SXG0Q+v2a4
kJM5lQfwi2gCfPNvg53ZOnlkJEx7K894fmlRg4cpKG3c600iaxynejhjA9fQS093
R2qHxfuQgRgQyQoGXkXLgYFg4xTwu/a4HZFhWEZCJVdQ6Qe4nrzdE9e7MwoB8GyX
+GX5lSU9eZISp4Ajnxany1GumJmkcgBz8oVqwb2ONC9kuxr003y96bLzedJiO8bK
hCS3DVrgbO4Zunuspbyg/0SSUWlAfy/kNPqnOvpiRH4DT1a/etu7pdGdLXv0Xfwy
d6JUILkrRGyCAAoLJSw1dbfejvAG12AworGm45ryRcpfmgzMqT9hArCryS2byrcd
1EEWKTeBoMQqXIbYvD1pNjAwmabIWQ4CCzXGCJkqQi2RH5pB/wAV8c0mxiiQLGSa
1oO6lFeakzfwisG8uRQCHqgY5cCdYIooJd7LfYRaYE7xM5TQgz3z2sMNneJOaY3/
EOueJ4qAFqEG/DzI72oqPDyBIo329kwffR94ohxnRoCixRhfaRtM4tVDQ6GmrrZk
NSCTGJ5OtqkVPGr0QiKB1utesX4DIPwEYFUNRcRmxNd85eR8gum1sKaKmrJvbTpB
QGeAY7M+nFpQc15nJKI2VfnXBymrj1kfictTKzhnMHR3JGM3cdoI+MemYyAiDUDB
xo6FxYymQkQSwOpVx5oLnuCBCKJXnCIHxhDIKVLfFWvHh55qgVnbT8AzhIprXz4d
U0MRsMTuKbTmv/mE8iHRbuPxlDxFvr6em0F5BmTDUjPBQ2pWmUz78dHwbmq9d5iG
bzx7DQ+nbih0XfCymXSzXgnf0J117MGXN2KhdCkaGq4gaPCqSGsr9F8ahbmatq8+
BEjDc2c67jPzsE+jg2SWdQwMVxnOp7gD6Y8+/mFXTsxav3WgZtw9Zw4Be/STg371
8WqggTI4yq3jjxAbDjqr2HiPUoFJg4og8D52jimU0/2zbL9K/68faOFN5UPiQicI
CHNdYykJL/QMCpOa8suQd4q/ip0XrT4TmTMr5nTkxriUITu7gIFUkcrzRTTp0BE4
FSCXZIyX47UaavAaip28BmUJ1pdAIBf4ZFe/bxwVRVEuugG/K4Yg+9C7Mb+5RC+i
oGfw7dhJCM/nfdQwfWCgftRmdoZS9EYGMvvayCgBxZEv+5WirhT7dY0NtVOPJgFJ
TaG1wn1F6KrgTriqZ834EnXaNE1UPWRDsK6mehKDLDsTQOMGY4koSr1BCR6ZoEyG
4GTGj7VNSsNu9XMStW2GYqBatPHud3vKHDjTzNJFdeD6+59DKLQHf8xQdqXcmIgN
hXxR4NYaloN6Wscks9ATPAIwk8VG4gHRNLZqmeYsb6goXdAkhJ9jxAH8yGPJKgjU
AzelF87qusp0fWbpaTyW6pPM3/p0cjKteQJvHnasUdED/8NOkB+dThRhN3OTEQUJ
BiQqisAqJLLRdHQaQrLazloel19a7SGyZPUElGJHocGUTnWPoKyDs7uk079rPupD
qpa1tfZQxEZXczvWUcwiFv+qu3kXechJYIElaBS4qQ9LAchW5Tlzm5Q5RXkLXwuW
3ClP4lVSnYEajNxeRUeH4P+FAC2AGa6dUNTOz+0SbLNyVnhBrN+7X7aYI14HKs+r
tVM5MHmJzDkmVvrFBeMV4nzwL4TJlkyj+MV6vyY1704p4bZht7roC9QaX+kwH3bf
SeCXWub/Vm015GPZWwELGNgEGZFJPf4OEKf6k81k2JnZxosgPAJL/ab0sxnu2K+Y
OyZML5opOUcJ3mHlrokyG8KrFesjmri3BQazgnF/ZdASk7owDyslQUWfams2CWg2
pmWngpxkVcDj8304IgIzAFhV01+4Rmjb72Hdm3rXKlEQrEVO4w8LRIWa+Wk5I+Cm
9rFVmgqFGvXPjBfwc2TS+tORkOmUZX3ZrJLPobey065Sa8SxsCrbsI/RGHAGYtJJ
LTHaJzbfp4KJ4BW/J2e5umaXcfGzcffL621fsy6cKnfYVPNN8YJI5nS3pzfN2P8Y
g27PyLdtP4auDVhbARJWyyKagYIzjBxh+eXwEwGt3cTBsxHzqG96F9uwV2p3fCbb
XCkBGcH+vjJVxOFwCgls1rOJ6Vnx08VnruaCXXpbiduFsrcxC+G8sVwXGHJpZGLr
Xwg0zwPQTJq9Dw86PgXLaFAB+aq7QUi1v9+ZWsRTRpqcPkZSFI2HgRcRH2BlknV9
G7M+1dcQ6thSryW6OBCwWt+PXegALopYzBIYn5Aa7sC+1CzxKsJLx4Ilj2OsIUf7
mEBD25El94Dact5zvUbYzRuK3Y0/J8MWLU8Mv8sCFyBPCtN4kIlHzADI2PPq3mYr
a933dPliMRnnldHDr2FcZxp44d7kKb/uCQ372e7SkqvtTvUIx4KxigUHhj5q2aoe
C9TnQ39YZTp391GWZ3y98SAxZvBTqlc33akEfBJkuCkYlqd6t1YM7ZsAiq/pEzMD
NZiatxZeV06/YoW6mWOA45Bs74WOq1+ul6y5YZbZU2+0ajVN5NM3cUIZ6hPbo1k7
iI09JjBFKGHpnZ7twqS54FZ8C9wh0N7AHbdmI4oOhJ4ocrpI761jBxhOicbUovz/
DJOXrCVOTQPFFYsuDDuiAQhmATG6nfP648jiUI4Ej3R05gRTN3kIruapCfZ4qv3F
sPxAs/mQwALrcMKSfR5DU0ZkJYE5E7j+YJsyWrdlkqRiokgbyS18tOOggq7h9a6R
Z0TmfLrw/ao0smPaGhj0RpyUmylsEzu4PsdlmQn0WdqZgpDXUIWtw6ZOgRQ8XtPJ
e/mCesw3ln7r+P/AUT0fgvMF+5R9nVq7ZXcXH35lRz/VjB7EyJKD/JnQS9eyb7xn
QGzd3XuG7wk13AI8qlcv1b/I+V1GaxiuCNHYNvsw7s7LxINgIpc3XG9HhPiU7nj2
rEA/p/Kht73yRtkYrtHXhAnOlFXAMeHHDdyc5z+QYaiCwcosIJkDcuIYy0o+aasG
Nis7WREmvYLa8cTMhEvL1mJfD75GxqStXHcL1XRTs4BIIdEwJFOxN4rjhnO0eyMo
bc0PCryhBaGdUty2W53ruRfVvY6oJfOVPlVXBW53rXHq5lUrTllpy6EPyUKBxbJl
++RnRIV5HgkholvQXWP72UJc+dIEjlSBt+jUdcnc0sXxf/De1XKi9E7G9CvtXoAQ
m2GR7ATqJwfbsBmiTbY6j31m71mTAs24WXMyL6aRJwkyehW2ZFo1uK2PQeD5/3Ol
GlVeuQbWSYpi7iXnutGydsZSKL5s7sAlsmaho56IfmZR91GcY4D4Od8DCWjR/8cw
RZxHwEiYd3wHEN7KXdW/89mX1+UPHc5Rw0YzXTi+m7P/iI2Gf9wPU+uiAgZSC2Eu
uTleeHjFizkvlfdy7saUW91omkXmo0+ObqHOEPgp5njIy/JjT4vfwahFeDSjIj+7
Y7khwjaOFnpSnGXIAqJhN5GWG82Jl2nN8oCWUY2B5osPd+N3seu9jGHtLTc57lbn
t+wKKQfMYzmn/ltJBsNhj1xTDkd5F7EiuKGJFt6rA0vBsrqtnFbbjz637bObqVGH
ir0Piy1JQN/GOcej/0WbFPtxE06Yrt0eNf1qAgBOmmWWflq/PIc9vrwHwyfaRlXc
HOB7kf15jnpd2tfQqwcwuVKc+Vxl2WUcghRYZn654nJ9QCpHvtpiwlBiLnSTKnHR
xejl5TGGqxZJR83YiuQDP4R3KitB+IuDyDp9Ebq7LbxlDTIdGQWy9zvz7k4M5RFF
/KlrnRwh+1iSo/kCGlvf7q31PcXsrllSH/BOqgYW1ntTMH2xJbKzBaMGLAuR2gzr
l4AO0d8BVPqGFxDUZUL1aDv5COhr4tlp+3mzUy2zWgwfgnU0HRjICm2o1DfKJnoi
zLr3hKfQvsGOdU1LKOdkPQo57jzQtJtnvUo5j3hV5eeiHbKjjqkKIIlGdyQeNkTv
jyOQbUHpL/0EeSblC8niBflDoORRNNUXsbN0uXY845eQgffVIKxbC1b0Yv0H/CjR
7dzuy854bCsSkPGBd16ZULEIEtciXpm4p7710ShE6tIAk/w96B9gs2pG3Ho0/7xz
6VAOn12i+UyTfUjDlC0GCYc/1hUkPCpEpNa3/xUBXKCtltQ4W7A00chW7WIapRn8
PbUXL6hLrYi8jtNL3cSQKqW/3Zw1WedPsSudcEU8YaLOjYk5SpqZ/zlm+dD7sMfA
4JDNDbE/7YpdTMmtZYwoJdfRSbo27oQtfTgetORz1F6+UgKq2IoiJB9BBRRz0Nld
PwmG9TriFU1P89AYpivjfhdpbn/qzhN9dG92mw296p3R6fDxKffJ6p4aLUDzNJPB
dJZQObwgzttGlAjeLIBZ4jwiLBYoq4cKb7NeLZ15lPU6WWO+puM0Vrno5EzK6kKM
jT8tHTseouwqOPLj5F0LVuzur9DtRBmFsZLrysCXrj8TpUeyG3XgyudwHeh/w5I2
VNEiBzFOimMALIY09iSO5v9uTICUjNJJ7XFdZTQiZbCI4wRgOgQLSROMBtoy4CaJ
3PE3AJWK7JowgetTHxG/0MVxjUv1xFjGWX8Y9OHTCRs9UC/BrAP0gLzKWNPmSd14
ES3tOcC04M3L8knH+gqmfmcxpI2lwOs5lEZqc1HQhwQkci45SQqxJ1F4HpZlQkeB
wJ40muG3glNuCueAJ+fUOu3vxgCE8pA1mMWoJ71iL+LSxnQSQdJVSoJ1YnXYsBbR
J5iQP93Aa1pycqv1y454g+CD8AwKyb0M30S/YiXO2yD6YAN3pjDz3dCXZTffMj+h
QjnLtX3JsgsT1mLxYnjEZqjzUw5MwmszW9ojxYChfoewI+4TAlvL7iPRiPzfmMVh
inDeufmuw7vRg1X28mQSHITj7NJIdlAlXZacg2NKObT1dhzw18dKCD2pDI8dHcoo
C4WE9u0usC4lnI0681ZPUC8zmRgP/Z5I4itDJS1UrfkfQEBcxENl89KoKXvicLFw
cZhBji6pnJtXyrnmL+K5X4VRdpLs6dor6QCs3cAEL5IwjlfJ8x3mjiBN4tFv7sll
8O8LAKRMP6jfv5qcUUh0IfmDuq5/T0GHvkFnMGhtfbMX4aCg53fCVqnH1dvKBbvp
wltvVnLE1YiqYg/PB6hwkBM2FSYMEUzZh8axv1mig6YBhoIlAmendSHMp1HE08Sh
NJ1bHsD1ugUaX73T2wxuox4N/pXTvlqn7ZrhgZzp9I1fSkLoS/qog7B4WvRcmeR3
JEqqAfX4LZiTUWNQG9mHktyHY2iRLYaGqlKqNVL5yhKfVjyRS93Jdjg+naZoD5pQ
SF46cTxnfx0YZY4nOWkTAjARoCJ5PjDbzpV2yobGa8w233JuupGuxpHzCQECgGKp
XZP2SMQw+RRu0hk1YKck1NA4NZP9fd6V9rPHxLSMpVHIfK7J6xm3baK1Qe/cz0AW
VXI1OdGj1fI4ZfaeidgA64iu1tVdz7n8Y2ZdgugTTcQf78ZYUVCSOktW71sJRjLv
zFPrWxk7Avx9pm7xVVY14sp/cqwYY1hLBYSzBdrCHhkk1tVHfUPlPGt3BTFyWutU
AF/iG64JILlr5MnGLXFoXFW+lBTdBpqdPBievd7zfmcLovAjPwqwCwntn/baIcEu
JF0BezzM1OGh7ftAX35n0nB+kACdc4sgqd6Rizae/I+xbQ9+RiJ36GXw3vOIjEhM
Jkrnt28f0vxwNhL7XgxKf6QOdeX9yEwLuvhpw3NcKD0iiZ6BPwYca4Xd5JFb5vHz
CzbHyk5gsQWpmlldvyXJYy5A50sNp4EwLkNhVC/jawR5nXlBbuA4MBwkjpktWtXN
sN8KL2glaffjhyMW08XSdtkDHS0VYVw88MAiYf5+tuEiy/OwVG2KjfAK0t6bbVx1
l7oT541HYg4Ipmx1oI6CWEr4tAvz4gJY0Wz7mP2rd7p9doc3HqyeJu0gdmHjcjLi
ceyJ3mvIilC3pN3l727wFrUkSqyuDzyxpw3jxAuEK4GPC2JYizPdgNhDkKdj71Ox
4ZzST1mftZVRKeIVWnGnOFedurBQkhM7puAybw4k/+pvFx6MO9ETW25qnfpvKlNB
llA6D5s2NhyiuvwEvaV/P8Eg7UWTFmReziwGKa/UhFufpPf9f8wALL52RFJlgipP
l/PU+GjiK7AgcYZ2IbLZk8stPg/odDFEnwV/6cTbU+9BpQkkAxsC24PmMWKN+YVk
rU5e6lSd2thm06Te8gh+kFzq1JxzeYTO1B9k4L2Pi8V1Rt+OwUQ6s4l/s660pOmc
oW+pUDpqitLP4zUN/RmRoW6qPkd1GEstocj5WmfMPHHlBEL3Sjos4nFE77MuoM0j
tGuedT7zJi+CSFyneuk4jqaYFXTN0Uq0LzzCURExzyGw7kxa1JcZMHUz/J9AI3sa
4jnBogq0ZAepxZbpb47lBRwVWAlaeRVFa1PZUaCM1Sz3xKe5vYvlkTM5k6emB6dA
woaQuwkzMh0LVqQtUtp1WFOL8e6hFn1IE+NlPQyVAs/ch0vNqNx4t1VO4stgM4g8
TMcmoAfcEmj1YHQCo9fQtWGex3g7fresON0IG5dl+kGBgFjHMUPhQrs0qHceDwzx
VXEnjpzOa7dYioBvoER0WajZKpH+H3Ia2ZvTQa4UuVOyHWuGf6XGUuprEjGRAvVW
WiMdXVgWPrDa9Q7x9Pp/D9GxSqpt8pmSvoG/GANK+KA4wlgQfG9C7HpEkOFjiqR/
Qtouk0DZnEyD8xQTYlsE893kQh6zfWYLYMEX1+aZaqCwLS33WJHA3QHSAn+J5d2H
q9pm+fy1jznV38qmp1/oit9yQEU2ADIgGikW7PhPiiHPq6388uEaWRBZG1GRp1rA
eCu4VYiuLNryTPoyw/oqMSDZLDE8hFW3/TvJgxOo8HIgDC8k6zED5jWyLdfhxoON
QXmZsvggleJ+hQp4m7Qkqt9IDGVJMnAlvmitPHonyo2KBfjSCD9PjpEiSVUn4pHQ
FrH81+ViAzkPgNZGFTUpWDypZK3FqrLXNkoO2hXgD4JJ7LzUE2QB5lL/6CR8JChS
3JZ1HZCiUyPQRPVpeHC5OodBnE8pAJGsehIB2ASuUAA8umSNXLu8FlRQIJ5IBWut
d71ZZKz+Wnaw0e/t+jIDMSGMWuEEFTwVw1yUj6soTlhSjFdcEPGwZNqU8/96HfWF
Rm0e62h2M0RYsFu1KrfKE4Nm7ZalX22EBTS8LOEcZWU1vau7AUaoCADyVQU5DqmW
Vpe3NUcUgTIM44gw+DEpBKeVsRGnIfT1Yv/Qe8wTgJUDtzrADEVtX5EjAao46UZl
H2OoUoL2eywdUeEc7a6AyDE+Pq0tldHmu3esAL0DUfzSHe+UMUjvw9aD0ZohRzgn
TCtXjWHsGb0KzgsReD7CPuP9evm1dXAurHnLfanwdM2MzrrZzrLFJUgiJ3FC19aR
K5DzCFTmLDpHZZqwucZlLJ3dytPNRW+v16UtSCgUkpisx2FkIi3ypPh2yKNqjN1r
MweWjMna+Mi+CAKcXS3VCsMwlrJHePGMiTdAckldmn5642IYsf7sAjSo8hGFmnM+
geXpDXiDmjzC9TqOI5Bxz+GsADMwwrh7pS1DZJW6cKYRJ3+7WX5v243ni1SFUVWz
1oHlempiHsLP111DfAdtD6+WH+KsS2xglgMLCiW2PrtneTAz2DPcwcpY9ohPqjQh
aM+TqjI93LU/kwVoba4xOnID9btjwj+PuahBMKhs9vUQ/XV4Mm2H6HFR7DZxDNB4
ezqns5x9JLheOyJ5rbP/3USCXkDlamh0uf7fCwWVj6vqlGTF+xLHeXBm8/LwqsxE
zWT5/jnx6RRzfxgmc39yXooQq2g7tWWlIbHF3ElvMw+hIdaDRdwn715j35XaOBGy
ESZWrWsnorvkGvKfZLpigVcJrZRI+prr6b1yyHMdr9x1rOMx5Rx4jxF6ZX3FCth9
e8ZliI8wbLsS+jByuokgXi4jTszMaErZS6aAgl1Vq5Y2h74qnBzyhbHONba/17dS
govVHTx50yU2D/I//INOpp7hsplHzPMNS1aT9HoPXKAefG6OMgwQvafqwKpyHW9S
lWbSvxCOwcAzWLD2XRKkHUwFR9DKIpJeIyTwg6sRdra8X9o1ymJMDUCLBf/1Ai30
bTL1tIsnnBRLtizxlYnPdcDsgJNLk0adL9oz/fRonzFb3/thy+juw0UOxybBM3jf
YKTamSixRGk1feHl/wGwWXHWNeKjly5Gyhl9d+iFovs3eP3CkNfBLoQZ72oY1I+4
+k4bmx2JuMBLmOEN83kkZVJIJnuK59ov/kkKaqU87B4CCre/AU/6Xk5XmrmnhtTX
K3H2sfCUhKopnkTGPTfa+L0BtIjczU6aPHQVidt4zwGM3Wa4h2MqCYqvn1G3NiUp
eWlg1C4RF1XL0WMNfgTpJWDltywXYG6Hx7G/3uCKX1fA9GSfc1lOmA2JrvmpcWry
PfpiVwytEW9XKf1VT9WF8ufNvhke61Ijjw6gtr4We26O5AUSzRwK6zRGGvlXjXP7
339i/m0HF5ZhGaD89tP3bQSDh6p01DtOEgMTyQc3XwRJRDGT3BYWpOgO07/yZV8S
V+Az5aL9D/BoXdKf2z1Syszfq7uq8CLlkLN1RzVNgQ43f+o1Du3RH5oD6RwDprhU
Nwu6zKwfxsgpDESAly/1lKG86J2iEh0pRuPZ772utgFqsSvXeDnyQx6nKSuPADJ2
RaM2NWIzNcrYXEWkGEQR4jok1mvrdAFl3aqgtnaB9U8IpDSYilcqJEdmAP2zj43X
N/W1pdCtPUXuXBJC/srAZUw6Xk1xpWhA5aCYdr/lDiBvOoE+SYzUZMCjoiIEbgZm
hWJAw17qhTRQanKldjKYYwrhDPBLF8Gr0Gfg0V/tljyY/x6Go3UBq1LAmfWwr7x6
60J7TEjYzG72YknH8mVxVmXTuzyojZlIylrghSrwPf6CLgr/ulWemRKKSEZDAnay
r9DSBb4R0rdf2DgJ25VzNorUX8Rc4g9DCRQ0ne7paZmksUcth8VJMwvzTGZFpl5I
lXhAMYBgJJCRGN+mHB009jwZD+EVHbPFpLiUunPFP6bF+WuTEoKsqNneUVSFI2qC
40twS7PxEaqRhB6wZvZRVr1e/qHfJQqpGgQYUcSobJ8YylbSG7Xu/lETbdkMnx5C
ZGRFbMpv8zSD3qXVYCae+GTk8PD92wOAMIQtTb8AEcs1u8u5HpRQeAauEUo2qUjk
vO2khbrssQafZIcs0yw6iPceK8Yzngk+SfL97KIhqwsYA4NrTAFPNdrlPObtcRzt
RTtJf5A6zo8zAK/2lv86v2cdNHioWJ4t8cZpDdqRVoQAlBOS3EdOtaxGq/OYA48S
HAnxJmhRcMqOJYDJ/BK0+mVCBqjda7quE1BPSoVlcBmR9gS6hYbqIp9+xJZtNxg6
h8AWEtbOmEt5tG6/+xeGGvq4xVuL99hvYaoWQczpPm7wJPDIICdGsjcC//LIqgis
JqgYndto0CgwP515znUOomE4iLxuZhqHAVAQcRfLWh0C0At+B7EdLSaIXsSen+k8
3ACc2e7Tn3fUifEQwGJoN7yPKGznTFmQlOdNyaRddhKdgpZcTfY3tr3td+uv8Xnl
LB/eqEoOgZlZAg1a5Jf9zI2pFcl7hGBGUJWoaBIRcwc6V1k8GkslVVh6YKqmQYms
VP8cc7UwwgjZ1JTetqjJXP53JsY+/mMVm0TJq3TfsgBL8zPiP0SDV5ff2aEDlwdI
XHZr0zi93L+YwKGV1aJ+P2p/vpR5HOoH7WBsug+Bcvb1/0s1ryu7WjZmeBzQqJyB
J6Uqv009KMZ55RFQroWKdXRXBvsLLN111QyILDYCFTNfbjajfNmBTWXlB0BLmsjK
6sH7jHebpFpmvLG/XMjxz1UI20fAGhqiAgN5ItHzgVxUKVGgiPNb+x5c7j9l5/B6
751cBghZhbyJE/OdLhTT2vYkmIuHtp9L9hmuKS7Z3Fgl9G/lTJdk/o9wpoSQ2i5S
dkrbAyHG+rnKvVa0gJvwCwSU8uWRY5F4d7oBeiWZOVeKomVVRItvvTEWqv43DHJg
kDZZrzRBaZ2rnLAmkYYGvowJwg4VrKx7PoIL5++KDyh6cO5e6e+eTUTY7mb/sy3n
+QCRX+++ZAEtmatJOFGByQ1hmB4KSQyCaglX4oH854YWTib22YBXeKedC9obNVDN
to7G0/I0+zrcuF3+276OyrZ8s7GXvFLzUvo+S4tQ3EsyTbo5/t3Vkq4OU2kHTkrb
4ku1SFXIF0nMIHq52Riv9h5X3PqjS7PW4ldBpI0JvEs+kYBRtO02nScrwSMGDxC+
gzZJRIsjSQq3Nttgk3GJS0ET0G4Sf1AKc4liDUGPXQCyHP1OmIegi+aKm1Ofh+2S
dOAtlN8FvrDAn/YRDZ59njQjogoE2Z90cHfK9xuQUpn7Ga6ocRQeMBJVbzCsGZnN
b8hlrZCKnB/v0FzoPRP0FVnbq1VA7bhwO3koucLkV2iK5s6DM770pLZH43MhzPJG
8EA85uMqsvSo0FZ/btC5BL/LJfUBaXAa6ToyLyekCPdpkF9JyxWMOY/fayfZ0y2C
77EOYlnKmIjHnoXJu8lecNlc2kaOJaLcAtaC8bcgNwMu2qQy8UcmVQB79exg92HB
OIBj69nAXFEAfnBamGsXZ4prHjR7DKriyS/MkUh8p6ADPRD56/0frCuHx4yvLGVa
Ru7kUc0MHUfV1modtyg1EKJFbNvX7p1Y3uV5V36KHNI2lV6wuSCp7c/EKt0OYG47
UEvCNmmzxWIZXr16s7CjWWeDuQ3QClUdNGLkBTExae7XS7uF/QOrgHxn7JkvHdc4
ItI+pyUlADZxcTAdLrn5xL6FrHvrDT/tqvmSfU6o42s2Q3ImU44Xdk3tcIL84bDF
odEO4ZA366oqewc3VTxOUgFqQvAjBvm+NsWB7N2jiDXhBtJr+AXHq+rP1uRVw7G2
LSGbTsV7/grFzTE1HP/QPrhQlHGpzkKeRJ6X/A/NNBAI23a4j33ULjh0oQadOrrC
ARDefwV3AAY8rMg1iDoEzeDe0Gx5REDNw62AVBNei8z2yMFyFzycp7O4hXaLEkAi
box1QWcmN8JNUocH6b6LjQ6jA79L6VTXisaz8dk4J9cEAohiqP+AQVCm/0LNbDsz
mHYfAC5LhBxj8RRc/16VcJHVKFnfPUQaqH7nltBx19htkXGUE/A43aZybEk4Jc9t
lEt/aqc2aeLUi2n9PG+mF2gooo042pejyyVuDCllhDU2H653OPxrFJPKLRRA3gLi
qvX2f33xYOBS9HmO+Go6c3sWQJmW0tV6evEHejzpjXJGYMEj4ArBnfT6z4r0ED47
4bLFeQhZNltEDmYT4x0B00JwwyAJ8L40XBMvl8Vi/qmHnoRhRcXW5ZSIbZLHgTKf
6cuGCbtC7mC3EybgAzJOkNzduojdH9PcqXjrEhvyM2wVBNtDIgMJYORxNpLOezxP
75O0aUE3JPeMZXWp5zxN70oAqK2XZKkOAA0m3uilVWzJTHbfmsWT6zneYa0WCThZ
i5lgyiomzAY192zQxmegfUMYPSW1HuqBvpiu12s2mUiCi1E0T0f5x3/I06eT97Ur
mOm2ccotpp9L1UCgiRIyxgJ97ac7H9JOtu/THt7l41ECyDl2Ab97vVHxvVO5otmN
NDN9MvXltF6J6vGAZRi5KdzDHA52fgj2pDcV+3rL4IcAI2qNA9qbWsV9kP1zV8u0
a1QfWGTvcgNAgT+MVPnw4rOWGiNuUcsb6y46YiYUwoPh/fi3ORM8FHPoqPj6gHyI
KAy4mMqDPodAf2ZMhmnZP/L/7s7SjognkDK8JbEs1oY6UP3jonDrdkdNnqP+LAIZ
jCJsKe7MMVUicdKhKW43nb5zEzJKZA7Jn/4KhJIMSEKGUiVbeY7sBZ3Fh2EqTkvK
tHNSmY7CO7gu9KveTPC5FKP0NZRo0ti/s6UTPZUAJf9+xbvAxORJLu/3sg+/7pQ0
LLlil06tSzS4qyQ7kwupDjB/G1KxNe7k4ZUP4KJ9M/JLbtTWO7lND89wEPjETwJe
4BVDHW0ZWJpj8mUCzMWD9E/5vUnpapuKERmDAdIqhOGQAw0SPn9WZAvvpT/l4Q1j
b32wEE8ZX/FDGVR5Zw0Odt9isJSjqR/3dja1LcV6cTBNNaYYcIYIZ857sVto0lcb
ku+4O+288+5OA5BUX3/8eeWGuuxU3CsoXJPjkDDcP9Eiq2Y3j0jEkAH2YBoXlxBQ
fHYH7wFOBEO2k5CflD2pCKeiZuB8gEMHFEMvSsuZvNHv7FDf26kC+fuN83yfGUrV
0cfwFGCi+GIIckJciCn0oqav1euxkSBd6shD3O3mJxaC0YLTmmspQh3L4CcG4Bcp
9tChp8ZgG2hWjBFGb2PNbjNhoL3QrqpWXhTXP6d8SiiF5u+gVbAJLGoY/N5kA1/q
kvaRloQLKdt71xQsTobexYB7mXu6p5KHhLgR8EP1XmWSU2mlyn5nJpLuGoAyCKIj
ZbDacZQ0ltR+maw9qeLaaXutDG/wAC7AzWlg/eKi0IQLmHy/55tpH5gBa5YZWYqW
aHUVhpttGarnJzJg1GPby2IfS9bFbRKQdg/rLkfvnSf11Jy+cev1/GT5t47/EM36
ywcED4jHJrjXYkA5DABoALZia6no6M4f0K4bTLbCZNvPAUYvGLFXuD5FwdqgUo9M
F7kMp0UMey9BNx8fNYeXlY8Icg0KE7bidy4ya/WD+VguNYbLg1FB3mFSV4ee9pnb
mZ45KNDW04eauYUHkQjgX7U8icUfJAGIhH+FnKTj74uRf9DyuXv1hV1wOuVsCWt0
nH9CahauAcRqQDdnTxzOUbdxNFbx/bDJ+g4KgDrF1OuCm3khBJqp4/9WHd8kHYXZ
z0zJqRCMrHf98Tm+ho4HYCMQW8VqBsZIRV8nKEu1qiYewtO12LCcvFLmyU+v0+6L
+h30iyol8Q2RlGk3ThA3rrFZalLQ21JlqTFJxE6rWPyzYnKRrf0pezSgEzMRcPS+
1wuvrafBHptQo0gp3I5aK+y0rRMQouvEn81Ho6LbHbPHZ3fQueEx484cBg+Nt/lq
5yiV7TME79EKQz+UsL+dfx3SCdJxEO0TJj4PH6hQIzYw3c/Cmaw45WRiJJjJbPat
lhFTqWXxavglgtb3PNVoDAkaZbisoJdwiyW5Pu8CEWhsu81n3MvNBaO1/P3dwgwf
24JjmJWT3dcKLkNGQK26HHdNo5A8/zrUKDxi6wRv0oknjgSFAt+kgB4TVJctR/Cj
6HxCqx61mdMfn+xJrx0UcrjXn94wHZNPmarx3ROQ+E40YYo+gJKxVuTle9lQADjx
vnvxj5rVNR1J+tnx2urhvM40r7i+oILU5cPWMPLHPmge7nWzmD00//9rUKYggh8g
Y24oy5NCLtdgDqlcWEhRO0FQi5qzSc5dF/64knNet38rZJNZBSsF4Mb8H+R2G+7p
4iGhn5E89NO6Uw3xMd2ypP6JXkdGZuCm8Mbi52Gz2bcXTiIdCxVVfn9Oci4sPS5n
eaEX1v96qrg5psAEiiVQDbbHbIciUhp1k0bKVSgvJ3e5sydVr4y9IDqavD/6vZ5q
gJ1ZgdIbH9NLarFC2jiVtMw0XKSE0Y2peZqnKwkN1UEe3/FGldMhA6uksaYpU8eY
6lrBIz3jIh5rO+o37wQAs6AhwjD7iThOuBhpd1lqUxzs3ddHYyBVAKQo/wT+ReaL
L0jOtY9nAqagsmkH+YH8dD0kjQTom6PljxlgBCY+eDfhQb2Xey32i7KQsBoeK4hR
od6T7KSD6are9ib4J5Klo2YHCNHCPo52NH7sRwK/np8bFdleMh61fAB5IwDr8Ae9
1+nr+Gbyy0B/n0acaLp+koBMR8UwMv11hcNna3cb1sY6VwnK+4Bmxv5qF3Kah9ar
AP/ywOjrwoSWAEiaj1/vWtrcXKPMO8c5rfJK6YqXTrziUOpbJNL3sEmL52+1b9xo
JQT9Dzl0jcU/7iphKzjiGUCrKpbJ14Ris2nZekuoMMcr8pka+qFhbGjlOD0Fk8zJ
Rqxu9riS8/rUkjcylJp6AS7fwIwEiuaUAecyVR6UxnJtk38n7KOirdJUzWM05ZLe
n9gO0COPaAIvWiCwdJDilZJLouLKRNm5ps1deZJ7mkOkg5beZloQPANZv+26sxZf
v7T3ZwalU6MQR6OZL60L4+LyE2yapCTJ058iL1igDkGMtcMlOfM7xcw3/7I63NkO
B5wCdqOMkGaXXloP6mLccXaCft4m9VSYp9rukFjMY5S8Qsfo4ot2rfojDPqHSx8J
Q1D8NtjK4SOY03bj/bOzU3/ymxK2p09hPl4CD+nJywMXTiGXAbAeoYBXBT2DnnE3
oHsXUx64G54KM3sBUwWlBLifesQOoED5/YH4tBmg4UId2JsmaP5a9f6tIK4Ffshn
2xIq3NwbgIgX1Ly1lTfaUaf9YIs1LgIebUliRvccv3hzVzgT2oRWga09Zw/nv28d
R1rlSonxMjTCKIErUNQBBnQrU/8joTNBmq3gol/8nwO8l9GRDGSdsyF9E/bOsHzT
+jTQhVNDMjMf65uWB6mhxM6S77FPGA7CGQGfjLKN18GhfchesTSQk37dWg7MItig
dFsoJ0+dyQpES/daM1rT6qcW6Rm9alzo38kDnotmHNsnJTLSUsIAGSAt3ToduBSD
oh7v+vMh1og/1D3LGl8J7DhRhxDc/lAvmNZvj5W+tcqNqfyirnevJ96Dt/cl8N4F
BsjEnFWbt6HONlTPusOQcZOFOcQL7G7YUKFFJv8dmO9gG0lLJ0m6v22gHwHb4ke3
KMRLa4SI0MQA7AJZPAqIMX8QDIQunsUwjN3MEwmzwX9mK/ApjZTX04YeifqGkK0K
19PsQiRTVNi6Z7N0N+G+qC+bfvfnM8R9GqE0wFYBLlzYSmG/h6xbZgEFsbgO1UrB
Fi8jdf8j+kWur/VH60v102jjWXSLDu75HlAGetU93eoRHmNjorK4EJfBRJgaZ1eM
i89Xnu4pqutXtsKGC0cY2BOp7qQg8gsJ0jgBAgKEoerVN8bxgryC1sreFt0FmUSR
b5VsKzKjjP4NrDJ68HFHqmpo57t62ifjlJid5edY1YHXpl/ZmVyuZQYmr3lEAegX
6Gj6EWAmhLMjor53Mv5ep4Gc7hYhQekAQp+lzTNCUllVHuD7iKgMx/XZZM5XvKEU
Q7gCHDBcmQZoIyvZp9ghCXlP9rQ77CC8lG2LlrJfg2wXTRtKyXzhy0yzozCjSwlh
4/y4vxAfgNa+xvrfV8SKzw1MOOxmx/WIC/MvveJ1tKSzFsDlFpGcdJ83aOtPq7fC
mSwVmu2XS1I+jLJ5jFjX7fS2gVPRyitLlJ6yA7B/Q8BknzSlxwipe/sMYL9WQYiX
+JVN3FhA8BV0Juw3eOR8+Cq2SMHO3XqPhYHcxwe3f4lYpgYd2zyncG6iof8gBYcj
lxQn6Sq7cSztBEC1+4aEYowmkw2lQzJ0iaJOaCgOOrI1HZFGRvxxMlbXug6SwL12
Djm/PN7Rwx8y9Id1ZMyRTXY3SsaLISx5BqX0zAtehhaXXB6/C6NgmdwZQXta8E43
wDS9XPxOLBk4X40CwK4Ut6MaEriTYGhJVvHRxcdtWAFp0ecuf0PTFluxYh6xWHbq
xf73Alt9OTX6BmKf73C9GRBOL15TLiB7KWVyGQmuRiQmig1VE4KzsWEHiTx0iXnR
HbmHQQstIlxln+dY+f+OPqzlpD0JdJauXpYoVn6uLSOeOwKTTQZX5bc0xk++VWzN
gzSi4WNtCiyVgazGH2vxqBm63c/dPTKHA/+R7+BWLnZWeqTB0uu/v6d9e8FY1rA6
5z55B+s6tkV1gx4+qJBnwjN0KuD0t11qXPPP6vSgtfD9XvghhnddfdQKhT3jB9Wi
Ta/eJ/98tfAMraSsw6ht6VNiehZX5u80b8bDbKeKw4GF8PizgHceqp9+XDw42ht0
G0ws864NM/UDHZmYekcn1MXREuWo3/Dvx0xS4/ndFjcrEZHxF4O1TuG+U2Z2iz3l
YJkk+yG0baP4rb/8VWK3HUFocWtchqrcihzpvXVqrJUDuor5/7BH/7DJT2svSTDv
PN5ZN1T9Oe5I8X1tDmaEvzIOdPIyU8vIOr3MGP+ukrnlV5DtaNxjdIMZUL3rQNZn
5rDLjrIbKap9S138g0Q2BbKBn/jR3ouXfVhjETWEXzgKyYdg+aX7b+nnN1Y+L/kY
b1B6IlJkQHEnrXPhohF3+v/cl10LtOxIOb+YysnHDRI9qWJAPTwEFg7WpRZ4qbPx
6NqVMMfxnbPozx9vdTmgvPGVZTkcijI0eQbl2a4cT0Vxop7xFVKxI4H2o8DL+FOV
6BdRzt6GfRei0GId/hbZyciGy97MW/FAWYuubcIFf7kH6AZrzkvFrdnxI9jpttrR
OvwLPV74KMIP7mFnUQBp+x71qPUG/Q13bUgTTwDrRu1xf3/NIRPxH/YE/zfntyKw
LG9r0aqG+zBos/SJ4nKSXw9gJMgNCw8xbqGpJx3Rn5f1awrw3RPmWyFK15OHfjKJ
GhzK9CvO5ht648aG2I1IgJjzxBgatxVdFKmn87un0SZ8FDEe57S8HQNPD3YUxa5J
LJiRQMGnTYfSmiSk0fTMAMTWE2XSyJ0B9/Hdh19BuepjqvtnodnV/CF0gR7E1CD9
4ZgzkOmRTYOIHY4tixoBEEp5UYXAsLh1SIZvb+wJNZW5h5Cn0ln6KMd98ABuslHA
rq4BXXlHHi3IcmTK+hfV5glWimPQLjdAnZolRa5Jc0DLI4G/5ggkXnCsdaOJ2Unm
1mu4U0AY91eFOPb6ytdpJTJ99T8IqhBol1ZRVKAwCPeumasgtlYQuc9ruC7xCUWa
dYWtzahJuxSJ5+/YUQhkKAQ6fD//mMgl0YOMB3qkx8/XzjiZ0AqaHOJxLqhwnCeU
MhxOUjdxsoEiJaM3f5HBgR8CeqQGoSSquLt7cSzA2rSKpDZthzbA50roLILU2UB3
I+KtIGpnKneVqzLP3psZ5R8HwzTmF7mlR8cIgfG9mecbwMYu3xcyTrjU5F3hHAM5
xknFSqKd0vo2f0YVQH99LcWx8dsT4qg2tlcjlZ0EU8Zaut4PDxgTcM7RCUTICzcd
vfmypNKtk4dRLg+hG57xYtDmjXT+GagxSS9ra+dkJbBgzhskyxYezd68B98yoxv9
kVMJPb/1TeMSctLSLgRya4BkoCnJN+ljZom7900SiGhjLzlMf7zAn4+PnqyXiF1I
xktBXiMG1zQ5PB1im+qJ7stO2K/WTw6o2SCjORkQjfqwRmKeTLyaKF0GxjiNgaTs
0o5LNZtUOI9fFXoZHb4zxZICVSbNHC45AYGH9yf3nQOjLKujCo9RiHBqjd7le9up
PfsdJqJ0CwndatPhpccHY1saKMsfoeuizNSwKA66YRX0fhmA91PFZi0uQTkt8WSu
dKpCxrcol7JD2fB5Hdof+0eTRdktXjuHMYNq3aVGjQVbucZ+MU3G/ugdt/wcd1JB
C/Gk7kbQ/hq7J5XBEQSfdqwKlZBb9CPYxnNEYUKg7dfsVa4eJe7IySo6yCBhjmFU
BAYlAe/lwCssxStH38xndNnIwecHkRVimCr5OHSq0plsFn513XU+zNsS1GUaCRUo
D7h15y2QIObzXoF/dUUdwIBaJr8K/hhlT6xa2qfUH4roeFsepykaPU/IgbDpcanG
2+Iu3llnOHym/F5Zj2qnJ6G2ls3R57dXmsIh/iLkMkcQWeG3O9AEVJ8d4tgdkFzt
d9SIkMT8M/7E+coHtBbP4tWmd/C/82x+ZAtKpSIC3L9iQ1y3B2ZoO13dp6rxdND5
IKgdZyIl8M8jYpWcx4tgiN2/VwX1DyfuO24qEUWGKcM6VQq6RvulSRzzZ4n1jQou
ijYKeskzj1hSfI+AvZPGiAY9KxUJ40DuwH5wmqElpF/xgiLpOCrAFFcDAG/BxON/
9ViT5EsDpGCLzu2kcRp/epAm66+2g5+vAenrFATo9FYXSZTz4w0ZgnsCJebK9BWH
odgBVHVIVry4Xjd+uFEaB7x9uVAMGvozP1wqla1WH4MhBUw9n328c2IxvolwliC+
0oxopESwZ1Ub4+buEeXeQiDjzqnW8XU0ZP2qdQ7giw/2XRXQ3IrXgCBy3a8p5y3J
cQKX2p0QdQ6wQE0Dom3VkSaQSQehlRxXWhHPcU5Dqf3L0F9oX30cwgq8ECu6Gi9c
ZV5/tjsOQLsuE8ep9crZSySSWjvt6CYyLkrQiEevFhF9vgjxDhA10IaI8b9txZG6
dapSgfLK9mhOrSJcfnhMtDwBcOv+W6sBY4o3fAtR0fSX9QLNnC9a+xtzPT5rSYY/
0hsgsGqVblbXisGMyZd2HGgtFlXkaN3B3g3EWDSyBOIqrjZJDjmkKcEAZI2nieqY
V8SCU1Rp4Ar3g9TE2hBaKJV5iNCrY130ShGXUDquct5FKUjuYEWuvdjYZOLakOFE
j+469n8qelfkdI/JdNn0HUJ4shB4Y3EH55BydXHdA4l62LQcvsXsS2Klarr/qUE0
APAkXcm47iui54INKikHjf+De8zhtjCG2DPZHipdC5B43R0UuBU8R6eIml1oXWxO
3QgYMRyPRMq66g5uSr77vWfy+ao8f8i3b3poxstPq51OQe4eXLyOm1koPdSJ2tAG
ucyuqLrghm13P8OfkYUHhNF7AtiFLs6mCO5fUwilJ5JOgnFww4I1713Wg9isCMyK
ZvWM1ISxwizRbrlJXcxeA5e7BuoRkfeR7+F5/1nrIdesEQhKt9bhzdPZN8ebpRZR
nqEGhTMDWrtidOFhgVZWgDyRidCuCQ7Zzm1w7NpYG01ahGmCyfgtbty5bGdVjHSA
J71CoFHwOrdga3LCiD0pxwFEG60oFLPzxjyq0BTUwmOg09Q5cXuRUMdNF/nkv1bL
gPmtkfebxgVcv5mQ6Lh0r5kvUHmoeO+KJhRPdykYhjoGzFtpJh7Ye+JQpujT016A
orj0E4W+BPH9xhiPcYBgnmJJf2KWaKLhmc1mR6tU73Vlq1j7TTj/6pbUi59wBtM/
6srPvF1wyfTvYcT7o+tjGJ2WGQsW/VrSlDazXaKqLQYpE6nfUlAvlwQ4JLlx9ugR
WaJ/E1SpOPZB0NXo3nYqZc2sn1CplcTMxwPb4K7xQWPv/BA8VRbXtdI0LQWwAJ94
czH7DtuGT0Og2+RFx0k/+CYNO9zMF/IZuCWzkkow2K1w3wkcdMMIeTBLcvKFom+u
0bUI6s2Mt8uwbEl+riD0Cd4/tr48cGlUPWlUwngPFtHNzoRc4Ln1OXmV6gdEiaRR
vujSsCHruRc2PZoFjD6FoQkBVyfxoOu6HgwZCEoow+2K+ouJamB5k8Co9N9R4GCZ
EqexIs7OSItWZvI9zQxq2HDIqs2NdycC0e1LQMCIUgBLa3yJFo6U0V52GCN4JXPJ
kLRezKkUgxH4/UL3cULa9szIxNBqzbFK+b8sS4bXOy3KXNNFV80/aZJa5odV6g2+
V7FYhE63D5bvriGtrtrC85NPExrDmGd4iurZlordkrxcW9D/XXCHanNUDgLHnsHl
NknbCj191wfvZ8JFUDddbrNG1jwaqPrby6MLdBBYLjJzk+McdEFri77www0p0l0l
Xmw0/TnaVPESpzpmSMvQv4qsl+hyErGwv0y/s6HJPvkxnVr6ICy/SRnzfpDs7+Zi
dNSEOkpYJKQu4FhgfHSwKC3odzmZC07w7Ke/Bt+clbhEqKMJ2MDlCDAzk3vBTVzw
rD47pskebMHElceL9sQCvqhYMifSZaJfjB98wat2iJuiqf2/GHBnKtlIxEh/Dy4G
939s/X9hoRSOkJmBNRlsg9JbN5zTK4z9rFiJg2eVx8MxCFl32GwVTHjlBeeYJUOQ
zKiD4svZyM9nVp+HWdBePNlLj+L0/jeGEIwBEL5lS7ZqC8ORey6w9YOvtI1RHS7y
ATUzarqWz4+p4U4OBmKqnwB2EcNtjzoX8i84ILmeeoWGLZ/J9mWHcyJ+VLyg9zLx
Hj0AnNYciRY7rnrDY3jh6eNcyz/1ZDEiHuDe4w6VT0wTUS1f+c5FBOTW1YzIIzbE
UuIXZEjrYDkWjIUqlo0aXCq/pSIG58WW7YQMCcLL96Ya+PvtFwJsOfgzpQJSp2Ag
k4Pq0/02IBPdbtxwpHBC+97BgHFFR27AOsK2dCbAYG2IRSXmIBfI34yrWsXgwPeN
rpyfgjmogJB85ArJOvonJL7nZ9qXocWFMc7RHTNUcnvr0lggOXGHTC5jg7V1eSOT
9ZAfTI+rZb3Bivy9k/PAJ+2CDaxyzUYIayyeEpjZHsC3jlKs5ruF2GC/ARio5uFB
47veXwcCaKmJmLmp96iIdBDRLDeVnWdpojPjp7A9c17+HSK98P9EutQiECCGiOoY
LU8RCC8sDS9XVY/UUwZWOCyMBP1EAudb3xqzOeDLN7Ry12oN15+AXv7+1uXDKPRw
vd70B9s1nJu+Azb3j3xHfXjZbXuku4q6Gj2DUNlkgAbaJIe8rsGKk2uQX/E6kNLy
/ZXMHtzhdgd4FajKV+D/fGMWuBHQtsxG9qjpwqmwTuS/IEU4+LQi5nevDlngLoSn
7WZJNQeRMX7kjynDvLnD4njtblle0z4zGuVEOrJ2hPPx4XH5LUMqrLiDR22n1KmZ
ripAOXZqGxo7ypcuunMmWCwyPnMPU4IdKJSbrHibHdGjuTIEGBSViVluzSdn2wJT
DcH+q+oVe33OT2L1O/0c5rRGKPzWgAYkIt0ZgWTVLSJn+PK+f9ewi0E5HW9xgjlo
D/NZp5bCyAsSwSXQKFOpf5IIS/g+IUZ8pyBOmXaeiP4KAFX8kcoQ7J8JH8K+XSbn
yRI3Nirqojg2L67tbIcEuO2MQC8+ZZGp1SwnyoJncf+DyrzdR/JRrG7GaW0AX0LL
LsD9MgLv1PJTyi5cSn80Y2faJk8Q5D0eJwg6dcoWVBJv8XEvI1uJhErNk53vaaCN
kVuEDlz3LqM8DlVRkKkd8+uqRs8Ka065zmXhNu1PmEOEN2YqoQhF+YtPfZRaner7
oJdGZTuMLhzDrCQ5djjBxVRGEK6C2aIXpCK2XfPeCaqaDjsS3biH9iXxGh2+Udkb
OWWJUX+MBagr8f3P6u4047JJA+hscCElj/geoFU3opPVOyfTl18OoYG4C9vumsQX
U/tUMYHH6fl1QM5GOL7vop0LKX8/CceqKR/n1+gtt0Fw/TF2inyla7cbKE5RJqfQ
wLuX/5n7SgCxi/02nFcldrIqudfLj6+Mk9+H0f0jaVvSv9Je0Fhg/IFk4ne35c1t
WJ+KhQl9qDz1n6WCq5M1/9AeuZxoqRcX7bZ/yf3NlUFKSyewKOfA7Dmk+5ajmKr6
bcEB1Gu5d3hcC90tzxabxX0JCisPSJdh5AYnzFHJ70E+rfzq/Jajf+UqFr6K/Uy/
1pZA2fmaPJQ7E0kLyQAIOE9DAzSZreaVde6JSisuj3+/PHNXZQDwIGnFVc8RmdVB
PsycGYviScW6+S3ifesUQ1mD7QUy+Cm54de0u6wRK1ruoVu/iWx/53l9BleYBfgL
jHrycwfhQeUSkfXPPKRPvHoh3vR7+pYsTXoOw9vw4TPHoLaM5VqRCWv1AXrx/Z9C
iTGexXyoWsNfAAw1J3bnHTi+w7Mvx1/Kh66puKB+z7yKyrML6aGn6jgFSdj2YmGx
qT6Pe6GSxiPw0NAQy6RPKxKY4/lDcBWXbWsg3w9qHkXUdYQLz2l2GyYcL1H1lwmb
eANGOwQ8EawFh6yr0qf40Zn5BAdTr52CGsDVRWTcrsONTOgamAVchJ6/PfdxCj2O
D26miYaDjzN/5DvNmAppzTJ64dMQoIF//7Fi3v+oZAFEVEHJAeMomobjRvCfB34/
9PG52ZsW9t5LtK2k2bjAQALQdSsW7cH3oSAqGGin/uRb5MCAAk/IVhjEXFUkVcHd
LDVvsXXcPH+ulJ7EmnDroDfDWl+1+L4v4Eys8Hw1pfl8oiRB6s02MnvvtVhox3fg
5/dtCUEh81GoiG8J6UD6egOSj/TIc9wtlUYrqOvelBp8/9xwWO5NfxNuk4eJeZ6J
UkS6gP4uEGoSPyw7FG5W1xCaYp3rBZ05z11U5eCzXEY+Ol0wUYoNvoHwrwpclCvs
6CtUXIkVj8a4yDjMYKr9ojEM/9iIqA0qJL2Pr4oUej8Ex7yCCuKeJfoqyfTsCTaI
fII3R4UxIPsSMrgOjsmjYkXEBdAZYrQphHmMtCiMFMEqvFfIcf+DajmnR6V6e7sm
R3zqs9LfPdEoCDHXDQWgEdhvf6veB4eVpntVa3aYHFC7fdWkpA2pTsQYHl6+9AG3
uR0ReYGpYFGPHad54HavvP5LO9yIj6p/BqIoPqyQ3pQKLc/gu4lcAWfwFSGNvMrx
YWKiz4/IlnWo9Vx97gJFfKUu1RdaHrZLLosHhdlgnRP6msI3m3vLzWJlafM7JBQ5
iMnT/F6nvw83wwk4/EQ3RRQvRWY/NPiEwJ1pofwu3DpYWBwjRiQWLR4JZczwfXBv
/HnH1battS13i4WRzQ2HcBDMhZLgpv8yI83m5ApNQVFveSQkWsAAnFTzk/Ool87f
DfKRhjjeX9xTq2dCV1K8Y0WmxR5l5qCKLF82Z+FKt5HKNP/PVHdXWknIGsQ0KNnG
W3Vz1RkIt7lAqmSdkkMsiNcq/dgFNtt7jeBes0w3ZDl9NETDMIZYg7bEQr0zGK5s
vYv7ZIy7GuAWkhsTSXCaGCy4LsqKK9FBijYfHm+VDSCt3yVl0t/4heb4wZ7wxQwK
VDFSBC1SjRnRqw/lDMOM98QPW72FQfiLgb3uBTUfQkaDy+J6O8wBPm/4TuVVdL62
Z9yX4hyZJlgpbqeqM3wAzubfem1vNK384SVp/HkLY8sHND65ApJEFHWJvXBu4T5K
dFY9IDdhE9je42P5xM5LT4jp9D8pB01K/4nORj7LDc3C0lWRgRufHQHQFLNacgvc
LOAhG0SpusgpnHIoDiGk2fJ9JT7if2LkPRuFL4Vdsv1xzsdSBvcLuiNPCJbTYv3i
jRmriWkm0yOXTWxVUa+AbDxKW3T01InDXcc+7RukdfZDzCTCj4kqIgN0vz49Oail
GiFTR8nWrHE1bDAY3a8zmwWziNeC9+68Br8Us0FyLZXSCuynJ46ye4Uxz0C4rV9K
PTYRP5MvresWhHN5fJkno6/PVh2bziyoYo41i69R68tqRL1WY2XZe6pr6/552riA
HiFJjMF9YoAkj8boZIqqoyN6aRCQP2kdKy6RISDVliVT316nfjzURdgSmHSBsekT
pSXYOhmYiwbLnIX739oSc23Bn3tT5UEreRu3lNs2/C0XeePyYBlR8/HsMAhA+h4/
aZMCCbiMENtRZn5kAdUW39ztiA3q5joeGLZ7DSKa6+blr6eYlIGzQSxlmdo1U7Td
qizLkFXLpzPzWMRidjiZpSyNS2l6Kzv725r+Cus4OF61CMY/09btfhyqRrsdXAD3
undFoWP6fO6cXklc+9yvltmeKFpQhGp9FcVmsH8HhXUN/gkR3zodKCea22xqgY6/
FQrsyU+f6KEdS3z6mNqtMk7q1/XUKJivNDD5UQENATSY9Hl/O6rIGmj0GRnpsXef
PMosWkX9SEexNRVKIVNzkWsQmKdbKZM6UU4HH5A7UO4m29YRAWecRbsuV+KAVESk
/puhYnmXNnLWW23VU/qu0EsrCAf9uzjILSS9AY9Z3gyqnX84QPy2NJHVXfzHADCd
HCGmYnk/ZlHQYML8s27tuHKRR2hHiXqPxiSFlQ/R2iRbwdbFJAK05a2+QCXcUf2v
eQJ0jTgrBewmy5fNpiGmUVbJP1OmzhkPQSMRbjw1bXTVK1tINrH248Xds+GmYgw7
aWGcVD+XuIQ9/rwoNVsrE3fT43DEygNGq9ItvtnpA+WNx1i5ZfsdOtXU+LfZgDtO
EidSXLbNPgl+Zh9iSszoQD69pV9KJ4XSRg+T0XqharD7NG9yDjRfAnzgYymO9WuP
1blBbE7nYINbCEJfEkn++ibqI5p/lDbq5SG2VB1d/WHVONP99ddtjfh/dV4UbKWV
b3KhvQThTKog5hfxsswEx/e/BwaJYJ3I3scmvLRZ+NSR9SrCahRoR1YStGDlBF/V
Sw/k6yEhrbgrliagrTMRCUqkWBEhzUhnr0j1ezT5OUfT3Qn5/sutl+QarJyHEGS8
MIov4HMDmypO4FxSi6SW8J7UBzq92gRgNMuzadiDDurtlZ0C4gzjf2y7exA16QjG
BhWe5va5yBMR8CvBEuPf7vIkAZdAjZe3voJmFSAh8jRhjuPBgQC9VefNd3Oq64cm
D21y+JsnjcfBP8Z+1t/MgDYdGC2/C3HRp5qohkl00khLQBy/2Ta40ryBW0EAzClh
bOjSI9ObQ+HSCQ4EDwSxrZY4c+n7Q0juEleNhypg4qZ2KqSK9v+MrpYLc6Pg4k/b
xan4E/aG3/CpQyV+RP+HXTpOHQJwssBD2ktGhmN5Phvpjx4triQlQKUV2TXK0W/h
5KBVOZVFKUW6ls1Ffe+/B4F9Zyfl9nS3xF0qgJyViZiLM8pEHObd5hUxLJJfvQVw
qKN3N0vXcLVMWL/gz5DizBB0J4z7ooHOIojHUxCmOwUXvJEhgCZEja3BqK+cfUmV
xapLUPV8A25lFnVMXOscv3YsN/bMQ5aDHKtCiM738KdIB4RFEAcleISrwlQcinLu
qa8aSnAm1Q9elI34cKuuAA+GH++cjXO2l9mIkjPkGLwCDN48PbXw87/XVpLZpsEd
qyKfaF/FCUdH/vv7CFfPv/2xeKvkfVO0NBM9NDMZmmvXNiXLmno+KupvlCzYNVKb
uJrsol2ZVKPe/4aItMgwUE66z8mO/WfiW+X/V8hVe4pSp7lLUWrI8FerpNO9hejh
rS1iCaaH3/BDVpSlke5DLKBL9NdtO2+RYy1zUwOqRzkg591TU70hZPib+GzA2I9q
UvJT1/eZ3AFYAo4wBmoKGf5AmAtEvLVSEliyIB8OCahjlPrXOtKAtVQ5m0cZJYOw
hS0lNmBaPX0/PZpG/AakMaw8ErMRgom7HFGGJBPjaDfkAvADylngze0tlF0CK2yO
n4OMLVWnMbb5MWHUq1ztDdnAtwOZgWbLnZ7K3GL2oqyWBjZDqOCZqDJ4JL0HEK6C
ZyBVLMKX2DXkyFs5uWKPWHp1/taIDVyjq6acZ4JbOJeMxrfhCUQf9uAGA1KHd6SH
/V9Op2n5DB6p2L0/fHsm6UKdRz2eSiMyxJI97cK441PCIhEFeVsQNgsPS4fr08UC
/mat8zhAOUOoAD1DfUTRx1KTfgszpjL5Mg0avcp26mW9cfdM+0WnGU6oEJHiG3re
pFGcB3O9Vh3lJsC5Ze2K92Y12fwV/kH0BqopunppsKMgSexieIfD9OjkPoG2zUDj
4CMbD0tY8D975Thhxi2pAxvT+K+NhkcToE0QjAM7MZF6XBG8jrq5DffdTd1+NN25
+NzaGFL979XErsXQejxmMr+uwBSOLsGunXoqKBmO62tpGfQtFCqryQnHjmydUKY3
LMAPEH3VoQhgLe26Vk/GprTKUBYKV2/hmzOr+jUgJEgZfVygVHgJBUih/TRw3TPD
E/W66F4OEV6BzdCTLQoZX5WrzYryJrsJtdgTX2g72mGwSE9HfI7ANzefLRI/Mk1R
sT7iob7CDSiUopHwJb001Z4acAqhS8LqV6vqHsUupnGvrv8WeUAjHFzDZL3ngkAl
q6yIWKwzCK0gCNoFLRzZywLQR1JmasNf56x1nEE33A+4STtccU9ZFbcMLRqRvyV7
vX8aH5Jculnz7GTYOBEHh33/QlU+yXlx2qVtSRUyTyyHgYjYtHC2tu+a/A6VLpVY
M81pZwszYGT2GkWbGILon+0kj3epP2CGa6X7FQIK/28etyUACqvNaRKBXt6JplfE
ejQM6ROOYKVVojrIoVT0PC1pTQP38xYiLPp/TiyoEE/5UGymzTtNeG6Il12rvTko
T7bSf2Jl+FLyt5u25falrKN+oEKR2CHgBJJK01T0qgA/8UVPlIunsHDs6AgWMLlH
vFNi8e6NEw+sl0e64PQgunCMwkqiy/hjUaSFLdnFkTHgNK1WT/GmIIokfC5OuD2B
DQkTLaAMTi2VRtG2mlYWFN3r7/5GH3UgyfbLLywlugFsjKaII9DHHuWh9ic31ZMj
wf5QwWUQFTHA/jtR3bypcqpWnsRzskb28QRUAlwcxKZYEnj4MmJxxuUPN0JDDMmC
zbxQ5P1oeobCQhspiCGUUQM3VwYRbGaJzGY6T39buQR256Z98f2E7DI8G7SAcUDr
Qkx/DfSTjjAQ9A/YULLTLADKH26xwtMTqJ0aW8kIxkkUMtyZAlv3q0tmr98EEYZH
hvWPH3A3M5VtC3FEp5hwXojN0sBiSR4OHNAEbmJiPzgIKNMFpG/qpwxWFH5PM/Ee
tXIONyehv2CHHrVqNlebDZQvX+epEOhVZU+y3L0coNqA2kqWxNORazAEbjcQaNwy
CA1fdB6RKaaQlzw37BbhIvCKgS37Dj35v76EbceTgb3M0k4ResPL0nr+7IqRUvll
sRi1G0UTOXjinhTeFYm34LlKesRg2OQFthg4PABU4wGOevK2lXoOpNfpQppcJ2nh
t8YiQzNOzJY4mRF7KzAOKdlGE8yfT9vML5sT9v+xH9W+ClEG0yy5jOU5iFG8L8CH
moO5zB2iBejjwvovJ053X9fgBHO3HipxJKTBhZnrsUr4+BpqysmkU5CejiQ7nDcW
ORAytxfvpDweYu1RxkDdP8NGkzs8uCwdBnsfSHdSGIy30rmR2SWckNJpTH9wJPpx
PWsKrrd2Hph1PFyf+hYNxTSNbRciD9WC4n+49D4HARtwuTPIcSUyrjKxUX3vu+bh
LWQYPG9vBp6+QX7h24tikEtTcvXEhyfvOLhRsF9qHEFv7LlGpmA9Ke86haWo+DIX
s/7z0juAQT5c3aapD/Ed2WoK/mJ5/iu1UehEAoeCwoI0S8CQU81xKayiPXg8ED0K
H4QeELJ+yj9a9R7ESuTQqNB8z0YWhdrOFGQCCnWwvakx2N0j09Y4BB5kwLhWKfgt
G5jiTRHsbhvED7OEFZjTgANX5kr9Kv/+5M++JBuOm1Hm7lLo9OfXDZGc0o5nJzX0
iP3YxUzKoPjXHpcxOGR8SNECYp2XOIBLFVE5RXCxdBFqI2oLLg9Jz2//IO1V9FAr
kIsB18faed7B86pY/3L/KN2iwV2iZMkGapNrGp+6e0bnUxPBylcjqjlMAR+CG65O
w9m2FKRxKrnaNUSBkcRAlCmSHhKQ+3nNcFTM849NDd6tHIQZUK4q+rz9FfYMSWcy
HazooLNcKzYq+hChkBjsUFQoEtluqh4xkwv8mLKsSMWGEcUZxZ9MbAfjVXOKSsCF
YaLedngPKPrxMl36l7VV35HiQyhebc3kCzg6hWLyGUHaUaD0iTKM0ZwRsVFEfBJ6
0TSTTwkGDIOJyhdpq3YbgKU/MdHRZJwgs6i3seUgfh0qC4pv9fLDmk3iUgc/U5Ao
dhT6ZVJZZ44vHA+kwQ23bmZQWUEktznvzt36KDjZltdxXgs08Q798VTM0M3iFHQF
01qq4/3IAtA3ypitgQucmX+ctoLGdelTHAJls9Cdpr1fT/esMEd1jy0zSAvpfkuF
lE3J9p6asY+s0R3vdYBanSNCzw0nLywtRBQ4MP5gseF8JIS8ZvfVyApvNMUkfLy2
piS858a1KswuyX7UU1Lqjcm00B/f/GqoG+iE+AyOKx+dmwbH8WP1iKPFCYljq01A
goZhf2tHLqqfDU3Hlxc2T/k6AT1s8x8fx98PlXrkOT6lDba2BMlyFRGXumXarnN0
pMXvxc0VMFv1qyK0HFKdmE6XQ/P/B66urIB+T3ee9OM/qLELoWsSVUECKaOs//T5
RvNBBod/d+X8AEx6koU2n3LbMgxbMuduxBzNABveiR6/OXISuQZECxK1DfA7edAB
xN2RCcP1+UyUBFRBYSU8plgF/zL7DoM7dFlSJy0/iOWlggqdU579jLCGho2PHm+P
+X9XsGWSPoU14x0kdVbfyRL1GkaEb0udlXa4EINaFEH/yn3zYIzm/WCWbuD4s8kH
zvY4oO9isXS6j+1cxygkSmGarJg5px2AxCXv67ha1Wv3Sg2zbeFl42x9nFfgxWAa
WPpHbp1+ciAaVpfs2K4oq3HkLDJlI5e0nXnn3Hk8BJna12gNwbV0unYRAHnNsyA1
u7Mb6uzcJjG4C2eX8qIivKvreDrMRlZqh471bvyyUDUy6RNoju1g7YgKaSBUE4TA
bMJOY36TfbAbUQ97T+YzpNuOrcQ4oCaUiFe532NMbqC+4c3ACBVkeZjmJLOwaCxo
tPZdU55jBQ2jyQsavaQJZPduv8Eb7y7USwwb5UhAADsi8tMRNxtpZyinmziox+kD
lNAhX5NfAJnoGb7q8i4LMK6/hFE2jOzz68ccbIOwaXFaFoAgzDYAgXA1GLukwvbO
LHFrnifA8ezbGkxDTsZcWuzLSdBRfxpHIaE1apuDuYa+XQbutR22UyAayLMa9cSn
usUyL1BMs3JghvR2AkxEQpQGt41AxhyOnKerJl19tdUVVaBjuFPKu6QZs//e9o1t
nd1PGXeoklQ+JyGH/3yeKM2rZRhASqIHfeuNFrtB/ERvEf+oArWocRFRIAq7UXSo
ezOB884YBIz1xGWjP2TpIevTl6daNV6YcgYfrkc9GVVxbLnB2F/4v/cPiOXNUZpF
0VgOBjOzX97NjKDY+mXTlhjE5enNeJxBa+X1XUf/wkrOMllUBxOSU64kL7kzSiQW
jhuI5w4vIPvzxkO6srzkMcUsGpb8nv3ob5v0LZdjmSVYFlgCvF5cB/QEs0Vwj+Hn
nxVqd6hr4eFA4e93VnahXcE4kLcSDv4oE0p8xqxuXJlZv9UsDisI9QriNsozVZon
Q7HPJhWjvVjWNNQ1IZekRfCPBqZxn9pmQkFvhFUv2r63n3BAxCDDNh4OHEgG+Jhn
J7Yk6LLaKVHb6Q7zKr3LUQyycKdyetE6Qz9pzkNBmJudcPW0NvewfgZ33xUiHJBT
0CfjG0oNNoNZBYkcaCD2cqi6hjntNL+zRvVQPErzXsMLtLuMxgAKVlo62hXAFO13
BeiN2qBxVPPRwMNBlQl3/9+8FC7SwMh6eMKQcItIob74GD7D1gSTKBiyf+eiaoUq
vpoPWFx8G/5DXm2ZOlFtvUSquXKROEfovslUQBSRV597k0BIKI56ezjRRrxyflf3
gMZ5MKxa6FG+oKhNlPZIgADo8mTJUvw9+O6ylsFOdcnFA7rv5fbk7b7eNnqbsRD0
QOTojVG5NwDM+JNtFpVj13A2QVEw5tNCnmiGt4xDr2LFXhfAA8GFuaVfcjSUygA6
vMPS19TOf0Kttea0kxHgho6kVs+mmGf3RfPWd+w3VJRdweQbP69UdQSdfR+fedj/
BfO8WOUAy5kXpTvGGtsAYymM3mTzULeMPjImhk2gRVYgMSJHRpkdAAVx4mHd3EE4
c1WpdLSmSvTc22ICE4UbDKihk5fieAFkcLSkv+64INkSPvhcRZlY/dE/r8hW6Su8
+RLuKlzc6Z8BkIWgd1/h0V9LZ2g27AvHGM9VWHjoasIXdndD4OhBGb047+AkoAGd
yp8EPv9myJdz64001Bsa1TQCYcQGz5Mv08QNsjpqSzrJo6bLXxMBl51mAHdFDLsy
lCtjsqyoQzJBtqMcPRSyuDlB44zlQoteh4Swi5RnRY/DIv7W08QASYFBl71/02No
fvwojC8rgTWUPomeQqoN3qIXtiiy8bUWVb6xtCsSOsETisllHyQ3xZGdRpH8HOrL
19Ln06ArIY0/Hm6qcBjrZuezsXlfiadADE6I3m27ei1wdPQLEOGzr9+GxuJf7rld
WucCpooYEF1r1cFHwfragnNSOtV+XbRk8JuWG3lelT6wa4oaX8hlvHqpIL//YC8j
bhl2uq45wBO96hphsaRXo+yWexE4K72g/EoEZEr8DVu377uvZdrvmf++aEbaLQ+r
w38HqWCcIcCb6RB853H0NVl1dyeIMhmFp6h8wuDuCRWaLrvMyKwBpo6wbZlkD5Yg
PY9+SyBAWYdF3GBNsdtSrVhb7zjbNBkQKoLaS7z2jwoZvWOm4JJ0QWLMqGP+8hlB
to2MlINMA5xTgqbHr1/FvRMRNmbVhXDqj6oJvwAk1L4TzclLAzW/onhiDzDy5g/3
71aiN/iIGwq1FGUoHf3Y9RLeSl4dJct83nA+yLq0434O3i6m0Fq1xuzGiw+1bmyI
sboRx7pgjRXBMyl6JNQYPgEJ14rxATtwxD3H1qhAlNaRoGQlrdKC+fpR4dEiE4Hk
P0jET3tkWcgQ7pkW2CEA3GMUHQmayzrlkeDeAok2rd17lzrtTMelY3NxZI82KwEI
IqQZ3+xQMvO0VweI39XX8hUbOsYdx+Eh9NlJo7nFxYBsc8VFKHTGjncY/fszNIPS
dGUFlZhtTHHgQcY1Ln9FEVmnzf8LPafaVhIB/9gUiUe9K/Ro8Lr9QZQfGdrYuubM
d67lDLwhTjCXn2Jh9M85ZM4CzA6wZDrCGLqCSaeG24q7aG3o7Vkrw334m5+LxqT0
aEHAoayw9bPwDcF7R1sKlqLTCchijooizsfwWvRtwdQ8Zm14IUwl7F5xtiRvINA1
jaXjdlP5Zz8hjh4M+wi8SMZQRUpSI9JfeOdi/+pHXv1TA5Xy9/mQrPIELR2/e/ff
yNpODcImamS4Zy2k9waRee19IqAwiPmRh/YQaEayx6rnUXpb45yqOZ4fWCVCWr5s
DJgREB4r80OgbsGE7Zt5/GQddTW2Cj9CiOFGb1IjRXPDuSb+vbAZerrzcSjWBqHc
RYkZAlC1AziQpyoaTSSms1gulaXI8IPIX8LxPKdK3PHQgNkqTmcgHl10KChDg160
D/x3/ecrp87MWrKh/yB+2IQ2SwuNWUXvBOTocthwH9xSjfkNYj0KKwzk81A17888
WL6tuhc/FE/VNTVWy2mokCAvB7mTGq2vTsg7bzi9yh51aqOjsm/oF2J9jT4/cD7l
qZAayh5IJ/l9YF837fkMiTmYSGu0rdMQtrN/XvtFTQ5R+RIzcskM2cuxkyvljaZ1
RWjC95FKb+iD2yqLjPwJj46bN4avlHs57PTLOIvZ68U5L+Y0qmc85WL474zA2/0/
paH2wGxM5g1aSffKHLnwFmWiCvx9nfljkGBUMgnrj8ZlqsykWk5gQXLRE0l5YnCF
qu/WA0Musc7/sfahKOa+OjwdLyAgfQ8o1TmpXGGUfu0hqKiKirJ4s5laCOPgYVev
2PEMWEVt5sx70adxY3xFWe0wMEG9kCX0gCa53j0ELxhWywAzArAyawMecUi8fS6C
20G55aaB4pIfJJvXYQwLoB+HpoAwVIEe7TOWlS57SqTjayagxFHYzOwgYlbvF4s2
tKOMxRuNWmpAPDU8pQAhDlm8uueugPBxTR80a7ornMbwqeX3AlKbEDzOVuxdo71J
u5ujjwdK/wDjAyrniLJlQqgQsO+t6bUUEDgTz79IkUK5spJvS4TaxvwdET1F/EeB
Mpw1ma1kbstzNBwTpKayTeN4oShb46MtYX42GKe5zkA999sG9iWgNic8KT2a/Ma/
iceCcFQ6PRuxUakYMbQJAJes/OnR3z9ymOXmkFb62avCQBH4xdoPOdixCLa0kdhQ
8ANQ7vVnTRLGrrEYV+eBdc3xYxjA+0YusM3ZbdCyWWQULgOlYBTQJJ+XJfJtVwz3
vbScAQYOxNXPeRuB4VOYSByKpnU8WGzrSwnW5HbS3SLPyP9WSYZfkQIfRbDqqxt7
gNRAWO9EUv+AzmqZFMbBAU6iZGi8B8ZNH2ze1NyeZSlDqhxHYfxOlx1UnYrezred
eGZv0SC5Vnzpo+kWuitmTk7XeWmEqYRyeqK/nGYL7UjT14Q9rZuYzBPrJUCADgzr
ES4SFtE6O8BGGecxztDnZB4WTcPYZUutRE8i4zClPbzYtQTUuVe/dVOjYR4HN8Bv
s5FjSluowgkngndnQtcA1GLZTrWjcOpjdSR3RGJkXI4Sn7Er5hxEbe3XcktrKpY1
7By1xzQcrrTy2SwTp9+F1Sw4G+wO5wnE5RdO0nxXa+76Ugqj271Ac2I1Na8FZFd0
RxLWnzloQHdkYcKzDsfYX/2y0kI1UoYEAoWPsfgs6ucs58F/PDkbih+lwc8MJjeS
th/ODIc6oT3uYz7/EXXlhrEdgio4l7IM4zhiJOOO4rI0+xrKzM4RwaU/sI9Boq0y
Y669MMzfVRfA5IblTZ5ARYeu7Z70QFTEW7T5Cdik4xGXcfMqfZUg/JdB+k0TBJu9
NrNgxTOGkQwI7W8bMQaDaJBjrffqJtbGXvr9GX+lYyAESyB3gQ/RHmG8SdnHRYbd
DaX0Whs/XAFHptUmprM/wstwBmGjISzBrIiBNSPAbPGVuGhqwkPkuwvfhDX+aET/
PMo4kvz7aoRSoSBGMOLtSJ3LU5ecwSD4Z48hbWJJJ8TAxVkpYN+Rj8qJWFWK6Kdm
j4sS6HolOzICM7kt83tTnZtuPP5SbgJ09/f24wXNCozKGpuhePvMDxJeCg4SaliB
bUrgB9gGjLa52qsopmCGV3VVCMyeafvhrmZ/aEppu1zUMjRumiLau/RzXz6PCOTz
4ueINpZUmdzku/NEOk18OGPI4uiD3+9MugiZ4RVNUVH+N9V4IHXlh9VU5YzYPi+3
OmTrn0DMmFhnrY288S7euoCsQuYFrheHJz5jv5vvB8h2T0jCZzY/9I0N9w3OoleE
1hv6XlpiHgfdaOGqsHrd3uuPwdZuTgt+fEz3kuCDzl3P6x5s5xv3EMLq0+hSjpEj
7ofrxANqZ4VZiSFzOEC9PHF1uA4DoKRCBBr97r5IjZ0ZZ8wZAAgHcDhEPVYq0oTH
eDEYDip0DlOP7yctVSVYroVMJaZqCJj3bkjlY62hZFfSSoYvCdtX/X8VbkN2zY6P
Z7HYd4v2bVFOyBG928/lhuYfASnhxUERDuST4TH6xUNOtNh59aS/duPsJwmoGFJ/
VnK5Eem8t1HTSAXx/IHykvTef8QV+E7ypLPkXA/SuA4KGiXgVCHERFHp3VQetnh7
fyFgH06ddcSJI++PiC5gpBl21i+Pj5vm777kUZjg72MbXBbJDCFuhhgquOkVsV5o
uopCXHkhKTEwZ1UVeP6QNjz+a8gKWXJO0nyeubbPCVisAlJIWpkFO0cA0IRMygHJ
FiGvGcRyiPSrZ0IFw1UMwWE7JHcoEOayR4BgX4TftNsv00njqSesm6owm4Jzhyav
I6O+BTlTkFiCjO07yzRDiD191wdhqhbOE5iePdmGShvpdWo8WydtLYP0XdQ5hndp
l0CXd2bNeZje/7q9gETjmE2zKdoQs9uQ5n1ZAY7RDMLI+8mtbxI/WtMvUjJra/yU
jAyk9CJYdar/FAhcit+AWuqissNJS6FWwX7tm+YvJ3SyNoRjY6oyA2v3or0tOMAo
LEGpo4Rv0uxVyar1oevY3SDTkhZyXf23A2BqwH/l267DxKfUQ8iCuRvrrTpAdgKX
BwVeFvxIltDLxM2PriWTuhojtC2CS0yhHMGDPeV9BumAYzABeGN1GfyiUmFrGV9w
miXcXASYIUS5JquD+T2HbcO++LqntYebIFR7for+AWKSz91u7DlXk161hMue7qu/
D6eJsFy8t1REFbI5ZuTqGj7zj+7YgFOHvZ9LEuLwSaY78q4mlxXLV+p2cGypnIN0
AUv8g3t22hBAis0NAq69FVC7c3GDOWn4yKB/bWD7c8WKR4+R3KkBzSKI1am+QzYu
KwZX2psT7XoAnH+i1GLPlTf3bPrg3IygbAxfplf6HajEk+v5cM7TAfKSUu3Caq0g
AcgJv8dRjJojy5WhUGQVwOFyMBvzX63pBVe/Umx1BI9qNbt8hkxuFDzd0qX4tJFq
v5gUUDXQBsexA+6lDtfcvAaoejDBLX+QKRat8SLYj20RkvS7jkMcAFOWpRVZJEOr
VIJCT8e7+68OqD5bSRL10q6wxpfgo5wLPe/CyRY9eHLrHszb+RIDXFvK8eJVSxsb
dKWerLyH5/kIxMukU76ZsbbbjxtHO67jGRIHxHOX2xtY5ps+XIydwlF0mZHZetXP
EWrRuFz55TUKD2M482JHXzS1oSLKdUP7lEuVQuw3peeYCkJYfvkYa6Cok+dJ3k5M
6Pk1IYDsE4/cBi7SaAWz2tKFz+D8wM1Fr0FvpbrxYfd8FP0Dd3fuo4eEAgoXfY2J
aGPx8cieVfAaS9LcCCeF8yw79Ml/lPMD0+hsovJxST4zYBXYF5Ofb7j7XgwwPbj7
P0swHg6yy3yyvWUlMDiBtQZFFkRMfzX8ffHUG/jd2Z8Y4ztusGq9WI36mTEPpoEq
aRQjrArcw6YIFiwHmx5MAuVxyuPPDBdxROiD2gpWy10QxenhOTGiGkO+be9grur5
deTT1FWuEIRJ3Kh1xzgw7km5+QPic+gVB5O8W8HqxA14GtcMstMbK3J/Y0LVNU09
WFIAe3ywh55qfTRIqFXnHcp2PdpzWfI+lhR2Hoqsz3KLvGNG7jkdislIcXdD1QkP
HV9Cr1F32YIJa1KEX0yjIStGqXHJwS+MfTj3MfH9ubJzzRtGjUKVcmkI2w9lY/PN
TfqvizVuLdGlYxKFAjQK/MLnp1mdFFRzOyMtYyhJyeF5267FFFhDmVGRiTUa76XG
2AYZ8PmgsWTekJkPZmfbnLwBf1f2StzRWeVeROHx/N9aacREi8ykEsOTb4jtvfF4
Dowgkh0Q/HiGMavfRqBm3UGyhveovGCzk+LU7Zp5tmj9PdkX4Q1n3gC7yAZlvAnS
JhaRXpxU6UYEvWvmG2n1VN333unIRhLytkSX40zqM3SUMcqetyIbPPd45Gt7N8mX
JRQc+V+KaMKbkbOmcfXHRZweT2pnjw77dvVdG1YINF/EWcbkrv+SWOUSkjE0Vtwo
xpQbC7dtY/2zVKt8E5AGVszLhjfKq5cr5k5+7NFbNMnaos90N244a2j+N0qOFhnz
l9LOLHS4LqqczzlBwleUnc9jXvwaEN+JBEH0jRVVXFkb4We/Z9Wz9mkBYfQ1FfFu
xUmqpurPsd0Ae96/KBgV+Y5Gv54BrJSgME39XzZu7RDFHezuU6jOZ5Hk3FZvq6w8
UXDdu7AUDx7LO4hSJioVAhBtDtuEA1eOvbrRaRsEWCLylB8c9/hE3BLjCJzn3Dyj
5BJGrEL/rqa3+DT1k5HXHQkOZTotPAMYMVmX0OI95jNlH3vtqG5y338pwkdelDm6
+4lfm6QyDSLtIsVodI+NWk1Bj9WGg2NQIDrGcDIdc5tm8HMGfPBMNqixT5a5MnLz
HlWsRgFNYSke3y/Cbt+qmdLkSzlx+iSYPxiIQ2bU/5d2nxibZCgD3IYwj+1sgoZ2
9gHt2L7QCArY8HFVrYe5rbghBPSBD+mcPqgk0C14dxinr5KaedKTvtBpWtJnS+NF
UR26wZ+HZV3MNdhKfDEyA1+cmCYCSxzC07CFXBXCZK2trF3NNTsSWiZSeWf5lfz9
yNmD1SxvmF3cU3xjh0Go55BCsvC4wOU04GxICZV5aMHsZw8Y6rMACPHiJgrTLvNl
NtHZO9zLvF/ocuRluTElc3LNYDq48bfuT9j19huZxLJKLDyroIXFRPKa7hseQpmF
/EP5OyqUgBlPPkL2/1+BAYruxLqrAW1Dpv/+r6jSVorgCb8ogLCRCcSU/GZtoBRk
K7gVc/WeD6GYBHvT7KpiUQcCS2cxB8ThQ6as4FkPWIKYkOeW4Tp6l/6PLo2di2mL
iZ+QeAbGM8ug52CDLNe9aYC6KObZvK6a+NA7glwW/rCtmiK0IaNzA/8t9VB6o+Sd
crezLkmZfOMba9ve67+IuoYCVet8mzrFABKTUpBiQfvPUvO002OkFDgBaa7u+uRc
ItXr6Qr4rf3RAe25oCzXNAqlw7RL0qXtDiAZ05NI8i0bbBIca7oV0JAwhieAkP0u
p8SsX8Jd0Sru0TRYHlR6ZTNN+BJ+zFMeuXplXsLAVciobeSCz+4Y33HFa4XR2EIt
ZpVvIZ04dP+bhf3eHuM4XL72JWhwgQ5udfXLWLhapQyhrfIZaGgcxRtfxIDe6e3b
dN/ntsgqMdiXeM1xHszf/n/ZKhonI4k0nqT1/JT3rMPK7JCUcVW5pSRbp8SLSs2o
a0XN+hrizA/1jDBsGo1SmS+VvdXIcQscNWtixWgv5NlqFJ+G2uSWAZpyZQpqB0cO
8ZcrGEuO99zdCBuDWKvDY75xMHep4RgUIC7KarJ1u2HT5q/4X/YzKNDairWQd5XX
22O1dxL685xLjd55aKHDyihUrtMkDurS3x22AajtR2IvA8UwRJ25RxdK8Ox7DYBC
WvvzNhFkhcznC4y/fwo9QCfRN494Ct6TAeRuhDwCAKngw0GcJbcTy66858Br0Fda
MN7uFtRBQ8pBxPb5Z3vNmmUS5ZYn6KrjnQZSMZZ5Cg0FXc0vtbKi5buRrH5IBrfL
sqBaLszN2iHpqE5P3PZCcWBMTaWsv/wBiU4FFV9ZJL1h5bhvCFg2NfvC8VuR1aef
kaSXneb0ecJB/yrWCtzcpqquN/3hbgTyM8qWHFKjdHhN7QvvGJB68FsO9M4ihzQA
jLRx8Jx67tlz71fu+SlJW8r6N7TnIh0Kmt3nUhNYMGqusOSfVTjS+X1J6el14zav
ybVyvVIuc8xDcKS95idGVwtg4ifPrGjTdoIXs1AWHnmzi3nh5KDxkVY4g8aSLqOY
wGPO0QlLCE4zS+kMaCl0niItSXnrTajuTwuze7e2r07X8O1/BxSLZwfR2LsIQy0O
eRj/O2exHPt8yiDEaFAHf7eZcCrCLkSlEGbImRINqjZB7HhiYmr7mO5/6d5vGrUB
zqWhZDtPVf3zmdVAHImEegZPfeN5Zo7r1gjvxpNKTm3QYCYWrwoq6mTDIhHKiN+B
n/ik7wo9nhG8aUKFec7yasUFQwgthzkfqx2RdlNhsY5hkje6WaHq9s2Q+yvpUVBY
KxxEXikIqk6ZyyoSAqPE2Gnzp79o0POTSSUEpPXz73vqbqr8GTrhx537oxacifa0
ZmD6NlHAStMEtUUDJvtvp4luprKqGKt/5lcPdbeDMg4RNwa77ncIkRzV3BaFJRAP
rBClZuEzJZhKVeEg/V3w7GLld9RkmpsLXB+92L89WpsSRbNeoFsLAP6hb8d1SBYn
ZBQ47pgoDu9bzidou3+iDdyHOtpRxLje281/LebBIC46C3omtIBJwTZL0lsTrmm6
yUua6HvYuF3vsurj6UZxUTg7BOR5cXKCgdDWeXdDh4RkmkD8YLxGyoYv4+gHxmBV
QYTG32kZw9/GynyfRAvotmeXJ8g3gqg4+N8pTMmBciUNDKSwHrLLQzFISOZV7vEl
v9s103kePk2XEPO1xaX2pFkw8py++L3IASeMQa/wBwdBOa+KzkgcLwnZloTMy2X7
lUTSimuo5gSYf9srGiJxqY8KFmVld/zZ6umvWKtW9Ebk+p/YZK5syHpBCWQf1V6X
s6AWvdkRWwVe7vhvTle/X1lO1a743EwV1q7MJMvjSAlpUhFzxEk64hkC/KUMuPos
UCpmrS6IZbglAyB2j+VOyYXVHL5wQJxoidx9F1eMNm4vFMgvv8ud4w22J/gaRq4N
XiZzh5ZWprGdf3DEDZJmPVvjFaujhTcXLRwWEeF9LpvIC2m1vWyGCPsScH5pxmh+
M6V7szBLwIR1DRii3e8+rzt0J3jQclc4Bk9qs1nvNn12V66ID14c757YqhbqaCrX
guaNf2EO7RDmcLDTKhNL1c/BpklFO4tWHkzayy7GzyffYjRgRCofSFw82bks4Eew
AL0GsBHqguWed6NwAfvCNxcW6quuBAWLKyc84kHJVNvrQ5IldQrHwfKc/hT2xNxx
XBicgHHvs3v0NSO/K9zAEee9JcvNn13CLUnYGLqn4AQw4HbhyElExP6iN8TEsqwe
qnPI0NKEUTHZEFBD/6HDG2ke/VitCXAsLF/As1xAiM9AP5urvYOp12FKj0d9oFQX
9J0sf18KuZS51T0Sj5NC/q0dlVgEKK9WcRr/Z7di8jm7MTeou3oxm/vARAVglLxO
HqXtwOf6m8ku24uwQLmeY/103TKon/fckW2wDBkdb6vEYpJTlJm25S5fK4zreGIS
IXMJwzdHD0BYbsSplSzCgd/qVEysr316ZM0cT4wJcTTNLdXo71Gf8n/ct1eZxEmE
ZgcJGjsAHqCTjuGwEq9gdMiKdkrZ7ThMKfKBEQxNBlnWEU5qO8921WATrgrzB+xT
BvmmeJS/Jd0gFMdmNbAJz6R/6XLHU6JSQHvU46BEaDupuYh74RCfQMFGY5tnB5Cl
uORqV3EflID8neUhC8pvfGrj6cuI78FUlLedD/fmhQetg3fLO3un/3/7uXd3E0Sk
2VsRmA8xwcgVyowqKqvn8lCqx4vKsDsOX1VB3XgVJhnT3LXYMK8jlS4FLAdo29GG
7cenrnXwF8qyRawp84fJF5HgAZAAxfRljmFYseNMwEzmVdjRENccIp1mxI7JqGVg
njw5YLWIjxexeMmQRER1UBkuoZgQBOCaMJ83QDgIX+L/1lfLZ13BBt5tDs8vv+oy
5b4L4IAO5HGcl/yjN1UXbyy3RTAhyHMA4Bv15zlDBNaZyZiMU1uEwY/sn9z7fhIU
7E+GS4dEMGmMN5n1UffIHgT5s5+9uAvSH1ORBkZx3ieF/wZTnoz+sRgJ1yuCKmSk
LfDFDbmbIvmfg3rmErIMmsfoMfLicBF/r3gl3lZ1N+q97jUu3Pum1DvoctFqaZMK
NeBrtqICOcfArBAb1Bvvf1wl1mO/zcdlpG2UAlE79MY2GeOym8qsKE7JNEobMY2/
FK9Ler3gEjzr93quKLH33DXzX1sSzqt0CsZ+4A+Mu5DB+fIOMpM7iOL5lULK+uZO
NZH8PdWtYvwkZShcQK/wRoeMx9PWrvHdDbKj1p1H2NQEJZg3tnTx/RgNWZhCbG6C
F8e9JzJbudusl+haCsuctQuonW9D5IuZ5zVujD99hVOiUADMlc5yn7FOC3FYIb91
zw/Yeni7exa4ZS+pZ9ONMDcDeuD7T6cp0u9+vRRW0sSOiBO13QX+RwqbgB0hP90V
qpS7jVA/jmWk0m0lss04/4DAaE7UUoM12MvD4+ZCxLch1ZjGCRWRE8QPjXZzf03j
g5AIyszC6OmSWON+Df4q4r6EpSvOBrLgF3a80BJcZTjWAUW0rWzRhy4vZ+oKnztR
8chZSs+o1x//h5/HYE/px6dZ03/fNMXsp0XjzczE7BYRL5UZeJKZu4X+2kXOQUh0
Twt5+XjIBNeW4n9VXFktOhGl+53qJD9CXhGG0lSxbia4luHGSOG00IOK1qiT6cOP
VWFfJYF/88XG9dHtVq+RRW5v1GZzXeqslswOBeYrM2XWm4JgJKCd78rNeRder0ie
EL4c/cON+pP2tJvcmsTqE26eH50cBaUI/hv3KTR1fphL39or7NEsfEM/GOo8GQbB
gfqIn0li3T2Ro1QjHE7i5IApMgVZnbOZUNtQpx+4DwgqgLVmx2FcVoifGokWoJL2
hIw+IWIADswCrXOReDL4DtYGwwXerlN0DkbLy3zkGwo7r0zHu77QKJZvVY6GthBV
yGzV+J/IPr9GutpLUyKbIs9sKdTnYrt3iafcIMBggU2EUMstyNn8O9OyWyFOOmv/
popKMoUVd+zR2H0L4dS4poRoWjGyJ4VxuZ7Vr1FsecmOH1yD5Fr86caUo1AfdM/O
Rafo0D0aAOLGyuqWE9zVNW5HTNtrnRlPMv5ptf+EzmELTmnolphqYPBtw8YvUwWl
8lmQyZJU4qJArp7gdYEXrEY25hnTcDmt2iHJpGspvcoR8BwrJAlmZY/Wm0caBQhF
ktx7mmMXDtN3Sx5q8DmBBfChqjlQZUqPqVttAKhtvZxRL3Tvf5o9Cjc7erP+cNsf
nb7k0cUNNw9nkupXui8x41X4uaX3mkzcJyosFM/Bk9VY9A2h8vHlSDujs2xfaJvD
+FHbLHk5M3/dvjqCzY7SmMLh8hvytT1v5L+lsaQOBYWyacEPnCy+xUGd14pX4ZAE
ArpDJ/gW0sM+0p8Rc5rcQimrgDlMLkjL4yw562nzjXViwrLtgv3h523yfkDki7S4
k1QpdmyVQXn3ZxgV4ybDt9zk/ogEs24cPP1bUWdT+md7IwdFKn1xKmyS3As6J5X5
TGIL97CH1j4j5rqYNr8HFqJou9yvqPAX+qoyH7FrSYPp14tZAnnuygtzXLzuvys6
+ng5YYvzXovhQcgGH5BopYS2QJpcK1gruAyiAPP/ReCW+xAVNsLKyPfKweZXcpcH
UgZ5H3sKGy7GR6aWaPCEkiTvAlpaf8vtoGjKfze9UtFMMPtIIc0vXkJAqBXA7Se+
7leHDze1BFaoN5/fj/ZRzy6WRbPEE0Iq3UPR+BJ4BtuJbF2cOgeWNdjbd7ZXL4XF
HfUh97vwFqoqnLbk5+jriqct+elaoBeiasXsfA+lgPiY4bZ5PV6VXVABkvmXSOZA
Xqv4YK6L7ETB4tP/VQDC6+WMqWUb2KTXrgTv6nI/tjUgcPyfxp4EftXSJrWjrokG
OVTQANF8qewBhBDr17jpb8v9sJXEKIhhvif5NgV0RdLI0/Kj42dWEkouszgTehio
z5dmow1nTvATHGNEELrEFqx0bNYUPPTn4fkfy1G1ZyQsigcrVDam8XsvwXnTDsQE
xgSqk6y2gJsZFHv3UNcEh2eUbEHSc7T8Uc2CvpVWDOl0h6ib9x04CqVO6RtGmsIs
p8wHRIHV7J5z+9B+Bw8UBpaOW4CD1vBBcj6ozcLFmjyTJUQ07hmXXzS7lWWyx8FV
yNeXbJT60xFn46lf3c9u6NlR/agjjmpUOhpVUH3O8kPJDE2MgzmYrNdgwjzk9TEB
th1rIAhZkuTf3+k68kl4PSVA5blsfmDH8OngfU+IP5iMN8uXT6kq2hmb02jhw0uK
yz4HgM3YN/CFwBa6n2wHT1s824ErLhTnsi9KaRZWcKrZknAGVnn/bEUwJGBCfsFd
4N/5WA+UHsLZdPOW5ANtTELp94vpZGww8B1ZKx/2xH4ObSZ/lmq0uAYkSg85c/Ze
bKceyeoPFoxPrYfegWz3NsLvFUw95OngXq1g8CjdGN/gFt+HrMCa5FFamZ2/5DXj
NifmH40y1jJuO29EfiV/LXOKqbT5yGniQCoL2rKPVaZ8PWr+dVHT1wrN7vCwZCAx
KCy7k1PuO1To4vYtfv7BDczBPOGO4ZoDBDzS3UAhdeBXujAlS+2gQSp/olIUfeXi
+DZB5TZcqvrVocD4zUFXP0Kw2LMLw1VLAyAYAV3XcErjmiRRF0ZHiwMCp/b17Gm1
gb8qOM//O18cZqjdDKFJAicsSdm9lFDAcwv59w1sA3r+6TNjVClrehw158rnyTXb
z1UijUq9Jyh6uc26Wdpfq84sNumBsK13Qg5hjFMRBd2f5rRRaIfLmHRqU8Q2cD4N
ynhV5hcZLeEk6iPt9Kx7Jol1jMHhS0JuY9NXyzDHVnNZfOXEyaOlIgi2bMoGW/g/
c7yuMMP07vs2An8N8vss4j+l0s5Bn7+EQfnee3vZMaD/IK4LzFKz88TBDWuQG0TC
6ZB6DknyqIc2tnWVoCP4JkRThRwEoFbXk3a2JoVR7VpreqBZPBg4YOKyQ65Lwf76
CiZk70t9H5zg8KJ53Is5xc4ARd9euA/3EBhaWQp4mRx2Km2MPFeSNk7P8+ZWrh/a
v4wNN3T2STDzslSPhoEgZleHCB2UGTt+G1zfXvWy52reTQM8ob0G9kTuhiAua08J
m5R0sh/ygJ0H59zbj/WC6DyALtsD3Mnvn4h/HHfkvEs9rgUICSQA2gVKVCDdYYdr
miKee55ZOqiTGknCGu/bYKMCS3hnjfW29b3oWqsFFKism0MX0zPr/JuN03Oaue3z
/kHc2KSTptKEPDHpZxSd5G2fNxXeGsOnpVmz1K9HMriGlB6cwnc9/5qLv8/WcWlE
Ndx954+KizgqOrjZm58/+eFLZBgXYinew18VqWx7xaTBIwkgpbyh+yllJxyOpg6K
6v+YZl5vz9Hcy3cXtPTSPho0s07go3oMs65tVp30mYSROkn6Cq3UvQ13VNchh3Fi
Lf3wnxC9SBk0mG+Xoo8aOvAkcvpmbRqGdN1h6f5NOO8xLzgvDkv5wTjQ6kfW0cCL
ngJOpvA0Fjt9+KZk9rSe4fMk/d6Cvahbg/glmeBvheyX5mObcB2+26oZ9k2WtgqW
o7fUW0wwmKbb5P/Z78hFUyhAiBSxaMdfdYg72/WeZ4/+bc/USAvfJPzNHBMHMNIR
eOh9W9wDAhvD98T/UI+ReUpG9xvmgbiy+PV727XC+MQXlv6Zcnye79hILQt4xqTW
vIRB0kGaC3Ss0Di/BtUOyuGUXYeratz8hGw4Hg1n5mu1xcc/pS2mSVzRBwPrD0jX
nc6PLJt/BFhq+5nQPTgUpCbAyAPctIeGxaoCLEZk5M+OHekB4aN9xfEtw+H5sK8J
aevnqPuaoXrwpaRw9OtACHer5YGokSTt4IpuKO0byvGDjZw43VTc5jgLijqYOBUx
olrzLKhYLrENfmBaOviA8F1GJi11T7J3AkRVAZqvavDMHvMhJ9dC80N4VpqQ9rNt
WJPCCjnyaWMiJSWxBjKltyiFkkfU4vpB1imMOEcIGMnO2MaY49olYuw0RwM95t5R
CqJ35yA8TQHqKmJxTxx6feWH8mwu+yCUhqax0F8MvrmTVp70/1ISUUIIwp2+cZ8i
mk/1PI1i4S2DP/ZDMyVNnbZJt/JYoqV66fyw7sc7tvSKu+c59iFc9F7Dn7641Jdq
6o7rMGmSgEt0UlEPqZ0xMhlbaMvCEfRlMTKPhIeCfZmQAy4wxPCLj6+LN4dHXquP
P4A7rau/D+YqQ7i1kYJ6zrmQgiHek05929jM90DqhB2tSVMuuCUs+avUlcOE2Mny
X9zg9/Lu1ZkMOesmjO4Zo0ERVwia7THKU3QQsCcrK9wgEuQRt4KF8IyOjta6JmSK
CXMGhNP+XdUWaK6BcUHshJBti9QoTqs8QdnjxQc0PactaleNbPwBzOF+kvHlnc32
RAdlZ7OH1jeOrsHlzBn9PuHCiXaqkNIOnaX317GxZoAxIDCrcf9cokpF6aZK3eco
8/Vke7B6b0Mh+oKpVcKZG9DObqEU88HXZ8zrAoCy92OIR0jSL3J4XyEdNa9Lztav
4vKD9F8aVmXPhZTVFGrmKMx5X0Ewegb8vVbRJuRHTzOxCIGUdHOOdEDgz2n2h0/d
J5NJSUq8F1v7Fb72JZydoVCvTDa0VC87WTSLkYaRP8pMu0hPqQjpXQMNKhMDb+9o
xXPCi3w6B3/4M+VI4FQMUBN4k6W2trkRCZYGbxrckVVaG5sc/KnZ28J7lUdo/7Mq
4/6HorHoxX1X62NTSFHb3jEOyZB621MGuqXD/Wor7+0xFRZBNoBHIzXTDDbXpyyv
OAfY/4UvpnefPh+zCIfrsnhD2YuVqH8zWbBnd82wKzNOpa+MhpgKkCM93LzqsOWb
LigFpSLy5Il/AVhH8JzGdx4IqR9v/ioz3Mk1OXr+VDj9ylNPhKiAXpahfr3dMndE
AN+Fb80tg6JTsdlGckeXPou2vYXTzNQP/Z22GlyAI+encSPrDKdexMX2Wdxe5kar
4eJhXk6TDUQN9FqnzGp6VzoysisXcWPpzNl+lmugTCrLVXa/duicRVVNcSzAeNuz
6XfAdsVyX1ueKJBS59RIu36Q8RPhoYS7EhkFRkBD5NTbgK9rHxMAKxy5n6BNGQdA
41aR0vFywDFRyC01mI+ZrpwcNHxuHNN4bHtsbPkH64aiq4DwX1xc94yEbnSKIL3E
qBMXRPOqzJBs1IpxMPX5/oHM/3aDbE95VpBkxFlr93ArQUK+YXzNg9WMn3A35cxK
nrrXNNkXEmPUw11p6m8YlFyv65I1pakRFvcPmy47pl6fqjX5ONmUZjtd5U8U70RW
kau2SHAGp20R4uZ6B4EBF3tXxr2vDoto966uh00D8sjlCXoNAfCZdCnbck2TeAgE
HyLIQ1cPz3cn64z/rrA7WeaXohMlDc1SQ9tlVI7iH8MrOdReDHbQSFDmZkbRNEhV
BoIYTYiDCeGrnijtb/3fIDBjuarKRvxYbI5S6lQoD6JNbQHKrK94muCu6rHQ/9Ne
gDUhsFo5Rz0P7xCpnosGr+GFjOGperqAr4vN/lnQnoPZ8AYATsrB+S1UMe1az0PY
TVm0EXGl3M0osDDBStGa6VSZ0IvwwD1XP7MeNC+YONrEMK0G5IP5hcoI0t9HfQwH
15Po+cx8il7ZLJDgPwZxqDt0Ug0X57kcmfNPdxIHMm1DR29RcALDKoJx6C8EisB6
B9P9fO8adRk9LWflibq3V4EeHckj4HPJWIMgF+2qu05/LBSqTkTmAxePEyml0Zjk
SVLoxcOpbVvVdyiFhZnxpTjAyoWhPd6NVLgtwKuDHMatCkbTV9JLSrZj+kfdDJMV
mviV9nlvO+Uaue4iKpciquJ9yfvV25P/pcGXdPbnK/Z4GytqRsNRpdhKJHeFfNnD
GefJlY8qopp8gXv+oQZR14+T7aDW8Idn7UIOtWd9d024SJjmjn4moa9beKE6JF1W
BjjNOZmsb5L0DC75EEdS0o9FENxlU8JlfD5l8C5nML/fKDDE39bHJ89Bdl0FtDzl
K0RlA6LV53EWaxnZhIxyvscWdjv1UWsa1p2I3gFuQTLQyAtxD/Mvf5upcc5oCL7q
e+zUpJ9SnD47hL1kAc7otiKYgMBRFwCs7iIuvrqTiJ+6n6bTKpVTsLol9lX8wzIY
1BtoeNv+v2WKAKInSZLxiVCu1mN0rorImZQfaOSAvDG/bdccfRobk7l/aelLnZUw
YF0hzGtE3nl0O4iVJTp/gELwTqr6Ecl3vcepzBER0MXCDk4AZC20w2NEndpFCUNf
q+EkLQ9iY90MItieaM7aWYV7QQ++Sq5SG98pe8mYXHCmWnqsEhwo4RKUQPkatSqp
bcSJw4TFgpk2iKfhGINjnOZXa3DzSSKUortBO2czLZtlIJgHLzxHq3YmTArowOm/
SRVCR9UW7Fv5NEV/yTAWx6gS6pL/rBntbME036EacKXgnJ8WeuS2l8qfQac6Dvci
ljNQR8b3JITRW/VosmKA9hD5oNFuM6A3QoUKcHvt2MHjsYizyUmxZ8R5Sk2gSjhX
datpyDHX3Oqyr3Vpo9iHWMdkkhzwFUlbHilcp2Bu/654XmFvuO7OCPR+0LSvE2IR
NRO1QLvh51WjbhBqunMSRyLnPH3VvwAxvRB4DMMfcmWKJMGXUWhKcfi8VF94j9k6
SyMUsBR8W/r2SrfNcfWizCnTyFcWfqMODN2RRE5Utzupq/+k0s2piSZt+35vkLQA
eBWKfXmUFHdYchHwupyDTKrRtQWbQ7rma/hJSu3SxXG9ejVA5U4NqHuJvjvjVPlS
AIHgjPjk6nhsWw7I2dUugVMeRGNy2tGoyx84FpYRpLBsAh5UI7Nq+PO7AOlQjaE9
RJA308kt8fZjNNx6mUKXC4/1ZCAmQYpshitW90B74pafvWqj59CzJcqN4zO47BQP
45DZK/UYXPGX7zXjjYtqgwccTgKiRx/qklSyrZX7b6byDE6i9wJdvMAHcUD60cQh
BWCXZjzHAXWismhXQjnEigN2pvCy+7sRIE95Pe586azGz8NCesi9myhXqdkThpvB
Dqj+EFdBLfbyoVrkD68ysfh9evjOjnfmiSLTiYIi/XE9k0W1zpVuLsrZmLG84Wb2
lPfkBMx1SiVWA6P0iER9gFjKXQGmSUi/QDPs8G4rBFF+QHhOy3TTFIPbeWdvqwxt
aLIqB4ezwOtTNQywI4+l6nyiOVwPkJA6KhvXilUJ+6zlU3LIhntZ8x6gfs7EVwL3
g26QbrBUc9wub18e/PAi9N3Mw6vEpi78LUbxCTytVFgrgWYzixfmePag8NKRzQmo
qh/I8cLX+DifqbSpt/6WQhrh0zYo7ZHGnH5XR8Uzr5wkfX/q0SdLESe0fbzF09Z1
F2gBDp0ogYyelbQ0lCrp62800cumdCWMfRh1Lr3ba2iaDUpZ58VkEiGZC8ZECtqm
4KUBgxO6uV9YfulP9Sj4AP58VjYbFswPUAUQz1SxB2NiQr/V/8PmS3AgjmB9qTz6
Uqjp3rHnM6HedK5+D5jrqWI1+a2dOXec71438NM3qI7qz8iv+NnY7+BVyQhWPVIs
JjcksBX+Pxuknpqelmtl/n8KmxvqtsIe+bvWsDBdJebGk9Fn3E8nbsnTtIa3+Jwe
Ukoquc4JkaOpghaZUIea62lweLe/sdu/fnuOMUIE8jLY3KBRvDZtcxaJKmnXm0Ut
wjuD+qyJoAqEdVQmofxzsMAUIcQQ5EMAf7kkOLas1NsGFT3sXOEQSSg46azjb2bq
trQpNUHVSmlVEUzRjkHmjCs4dVsFMz9VEeXXi3TCGtOOg4MvQr9C9PWJ0blmdL1b
QpOvGQDxfPpLD55LL4PshZzoP94tgxB/m6H+0Q8TV/ISb1g8i8pAs5SVIO2Qr24r
p+ftPKEb9x/tqS0xiq4DRGw4z6Up+aWcGhDa3G4BZ5lUa1sI1K4bsXn9I2O6qz6c
jQXtibQgPA0/3I/fGCuzm+z0QKroO3TiQFSdGgtMuwcMaahHjn+pw8pcim9Ft96w
6Gq8rBnE/Qyrn5ViDwMKwXD0Vw52ul/nGWu9y4P7fWER6xhbDlySy2qw0J/FhrJW
c9Nj+zMH7jKuO/jZWam/HtqnB/LPGSfCzyw50XnzW3jSxE43KB66QwJYlCYSnvON
lStyhVBmtza2JE73Bg+TjfqWKWwOJC1pBxB0vQmru4YWWgcsMCbeeja47LOrkQ57
m2cO3fVBS+olcs+woT9Gu4hdRvcs6VM55Zbhod7l7oDgQLXfAedre6MbvwW8iwWY
1NClC0NvSNgeXO5kueaqmX1MVJBp1Dhr78Fd+G3MdoLYuoM2aJgaSbna/FzOMURT
8wFxqjBWfZkEBAmnB8pLWPQAR+q2VGuwVNAx37aIwoiBS2X7nzatnsU4ivvpLaa6
rs0UwGMq6sqjQ6Wfmy26qHap39wWmBrEhTub+ftleVdBnHnj0YQW74aIg+l8qnkr
Ga8OqLQ7V7xrKhxyw0f4aVNfnXzJbhAHj4qKXg6EMWmxIzmnDXp+nXvPUZjSJtO3
hTdhyBmrAskPqGausf025a1+YuclojOBtiPZkT3fDg5x6zLJZS2CntZgGz2ZLK7O
/LLju/3zMysCl9Rz95HrQ0ZswSujpgl8pSp5DmG/aaDCx+GSPWCA05h70fFoNmif
OnOVZMNNVZC9nl6KmjBQH80O0rm+cpGDePCbshTZZnFOS/wbjV0hf7w8+Ab0TtAv
kwd6CjRsNQne5k+X1kT4qmgqvPMPfK5gF2ReHBUtaItyqg9bdK6+dygJ+SkRnaCP
ZJ/Kr9/CpLUrqBcUKsxWeXtCzLBlKDLt/toSj3tn6Vq6mTwYv82XkZDa7pjRo571
wWH1m1EjMbguY6Ojtk5Ntbtuckr/m+M55bDrQta7PyF2RIB1SG+hXMiaPa0ySTpo
a0F3S84s/c3YU6cYXCzSACetD6MdO84ue/zkHhYwSarp36Fgqb4OCW4jhAfVdfuc
vZCBZN0nw1MV0U9LzZDZCSHdXbs0pmwy3H6+BwdJ/EnJKIAPnK4UtTV8tf7Dzay0
oVHJFJwl7M7vPbUT9XuYz9PSm7VjcfsDAlzG70Qjdj9uRb572Wb60DQeB5uG/Tlb
ln5ak2z2jj5neEIJyyNnNKh6s3jmRyntdO8uxAGoLM9waZ/12rn/4RodtSAEPGhk
AM9vGjGtXQvE5rXrNLdh5sxkC7dT0CbtqUAFmn3E2T9u9YmHUffiTCcV5HM61/P8
KFrQIo2w+IsyPIBJ3KPgejfdjQ9WEhVtl7fly7PIdR1xmoPqNj1muGuHd/iKMimg
OoCp0DqmaTT6yS+qq60E+jRmEocRbLj0SD/w1+DFXz/7wnXQnUN8NwvMwqypjQwg
oVMDEyhBn4z1jBXu0lRNvv0pIgbrQIeoIjwIeXEPtK1jKsoQENxorCAweSZUUyi/
mLvgPUPgomDJQn+L1NaXwGdrPnKsKQxVXS6rGOVAzny6KFGrODC8NGcggMu5qg0X
7bYRQnScCxbRuHlkdjLwHUS0zY3ihtXzlav/M7DXifWcWSYR3BnINrz0BQqg3JJ8
yvHs5BPk6a8i6ndZjUrTXmOkuKd1U4HsP+sEpT/Oj20YpwPRpP6Zm9feN8rQBn1I
flcdR5j+QnKrbNSFDQ792ExD6tqCmMA5p/lbLaAVgza0QyVSGa3IO5OqM6tCoSKO
8rfg3b/T2haeG6BHyXQrwQrlA/ZN4lPYa/NpJW0GqHTtA6+/E3bjwus9FpBWCeoi
hSIXBISG38mTrlIJ5wrfZMGqDFQbldT2RmLe46tQz417SJSVnKjyXbKqN7IpOgp5
JrsTtUKpDOdnqZq9Q2yBzXmhuYdveOHQW0DVyjaL4wDPYvLs7OnQHD4Mef1T/x2V
Ajt4VLs4t7+8A8ZOFcuYn5/j1htQMsZbm8tHgWSkjD+ZpBAW560DftvnJLY8sdT0
/DYSva5e7tY+OglzKKwSbjJFkdJpVN+VBFwsnAq6TkQflFeX/BlKmWNnn0+9i51P
71sYsLOhEMeEIZv0D5Ayi333/FNH7o+QlCDWboK19FcWX0RUW5W2LKtSWLI5wD5R
iRXmax4V1A8MWy0BrfTTD479XukUJT05O3aD3hP0RYCFofsc+5MsQabn5ImW+XaL
6vX8uSIReFdsnsGivsDIztdGaty5zEX/lspZOQvK0Ooq7Z2XkrM83UexxqeX1z+r
RQ6DYBa9B/+aUI+6S/04vCY9huH873oLEnOBLcX+HR4aTGxEQPk/ZS5w/s2Jghm1
uTLFkM3a/XZu6kMdk/tbXAzKyljpC/fv7pMahfKxRs3OGbSbthCSnbje7eMEXt/4
2wIgMW7jn8gbC+NDAa0UKpiuQ2XOxsS9kFPbS43UfZMpjkrqKuUyKYwIsWLr3Zub
rphX1lrP0bGMmsv76GCeqpHXAVpPFwVqU20TkX9n1/PeHhzvYU9Moh2aiMjaZafc
lamCJPIt7g3KFPsMVDIks4ENFdeBQasiKgL0tgCTOHmyjmpDG/6kO2Dj8pAIb9mM
Bxzsb22YDwXF6w+GVLElfojqTk9K0koleESSBYgPoxr4dKAcNF9SCybKFV0ch05n
yVcyAf30w/1MUX2Oe1mZu2OImzUeXVBK6kUJtq/St4lkTFkSWKaj9ndbD2cXQ7Vq
3SnLQIaZdWCZt4M9CkpeTTENpL4K2ktn85gWzVd/aszThcDuxjW+9VP5WQA3GAL7
JkcHO4yn0Lq4WGTmm19MZSwtQ214U1jyI2e9UO5LeEU0V7jt9zYEuWednFud/zcf
Dy8eaBfqf7OOJYOwW2zgSuoJi5FQeTADapA9/8laS+SgfLKhTCgxkZFPJUGYV8Cf
auqp6BH29uu8oQwed1JX4hQGOKifWI/hIQmApKoe07cacSrOSur6OGToCU+TDtfg
aqksQo17KLiUKbe4y9xJmRiFMv3zSOA1333RhrCjW12AubWcoqxgLvraHrPfR7yx
IjKbx+IOgAshkUlTiqgG1wOvpZPbFiJjlsB5XbqGCMwpj0SEwH1SLv1H2du1gj6V
bmeT6SOYqPFdeGasyRdd43HMvsbtHp6dSOve/wR/Kk4Lqc3Y5C/Lb5rZcnZmnPp9
/aOpzrvB0GWOxssuGec7wpPQYEMsf12kUrPc3hexrgNXKD0Bym5LCO+vOhJXZaDC
sZh5BwPQbtnTDRzSHL5MZhsnGcXelinX/YU857QD2XbnTloS6OG6wsS1R2AA3MaV
tmHAqVZxI1H21zMX/vmuVR5ZPOJw9qiJJfgSU+nOATmkRfcJKcNIZYAkJDrW8BPx
ca6AbVDwesbV3Nqux2rm6+QNpzujCBPOFiKO3ESF0242K7To754Wiqms7hSxAUrZ
BGxbxairHBMgWJNfHks2tqCVPsnxiL4QhcxXAQn51s7QpPTjFjXf745AEU1Z6ujb
E4TDEneLMmc8OgdhFowTME20l5VVshb1g0TPS/qMcH75xNg1RyOkJmKki6dcOAB/
ikZy1gSsn8w6PBLF/4iFYAcVEFGqlVhwX+OEWvlrQtr4WVtbcoU3P6nu2O5eXRzj
UYWUR7zIxHIW0VgKie0cY2GMI7+enGovJG7zO4xJv0ViqS/5Rt7CmAXQ3IkgiK13
dPos275DhWg94pEnuTcigGhd7qp7coLQjMM4bleYp5s0FQHQRy5rd4W8t1qCO+hk
ADszcSCl2ggWhW984SHCNcTbLg3pn36SQAjEsJUH/WL6OYa7GpA/nl/tMA5bPwy+
4iGB6c8temhcq40MTRASHiD0qdrblgwjPBakvfDQVCEhjOv0/lv9nXI8E9sJ5GSJ
xakC1J2qE+gsAxulzeFki9x8e1mak23zpKadrIOMlyUoZEKfF+IjD98KrNNzQZiP
b1Y0F3FRfslb/FkwRNnwoHXahRDcxn2E0sOc5ZM1JUs3EwPbfh/wFtPGp3tGs4pH
iHO+Tr4LECk6hqjP/e399gjt8jhU5ayCOsYMlVCaKaOtzxlH6JUOHbFaf74jqzYG
5L23nTBNRS6Yt6kDx6w5jR+IS+k25ihiM6fxnsnoLgCgiB+Mw7fyGJ7IjcQH5peS
DzD2TZnaT/kuKJWhgcFTBvrB2QwqzVMWa/FIAxfPG4U1taE1Wa7tJd6EE+EqStWz
kISk31+FdQ8V1GJM6w9ddukGzXv4VHgiUdgTZhExnX2ntJxMIzzeEqcRxHd4lcFY
jzJQ1XsWHlR5CORgBr/ssQtiGSo+sTuQbvUsr5+zwDEdaI8lkTs9NamEtyTnkax4
uk81eC1XEzTznaJ2Xds1zBaoCSfv05fcGgwRYJi5mf5eqyYYIrJqgDT7MUyhzagz
n4YvAA+U1Zss9NZEol550lZQIWEwN9F3U2E1TEnT0mcw45JKEU0POr3T7tYvQwgv
Qh6sbjnbNfg3fwlulWwVXL5tw4/Q62Uhuu4YLzLRYG577GWh+zofmA9ZUFTlNUYo
zijFtY/2Ulj3/44B2/h0CoInRTsQV9VHV9V1FiCtX1PPWhj3/EaseF1/SWezIBpM
nC0BMFkC9fTUAMszTxRhgSN49AXY54XkgCNPsuRNxGcyfQwM6Hsy5skQJVJ8+aBp
urgZboiJJ4Sm8qQ3HugU5jbe2IZf972HwZ8UQSv7VdXMK83prHFFkwF5me5VLOy4
VpD2/0rTPW/BbiycO0Y9D/wlV0/eePzy1rfAx9k0jajidgoMiS3YUAuRSX98rf08
e/kjTUmzlxLiPRjbbGw1EIQ+p398U4NzLRE9WGKPFyouLEG8UrXBhG1YAQ/SAW7O
EV3uA98SdKDLhvh1Ih1AP+9Y623Bh6Ul73TrfmGm+bvNVJCoLlLZc56ovsM55AZm
IdaTm13wt8626G7S7bCZf4DC+9ZsLRikZjjkvYxYpqWXQ1sB31qHF3+WEDatEGhN
4FwjOWkvS7rCm3iZjwkXrgoQY2+xcCCDtx8usSpQBO4ljlak95ReovTxsUYI4fQh
k3UZDSC0DG3tSGeFIs03ayi01ebeU07hNjbZu51xrW6xCQUEz0qP8X7hXnqpjC52
jr5n55Gs5+cyXI7Tf+ECfhe+ObRiTFBwxHc9aDaQ9kHd8kofuVplFJjdshwJmCVC
6Wf4miH0sGeErMWiiSNmZR69eSmF8r0tBZnqdYbOO4QEuoD39CWA2pT3kbzrUAxe
ULnZA+4L9lGuoXfPFfE9s4lgS+7Xm5wzBJYW42GCvb4aI3z4+gFo9V8x0W6rAN0g
h0JZoDqy8AA+gsAuWfqOpJdbtgfHxiPIGWLvg4LjRoWOpksKyLicY5EfTl2EEQFD
Cr5RBH6sksfPy7U8MBuS8djFJo+kRHTJwStZy5W5MHBwuZqaTwpovWRdkgcBEZuN
ToVeRkCvBXk+m4/ztvZTBPPoCDYnHUPAGtd8St1OtN9crTESMGuZztsa4SLlD3s1
KV2z5smUSoo3uHF7PzcKX8SKU9wcNEHHkTtSPSH9EKg2Mmu0o9/7dkGDLMWGjBOr
OeHPzHM0s/Wc6SXnl/0f8W2GWplDfUkv6MR151t7ZXBFa6zQjR3lz3yjdyILShOP
0yG50jEGZi+4FAyOTG4CGKKGbI9y5ArSGJVWUveOUK9y/q3fd+ahRBTZauQEKSe5
DUbDmBBuOL/VMoew7m7HRCrShLIlqffo/fznWfoOEEzsFGQx7osqkK7/0ARmkxS5
Znj0g2vD6uwajL9OM9BPryJ/4lQfucNMQj8p8LA/YLZfgnHriJ1M1jIJ7R9nJLu9
IMmtmev5f1B1Sm3LFPfMp3dMF5zfCjEgNd0fGNl16UfL7huTNx+A92AJfLLWHmiD
2eASeypYpksgc293a+eIqrGx6k7kODIIiRGo9KefocpyZlWbZC+rvD9cZyMrXlTs
DUXnRfH2qXuBq0quch/2adtzoRgR1owIQYUXeUXFtJRmXEsNso+s+ShjlUW/DqDz
YSoh+grQ7XsTjBJh5WkYWs0DCnJjKqlaFzF5RWmV1NM7lkcVJWwALudSPZ59ObNY
pDB9qyOYoxHk9gg2GDmUTOocqy0Apc5GxWQYwBHxiSTwDGxtt9DBsDpjOqpe/9+f
0H9T0/W4ZDBzwc5DIerl0J5pFesVBw6/L7gIPgY4DLGk5FzJ61lxCsKsfAzzQaMu
5PSt7BHZdPPd4UECYoXWNk0y8mNYMibbD4lmOK2tzqLtrucGgcTeYh4MA+y7KI8G
QcqTtjuvMnS+b+J+xEjc4D2UNqikWYXdG3B3GTuF3uGGmtc4VgbWHv0aPAFi39Dv
KCp/sgbIq9QZX5ii4Eoahgf8Hd9HhaEA6vyWw6ENE+ymzK4AsuZPdTUZlMHD1Hr5
t3CVYprf1VuezCDNrR3ZoyIZ86NOkkneh6OYZM39VV+miGMpESp9pZ8oQzUYGEy7
yA1H3EZ785R1SJsae7z+6DUE1lkbWY9+GB2R2M3OKv/o/UyeOBmibtQnVk7S8fzn
+GmvFtU4dO3ANeJ+UxKdS1lQ3R4aO3WL/e3hAhAKosjD8hRWS7/Ar7OGGi5Xo0Uo
irPJYXJ64O4k03oeKOK484sAAgjA/eCAdx9k0og5zQvNr420cM50VWsU7QGB8w+7
mzBho9KZ+jENU5owgzeFh9eUmHCFSlWLlLIpV5Y9boNIiottXd5/s4BaQjBlT3x/
gUNJbp9GdFDVemHm3u5JydYJHc7KADE2jqUnIyPbO24nBtYOL0BHCEMF6vmmLTmQ
xStsl2Swjg3g6jsCt+FTR6gQQ1a7QHx14P3thKS1yIlkOmgHe8U3XjtKlaLrolC4
QUid6UAQdTxfa0YOupsam0oQTcKBlt3D2LBKYlLrS1RbQkY24QqqVPNQGC492ILH
7TzIQToVlnDI79CPUXVfrodTsLhlOuEhdoa+ijV5uKkL57g5PZVE0NNBwjilyvkJ
59SokuyTAg3NtnBe5ys0F8oSnIs60gvby8h1SDnj4ftRC6LFwCM71agbFZ2u9sXn
4twaloxHf5Cl+gghS/zg6zoZRaXLoxK0ljvBLcvTh7iA3PdxYAsNKr7N12VL0Ib2
18RWI+9V3C4Pp41hFCz1QEjRZiVR+JIIZS1EYS8SgUTbyB7wEb+0ei0+3317VRAq
PVwUZUPhptMxiVv0qofgipdqkiVOugdXBp1Do/0zLDg0aOCLuc4XA7vYecJnKuuw
BzExHPj52V7btFrXRE8X0uObbN14o6Tx4q8sqXpdAMIH3a865E31RvQXoVJqtj48
9IlTfwDgB1fkyB+v47pFof8RhCFHfxnU54RrMuU/oAA0UybH7B42XSQ/8SeJ0EFW
wYqGH97GW3blDeZeim1AD4zYdHOJiqOR2UDFvvmVqJZKWX17n1261GZ5UagkpzuJ
KE98nWM0pFkXA7s9bL5JiZQXxSCP+mgmUWlJmXryNbEXG50sGph/+e1XYAqJPPZd
6btNi4xfcBEH7GKJkjmptwOKaKsAxdzjoWQCQ/ijBMNOkzJoQbcIyqO2a1mhXYtm
Jj2P3T5l2uwUUUAYCeCegdJI58Z1gTXlybVNFexQUycEPIqvmL5GyQEK8yMdwBv4
wNgxvdZyrpNx6VMmiXk3Pr1rZIRliDuBe7OkoqC2Fl27sPWT2DhGMUgjioaZA5dA
NJ4pkp/6h0umkc+CZaKqjLibByXwlu9Rz2NYkjtmFncXwZXWuOPXw6xSA4TRjnGr
tss1CMXSfw1mb3xjtv0S6r01nuEkNgKRGuEWCmoSGTGmL8eBwE7MnsjYOi02qE97
YRcjGuCw5b7Qx0cyJ7cYMdIas5uD6x+xrdPEfFBmvBkk7Hp9FC09EqAy309KEbeH
nToi/WDV0ijqM5yDHJRXpe0PQ8YfY+8+yGM8BQisqis5CN4PFMyS2nO/V4mQpWN+
WlTjfNNa6QJUFRCRkWDGsOFLIfVuYAorRFjiFRlz9LZH53AyHQc2DHYfkuzx2qMx
Sumrsswp8ePTusMM75VI3OWKPIgx9VskJuG7s6oZKcgvd88AY04E8erWppucP8LY
K15egZf0+CBEKrS+170An43XehwqDICmZb2s+GkYEyYy9Dv8ooDtf44gf0sK87Zm
cusijTjFOhEHSiADtyyBpOKySC7pGgVQRjAJB69MpsTPvkNwZv84yB8r754x7T/2
8trYTZyLhX/sOWy0Eq335KJs3EyKReq9fxoSxfNKrOT7FKbnoVcvakdghBuwBkjN
6b0dRVNS0ucLLD68SrEkP1HgXa35wVidWpOXmvLdu+FPCJStFC4iBxZpQ8rur6pH
hJ5wmzKSzUrBstHHaqzDSFrAvIN0wjAFV+SUEdYuvgl+4JgvBfngahW9xkJh0Awr
1ZxqQm1y+mQ/1O58OlQb4EN8rjWAfocAV4HAmeW2JdUUm3N0bqveDpFQD6W5Hz+i
f2NEeOJP8h2HYbQXStRD9lfCB+vnbvyGBXv0mHk4mHAP3D927RC5WP+eki9VBsKD
MWTKod64aQ4ZaO7tXBcxPpl+jncYB8Li48pQNbq/Ia5r3UZXXgsMhSQER3n5+maL
UajbjaJMwTaLdr7oYHBDez4yLrjTcoWoLggAc9sDQemVCXhjyuk8StYfD+fkFiOa
L+Ecgv4HONQQUK74AM+c9HGJl/j/U89nBVwwI/bsotXbt1WOsv6qRI5zcuhBKjyv
nDP6PPl8eH6SMH2SKFxfkummhu5lx0wk86JLAqKRrmoWjBOZdAAftEgR6aOWhKcc
mXdC5FdNVvnpN/OyGXSNG2STBHDWVCCNOYUxitvYgH2150gb2k3jS+2xX+0FQm9L
LvEY6iUbP38/kzPxXxZzcY5ScwI70lH/4OXvUGEVnNXA21URNcoTfxT9TrHZtNzg
OflkiCHckjqXiOTsvW8clrlEkeB34x3mVOdpoKFJNG6XSsearw+HbPm4bUp//cc1
tPy7V3vl0/9XGW64DDuRSF8iwVLHzYXmMCt5OcsfbX4egiHeTcIwc3pDvlp/yebE
vEUjllNRjT1dV4Mz1SEuwVg1MlukLAU5Bi7reE1qmhjDwB8Ht+mcATTU7ORhi1i7
iOw2MOE9Rr070yzu3MUEGpi5RKHRBBMgDVhLS4cAL96WqoHaPU2FRhSzAJob6vVi
/q1E4xaWZIjYRIHV4Q3DWaOK0K7om7UtHEeyAwqlMA+/CaN+Csg+X/CkdTrNW2tq
gdi4II9h+x3bdwwiGnDx5nuWBKcmGq3EjCJ7Irmyx0DNEB4u/CFD8mMiFBjTVDKf
7srqiEx3b+tT8lRO0t/slHQ9Bxi2yIALnoELthNOQOivIElJLCJLjBEPGE9VBE4A
iNSTx35/4Vit3K/NSlBAuKKMwMWPJ56hlC2r56rJTM4vcv10NZGR93z1UXoJoz/9
aBitoO9UhHc16bbMxC3EDuGspFOEDI7QUZeSf0qN4oyeqtdk3qINjS/mwFLMy5LU
hRYUuY0IVq9Z7C6NlVwaWRsxpE/IhCu+1jESkVbNDWyG3uAjUJMQkKLZS+sZ7Y+R
k4p7bvIZp4YsMZB0HKuZuJxkLP8nTtH2aLH/6MnSm4DKruesI8iyDzisz2XfuNbN
zrnyaHjKd1GRNebqaenr1ZFtBSTzTS29wEb7YZOy5rGe48J7YiWkvZ+o+wBMGGuF
cLpYUKY1HRK8oq5a7I4GQ85rJwtaqQqJorQ3iB0trebrTixidb2WeC7K0VO4S3Xi
CuRzY2l/Uk4LtfHqVTULSXd/P6GMMxA6L7rdmikamfFGuj7zaXP+qEUNIdO0Ou14
vUUrSrlN3xR3pw7WM46LQXtnKzyovFKM8THFYoF3e6DDiBWiUED69J+SduoVZS12
GiLnTzIletCbvwmTDXOx+jo8F8itOGORblZrnvxZXb/dFFBCbki36M3F3Q9F+nkh
QuZ/p3HgwnxRy6/K4xibBqyNec2H7aXQr051C4ck9u/PxfolKIqZgZQHFyfHt/m8
cJEIKTTLi9eqB+3evFYKiaOW5hkHtVhfK8MvXYuiGMW+G5PuzEN7WfebyxtrDl7Q
cftUsIzT+EvEeOnjxZLFiuAL7N7wuagtLBDT/ZyNBtZR1mtq7nj8e0uZ1S7WZEGj
DSrTv2Xl8UQNvzntUaM0ldqLm+ZRqteKFLix4jqi2EywKdinqaCBynJ3hYMlGS4r
o1lbhVeFD/QtmTKwJJvTPq/BR5lkHSO9EzAGOBp+1wDmCU6wQMUCQxCUCDlxe8Jg
3m0Yh4rf5zFXvSB5wdZ0ZxJPCaGE002nYgzZOxY1Ah2ZCqybqgZdVGkYgw+/WC1Z
GbWbuYOzezzbrB4ZEXbKg3/aYMH2YfODfwRJHtdageRhdvcobPtZph9vEhIFHubU
/21sT1ShBVBPgMoGRTZ5yRaCkl4m5+Kps8CeBHRlS1DkCKW7OqoAlGM1qol/inqI
fE86419SP0UnUoOx/KAgDr5V3SmzydjPcd5Sx/QuMK+9QK541sX1bq9FkbchhURp
JFYbI53KxiPXZLgksPAIjX+JcRVu/C5/OBKO2uqP7WtaBYtNMzAl840G7RfT8PdX
HMyoR30FV6HwMcGvxGfkwgIBQrhFRQoucQKZze4Pkl7H/mygvzwYD32q0/s7H/II
ghLmXvOWJC69cex45o3gNFoYuyLMCBoWujtssXA6kQSrSrDHTFXhxR33T5gYPCpP
mZSCpv2pAkR3OkxHg/nXUldfjmwQMPOGyF5hwfwUvSKyBYEJfjZW9kmTVjri3osq
zHu7Id5ujgDehEzGy+5yLor4IiyX4QUxRweES/RLKuGTJIGhK6jImjcu9O2GeEcC
HI0bKM46vb26J4j+pGz2NZRm4IntPbpQHks+gd4Pw75H4yfPD/tUrVWvwRqiuDtT
zwBxzRDLDk3Tp3qHxhP78ofqEJh9nufBjjU5I2x7BsKDt160j/vqcJYC/R82OQ+9
DjKndo3q15X7ZXKnne0ZqabzQMHlB6yX0JYQFdqJnYpSnGSfWxuQppiK3aDLyydw
ZM19MbQf1iPkGfExEnr/shnYINh/4sJo2ATz6t/pD6/tLtWkWutHBdFuF9vwDewv
5+Ja9kvOggMMGU869lP8l25iUGTE8I6h/VE6GMlIuynmOWS6+q7OFreGRN46zZ5V
VI+O+p8ATrlJTT0b2LkL/3k0YBkV855bkADJ/ef9NZ2yNm+hoJssIGHvGxv2YXW1
Fc7Jcy4ZhGMBQexfh0q8RSXIcQBbJQL64Z5YAjrpkZX+Tm5iCEgOPaQYX1Jndska
kjMQp+gQvMzBSn6CyScXivZiCy8SflogTNxPUI/nJ5wl1OrYAbNFfcwlUX/wkSA2
Kf/mvFG1uXP95ZDFKbEjlYxiOcKEQYKyc7WfKUCcTu3243eZBdogGkB5OnVqAlqd
lJDnb7+qN+QTDyoKw/x97dJ4/pIhRUe1scyh4Hv/jUHAWvER6XMwoileFQ9mAaYO
H83wlZENh2TH5PAK78/f39K+/b4xQbV288ZYybMf0TtgEvSc8jQOsMrLVW1ZJJRw
oKmbrxKFewKMtMJM1cJGu4zT7dkQvtdPWgLKJXhN/0HV0uP1XSbEeYCsubBJ9kcd
q13leCJ7+AEARXhjAGuCAY9bY1J5ohbPDvvQiHy/h3GRKuez8IJ3oHB1/IHouOge
Fr1Ot/Bnck/LJ9IIYf/aNXw/zdkzRZ8OgbjRdHRM/TPd7ByYrpf8AjNOE/RbGahF
+W4I25tUiAwZwJwckX7+HH0qQStuPX9Y0C6JQDsA3rAjhYXWeRowME9v9rS6uGhM
vUJEQ0ewP1JKCZSdZOL2V8hjr0ak2mFkMwe3sS9HlrDhykhegA9jkzGc2t5zYrN8
0Tx0f7hwEj+3eV7UOAQ7Mp+JHFpk+PWhfan7gPpFd1Xb517R39B8LsZE3eCMs1XB
aLIBmL7elsILO0P/M9w9K/9/YDBWV5xjlkrckojNsHqfbuSwIYOYAvONBpxL9/ok
jeOQOqSs9CguY3cH/tEQAjw7cdKYz0GvCmPMa6RsdgzGsM+bn4gQ9iJlGvT8f64k
giVLq12LyVaApcLZEW0hs4N/+EGHk5xBcyHpkSd70gTjoBXJnedwVOYnrD73AqLJ
6HIHOLVc+1YHZWEH98RcWXM1NLhrs3nitJdHb7sgKjPSSgmBgmOm1Cpl+lkfA1Oi
XQk20t3VUQS8Oz3IymSbfQEJ9SotrjkDGva9f46EV9jfrAA7xl/rF3Ttu58/cIUX
HhHeYjOWR9cTRCgZ5FM5achTSe5Umibss3Bq3Y+RwZiYJU2lVaL9PYFIw/rxt2QA
ImwCYjGY2LU7Md8olst9ArmTh92CkhxQNgIWbBPt2msjjjFwM0dF7Xa96/yS/Fjg
k+UdyZNBp8nCa2Yn/iVv4aylAfZcjldNlMlBrbNEUlfe6KNVaTcjxhZUY8kReZyh
gSwfV0uY24Ui5m8wJ5gyPpS/u2mYA8z+qRM+ynd4MUp8z1Pu2YMUEuO29UgNmwmX
c/I7Agn8REYtgRud2F4JtK8r1ZJwntxPUG5+sJhLlM/p38SiMJ/wDF09p15VYS9k
RdboQ6XJnR1y083sE6+H2EXP2/12xGDXKX+fK9BFK28GVCHb6ye+2AoSVn4jjpyY
rIRHSXqD+4hLtjP9c7LYmlgHkYma/ahvgt7NF8hKrUcXQJktMw2hbCv61CDQzT36
LkCPvPEVS2qPy2XbwRrRoK9JluCaSoY8r9H0HRpwiBnMpHpyVn7Zrko1B/JEcr80
wgP0XVMzoYKxzka/A/B7meW8FXx1tjENfzxEiGxVJiSKptSOaz3k5uIGCobmKLRV
x3kqXw3/Y6iW/fnitT/PDwARdN5kwLV+A79D1p9XuTruCMY8bOWlKjMRo2O/ZIUh
kCKP3vG2vIDJvZwHUPhqkmkC54ybqeDA/a2bE97zo0I4pAh3dvbguh3ONpDoqKgm
SybkvXXtH08LojXIMblpXD3f96zdsOvrJOBZsmc8G5FBjuRgdAWMDDN53w/853iQ
aOekDFpaGYJ4P0JxbcBojccE/ED8Fmx5M+iOVStnXtWmh41x7+9ycNuAmtOKrPIZ
BknuMYmS9IP17Jn7K4BkFXbM9HnWo0kFGaWRvU0jAg5lzWlGYxMPNurk/cVZcUnw
ZLQAedih+BLz7ruMtnMBdeH0N3RQcu24hXPFpKnbnfj4Kt72TecrYW8Qhd928eW7
AegYFk/dCWkFVXXsANs8HUx4fK2TXdi+AJO3OTGmd5IZrbzrZUWQqepEGJC30Fj0
pCjwuphVtlgz71L73mV8Qxc3xIm7c7NqMA5zdl3fL67bKa2HlT5PiSH5I8fAeA61
Fa2EMYjD+8F8cii9/E08RrG89W7lmQgHS/BQSqAbyl9LgL2OnzXo9ITBKnow6ZSk
/l0NsO6umHvlUxR3j4Qf49QbIL/D9TRamEVQG/29/vCJY7MhiqbgvVhY2KBBkK43
M8XZZiI6LQf4ghg45jqsKY4Q1K7oVr5NwfTb/FZOmoQVX+ftmj49dFBTTJ8wGrqe
UHt4htPZ4oL7MQAPJSYsHkBDCP/Q5GNSRAANSI4xL55tLvjqhnzoP16jHILKSJBQ
B0sBG9QASpw6e7j3yQ/QCmnnmkLjFloYko3HoSuFAqDsY+gBfT+S/HzmO+URb7wV
XKx54OcmC6EiKFA/L+Pl98CCCiFXQ72QgDYNSMnB7R7TBQvYa1LOjLs3JYfGvA95
jxCEZyavbvzxTsJa8Kvdlr9h26UW1ned5dS+xs9xHcLN/KhnkQhQjjcD2bRVjDDR
7GkkIa9UaR62koyFfs5s+LKu6D8fuUSNrrYV6mNiAbgULRQAxEtu05xy9v1EFASu
rrmvTo+Z7MKrppc+NyEkDQC+BiDNP+zwvKPTia83tIm0XFCsQBpLMEktD1FHdwWT
WowGBSoMC2tAKN4D1nkh5ELNh07V/dgDFYcJDD19qJvSfuW/tO6tl52ut9UEeSU/
mffqbl3poiNr6VBulJdpmm94ZJwx0r5pxWhy/geY1iTifsXr9q0qfvPb/u2NYYRy
U6Wn4j3tbtCvVoZJnJjkjbL05aijIU7FDBOpE2c618gq/GXFKqosDr3Hwu+XQT0L
FtYpNznRZC7Sg3jKxIT4qBvZ4aD/+7cLBKmFWQ0mOSIr5H+kG+MCEuN6WtQdWllI
6kL5vKpNHeudSfUNOrl2gCpeIJcutu+bzKsT8NF9k13Br1jQURde2Ds5WhWedp/s
rH6LeXPsbIncGHzq8ZymOqC7Cl410ld0mit/zWhEVo/DyNBKQpXYXtnoPD8+WiHq
VaLdk3rIX4kCY0D3BikheeZ5fjjEUFrldW5V92hoR244o1A5+qGr8QcdXHNkA9Gd
wj8UpOOqHuW7H7i1FcHsbYMUngEOShqaTH2tM+v5KCy2LpXqrZMeyHjL9/2FO+uj
uEt0dMaRHCvwpCFZyXuM0pdExc3vl/srn5NBfc5OsCOsKXRy76rd4QWbBWwrT22+
AmBDqKAq1V5by4j2K5ywjDFIgYlf0lhe8EbQeRlb4YyQfxRUCBZaRC6jAzvz2Tvk
Mki5N/ZNr+VlSbsB9kuW3H+kuOtTUTQFRf3axnAUMLuEplen68BRd2SBenPCziI3
2MEwcmQn9Sf/6QgdQ7iDEavz+lbfp+QIh+OEt4kH6kjCsnspPaMkcxO/hOxx2SSY
WwNxoW6c12OXtL94t20Rd8VLKHAY5Nrzl1MsqkfiTiDidNb4G4g1M4dxvwRpBUFp
Q8ogJanJ2e8UoLTbr6LgXaJdHQ1polLMFY0ReL15nMfjbP3Dimqh5zoq27HRqjaB
SeGOYnTu2vXYQX2kidvbRNUCsKqfB671brFvBH0fWJHpBSozOWZSSdvqiJTw9bdA
PV2Br7z8c/5wUEkkOgrDaDuk5u2/wUzV1Vx74IY7rlaEV4HdvCt2DQL/5RLmKpET
jEyF5I3WASCRotqg99OcYHdLH6psWqiTe9QdJCRrgJ1hiNAxh4sDqhu+LQ1HWo/t
geDQAsQ7pHjjsnj8BUfpRTBOE5MOlVX8u8lL0/PO5ncmGUT8lLXxNe5vYZR3sZcq
UywnoD6GkUmoeUrNL6nS2ZwzpFt/l1DrYO2VYtXPz7lUqKRqlWGuiNEPUfMXVIPQ
AN37Xkhb+xzYAGKmV+CsOdy83EBHUDiRZzpUW9LyNHWgK9gZxIYKm1KJtsIqv1ft
oXNOBs7pz6aRwSAneesTtdCD2/h+mn0PZMROiV5ayNGRSKGgZaAAn+VrS0DwUWSV
tlZW1ZN7eSmy+kUCdpBYjeGe2R+GmMttPNkKqux/oYu3yzJHQGsaCofbZLQrgm0Z
Ik5d4M70NjFDvU4m13nEt+FA6woQnAzoFdl9MbSzLIi99t+yhG7qu1+QWiMSCVKq
xRY7j4stbBFauDCdGwa8Sn2YjsQzZHSi25eRPMl3E6RMbfWGE3oQeZMlMyo4PF/7
19s5671g68ZrwEI1xr/jt+xvha0EgWVk1CZmHsUFgU9HIHCM6lWQj8JkbcWof6s4
uj4mwfqKyvhrB3P/T6vhBtFyHGi1k+o2ZZw31j58+U0u2aBMzkCfLMhKousBi8tL
3QQcdDesmeIrGKX/X/DX8TQxxDIfsksZICJsnjhjcUGgOmoCa21KvqlZs0G/3Pt/
CIQeFh+pSq0hvQEaIG98haC5HGa9Mo01la+FoYvfZMfXcUj+nqMKKw4VIkUjS0YC
sUpmoVoJy0FM79WVPMX/QahlHG/S9vuRUubJPy5WBUrreVflBYYZqigqMQfwNuL9
5Xewx+oqoMsTDqXBQ4a5dcaGwv0RsbzpfViCZKI6+BP+KsMzGe3Jymr4g9pfVDQu
nW0zg8vBmcAHJe0N1cEhg0m14rX7D1XaqRYwtLOYKqfnuz3TJrC2Ih69PbTXrOlg
0beDUt3IKhxKRkisH+NhCx6jy07IH7RHZ0eRDPlo8ZLM+uZxIXVHs+Wy9DFJ5Hv5
OAMIT6r+cNvTVSA5u2nOmTdfvq624N0vzA2F8+4T17V7Y27kJpz2BydduWtO2krr
F+2OYgyWnh69evijI50BL6f5IU0dFFP1caGx4gLLKz4nj+k6Vu3z39zqimmogmOW
zgumNBc+fWd8QGhnyzPSS4IjvSyUXdEJqp2G7tQSjC5jG68HM8lT3k8tRx3pRp1O
r8tQOaq0gbwYC4Ibc27Kffmg9+rL8dHi/ddiIgrtOS7F9oN7xDj991HJzdGZ1boL
KAT0IdHSE6PwZ4kGdCki0w8Duo7c2FwSUD/Fot1hox1awGdoZsWlANo8oWJG7XuR
sX9aUk9Z+msc61DWZbojELVN+I3IKnaG3zfHzvDSKJSNrrl5KCJYIgIMQIUuzgYb
24v9V5rfyth+cNhlFiGsOYrQI9vJIvsguSnaudfhejHsEevDboXj9wKZkr9GCU1l
JelUGX4LlJZCc/dGQbbSqr15ayo1lEBf6DJFU9wwlh4AZiqoKFtTnkZJQRzpubmG
LT0iEyBu115n8EApKE9XxQdZrnXnswpzQFsLRbwCH5QOD8psIyBU+VF/loCL4ef6
T7DcT8A7XjZwfIZ9eqdYrj4QBmB4jHwugyEC2zCr+Qt8/yCbwjKrnnuiFjrnjqlL
F5lHuBKUJyVf3o0a/wMdSAWfIiV/nG12FV3f9IA1mb0Qz4yy92sJLJxmj8+RMz62
yh/OuwccKi1FmOpsORCN8uBmRo6Gy2xc/MrfIDGolD4zHvIyd3V9jgUMN9HlKKFr
uSOrwJNvuTnZnjq0zdxPgYFVJi2PDhPag87kJ1OXAJGfrcDz3IMeGUcReH7w0Nc/
rpZBsw1ClqYxXpCSGUWabj+rNjqMhA0QrGxebibBiG36dAg82Cpp/lY+8Wvvk+Rv
DXwaV+1Bp2X62iqfd1sG4+erIUmthp5ZGSyQ/kDKXLicElpcj55oRY1z6+vH2cbh
QKMnERI0l6Ug+fQmgbfuuLoyBObWeLSHEy6lbl5AQ//ojeLS8GSuwuU/qVb1+cD0
wcLfz6d/RaULUnApqa/YJsOknHowLikyCLfFHyYHRNTORuUxaV9qcKp5bFsgTzMy
xBihg58YHdGC8emOiycMDuKaYCltEwdzoe3qxLMcyHHnUSLhIg0AsOZHy//c8rc2
zrp4WZTby7O9yWCE2mmu3SUjkDxlM2nv5JAy0l3Wf1xGItB0c81coa5ueoCWzETh
7zJhy5aP13mbvGrhQD2VtMC1v4QarYUC0PYWZHcCANsvuPtzxERRHLdpIhp7xqBR
VXCV2cYWwChBMSriRFKCJYly/axzLPvgj80PqNgVPzrz19UBnJynu1gX3965jVZI
392/7kbtvEt7/yUAxgmW+RWLhzJSH0ISLjpYXPKAzxLwb8QzIWnObt6zldbKNKMr
v1zeYsDOUHhCZAvWvvSjhOzuDiGUBrYSVF4LSd2I9NmQ+gLgH5evSkZIddvpwPCR
ynpboxe668OCxxxalJyxC4OEXpBkEhAq1OOhrJXthn/5scjnJCpz4P8+gB6dDcgy
Tuho+2KAgTJz01PGZzZdo1Fc63b7QMWEdxD3IXxddFfnB7Aw4hakq9d5ktkhtdWh
w7hmSLj6ZV/BKbqyRqnp03lXQoKqUEf3jVz0DaKmTlwfSZV3yozlLKv5aeHmrHB4
O/VwZ0mMO6UWH4Gbg+tKLZMZnSv1Ytq2POeg7REqVYz/qxFQsXJBcpUNZn6Dm4Zx
uLM1o6C3j6WmTYetyGYUGG4VnCGcW1GBmpa5K7ccb2VtcYxoR/EDcJOrhjxnKKTX
HwGRqGxZm0KVY7wb0oZOIakxn22CaVT6yY9fsAKztSM9hj+ZVjn4G7lgMwCCZgOS
8ZCAJse8W6Yz/MXuSpbc92ljGk4aPAI0QaDjEIMssIRgluEZafm6SGdnHnRNyX5g
eqbIkKJJRH5GbmuvHurFEZC0v2CIbOe/X3B9MKsZkBMmp4fhxgcLYHFj1hwn635f
7EkfIlDAI8ZDuutkpsQcNKxtz2J/Vn4ovh8cC/bMHjblqwZ0MrV9toL/pnhN4YWE
MCoPj1uwUexE4dBMvfVOAgZdWTRJBLK35wPNIeA0u+jIW3N84QVJK9XVFlNvW0Nx
yELxQAuJDNL3sDku4ESsyCUPFdVeGtz251wY2D0ZgjkkTHo1jbv4gntWaHT6yG7N
38xqZdrV0oHunajjavlo5q7dbU7ijpOWbl7rZzHfGIMAfnvK++74plgawo70h6J/
kUdq85MEVK4i2GlrC9yn0T5KGJlJ3kqja9ui0y9M/nTwbs9nRp1DeRkOockDCerH
ZNAqUpvWW4ZVlsHoIkUs2DgQMD51k/d0/9jANiTT/i0TVhri036A0oSAqAHmTqQt
xLtxa0dAeDHok0A99mlqEqAy2qauX3Tvnbw0IomsTWAOzAH2dJkMGuyYr7GCceXp
+v/hWFpLn1r4MBnVzKGXeCmMR/hki4sTNqR69slS00zeBbWhaMZHw7CpMM+00GYN
iaai7Up2BTmfhqWLg8roPVpde3uwgbAFDTW67rAAdsixcx9rkp1kaG2Bs2j47Bok
722ej6gIUGWso0dWxr8wU8Qigae2f0769DonR0xlt1PNYfXQCgngZw6d75B2ePF5
94yozts5b9bFNSjyuK2Uxz2K1XM/yNA088ltdiuddbeoYB0ku5OVsf7EuE0QEE91
l9rSkTC0LtDITX8WaGqi2DFnwse6Vhxd2Joob0kU3kfS96xnx/HrTvoiUfFzKONc
maq2cUrDUxkz7DQIsQkCR265gF+a0r2ZgAEuL4CyRURKxkgMq4uX4INi90cv6Qbf
UBIwz3+Nhf5zqL1kxoCffzuxxYwasGyG/pdUvhSp3QlExPWgb/gPfA/GUOhbLUoO
G+ob3QXWmQKE7USg2kwuPdgxwh3hd/YaBJK9dycHxf25Dk+XcafYdlxnKu6n5vyq
ZbNhAzzjwH6YhVp/w1XqIprfCT5JVVNivep4lvhZo3oAuEXaB5wYkqO8cS2fm9GD
+vucjZ4dBVcWFP/fy5ypLyEpjd8fsUD4vWnxEy5xYfdIHbeu2RjLZ+Kj757ZaWrl
w+yHhc/CwqpghwQ09V6k5zAY5lhbMlH2umiVyvwLBQP4tHvILprf3E2xwC2euuZQ
/mKhmK31b8zalGHb/AT5teeDy8JMKqqLEURJf5Kjlmsl16ulmNHBMXswl8XibHkE
Bt8L/2x+F0TluMgejniIyvTMnAqS6GvoURB7eW10SzWPW0GgJZ7/eTFW+0ZW6W4U
YDBmHqkITCfDH8WcDhvSXgsxipxneEaEs2hDeoD2Wno6WCOIC3mp0bpkyOHYzxUF
OMvb8MgXq2rBoXPAKxGkLonHa6iYPzfcNJ1r3ZC3oiYwWqm151eprNsoRV4OQBJh
MG+T0sdROMkgIreaS6/gQdSQY6Lo72hfKLpSw/EWc48IfzQGhaER0QkXcMzQ4Eoa
dYwLoujs0IeRr9P8BU1NAEM/nEr+cO0dN5of5WP2mabbcbvQe7lY6tnDsZduJ+yI
4YB7RVd+qQcrMDr2n5ZqAcgKHSpk1rWl6emcSOKZYEvObKndhDuTf6dJEYMUHh2L
aPmj/JA22Az7L8mtkPs9MGJ2c/HymwCoy63fwiincdh+k7XECtDDXdfTwguMlw4E
4hc7D2gZrBTzscAY5hj49bwAjP6DQvgPohJ4cHeiIaCJ1ZFudLB6q98RZx/bDId+
BkBIDwE0KObxgkaxPb4I7d8GScuejR4zgustgmafbLnZ46Zfmxqh/C3jE3w5+pJe
cuYVkLemzbc8MVSV8tw2HXxXiXAGx4OJsw2DzWGoBn+MlpDSkmC4h6y1QrobU9Fh
ElQJOYqgKbHfxQ9AcYZbKDqGWt0ZCd3EB4hsLA6UCgyLG//5ZlYaevAOm368zlRa
W9ddFInW4cXgSDlRhyw9JTy9/1mFTcxiHNRiPTQoD9f/HHUjUeCOYxkZdznltcAl
yNsRoX0WdO55gjoOyQMEQWZ5hN5QJAADUvue32MMDcyYiap0wRvQCjPWED224TJJ
DhZRRqAzSfFLFgnJ9g6WuDEYtLqzwacQgYcWwnplqWqsh/k6ccgakbZgXntZWstZ
z8LoyYpg+kW6NJSAmFsXGAQqw/poOHp3ha2HCXOQWVQR62aLnUjoDKBM8YWWQF4c
Q0lZNihNXslPIpWWm6+MsvLT9LEvRlI1OStFi3Fe3Xa6/0GKF48MDZgQiErJtCsd
8BGunXvcDkAOuYRIluOaxSCvrB8U4Tl8MimrCinMNS3jpOYnOBJTlavtNBchbshS
S/xNIqu+aWwsvYys5BqaZFoaTthhiZRmY5zHAuPUSWbc48Bg+QUxXi8Onlp/u/vx
xrbW6gfNxwBYMGm8tSZ+48vWA5szHABYhJK+8JNGDtsDiqZXi3iLTmTOAY6W1n8x
sGr4bRXmQHrcGtY9aVM6/O2eH3JsmWezWhCLiEO4BZE6n5rCDtvjBilV+c1wBmHc
sm/QxiUZszTr9Uxiv3gUTe75xaaPieUlrQcyoJlmk6r1KfZfCUJXiX4DAsLL/cEF
rxEHePWgiC3zEMvNF2hVeViYTUzKah/ViqwgYE0tvJuh52+6aC6X1djt93fi0lQ8
VLspSP3y9MovKxuD5eLD6ozju1GsSx0vVy73dCArFeQfp+iFaKfzW8QfzUduSrM5
68dyCt8heHOi4RvUsNPEyqzbSa/KnKpO4+r1AZl6egql9ZkVHBK5rzC6z3ytJqQ4
WYT5XdYYZwWDsoTdZUFkRswP5Qain/yDvjUVKCMycMxIW82Arjo+IoqJlhta/Am/
RzCmD/KkhsKSFpSMt07NEZN7YTBhbYNxS72uzJL69njJQuFYfqr2t9cEIsO78dcR
lZHVB3IICR34KM7pEfw5pVSKLXLpkh8zLYzq7o4iHBtb2uoZWv2coX52eZoQdrC7
/zGdKnX1g3ngMwjaPSdxgYxFC7BmNf9PGOcCTG1ruifrBVeukkvRObRKTlInfxsH
g9+75iZY2/hb60x+x3fDcMd2soD/2eYYy8KaB6ch9HNpcfgSid4471JRULlPxHLr
7pGeez2OgHKWWizv5kXu0B8clneqfbDUor64w/oam62ji0+Oi3wODqj41e/70Rcc
Ov37XmxSw8tr4bqtr4fxf1gxr/QX98/xxfp07DnWC7FwBjCe5WBX/sVbc7dp3muW
eKwGjlwtZATqks6sk9O6BvROJ+pfuixkUQTvFN9CrpK6C/j1jP34oIcu0ngj5nJE
TqdvdWr1VoW75VSZOspObAUaQcAL9Jbg9O2AmVXYJlhy3+dajj3aRDaq8RzREGap
/zR302gpdhagwmm5c5f3NrES9qiSum1TQbEVl2M+pmhEF3pj2uN9KTcE9kf2GEE8
EbVhABaMQ02dMKAjKssz07V5Q2XseomaIf6if8A/xrMjYfmV/tDBgJE4i2fIO1Zu
WbWo9DFxG8Ofxu3mpbRrlFv4i+siOpclcRKdahUCdUiJucdn0VnCtIJE0hRRF13Y
7k57tc8iVCc8+6mH02m3yn7Xe4eug4NgeYdkqECrbDitIyjtPxtDCsoXyKverBJp
PwyN+22F2L0f/GX8rvliilh4rcKytLylzMGQqVpozD9RBCNZkTdCrGGiZewZKMWz
R+y+ObX0+Whj3FjC4SzZrrYD3M8MUTByGbYFWUFaFF0QrvtRJEBmLSJj44v7qloy
/x644WvQyROyxB+c1buwAriIk5Zhbdr31W44ahOrq+UI/7z2yG0zEgY4DGSHoi+8
d+khG3xPnEBQtxlkAodSVcgFPyDr+w70R0vmKsZ+ms4ZOI+UAtM8P03s3gJrwc0j
ZL9pFM8DoDjxSZ5qOfDOewGV7Iaicis0xe00JGaTyaktwb2DTu3iPml/H79aVO8C
LLtawsEcFbLuX/0CUDE2we/ku81m3vPm8F47nNzUzVM239RpvpwXr6G1NNvgM/+j
pP5c8JJg2ZxI9QCTD1Oh7Quh0ZPw0DZ8MGbIzsUaCE/wWnCdgaMCdjacQmIw5D/e
o0ffWZEbNHlRARxah3z7BAsz1IMfBPw3u/GmCWwYBXhzJE4X5kboekn5OPGsTlD8
eWsWRTxAmI+52nMdgK5zKY7/cjtRpsLspcsXFXG4p/UkabD9+nSGqUkZYtyjIl1Q
oEo9oWk5O6oNwseC4TemL/l+uwTCSvakoJmkEdZ8uQT6rYx9+6WailDZWdFSCWUR
z+KgMD0sKE/oodl77u+pepL5LzpoiZkUXakAuTgOTnAuHwU1s2E9qI1AHTLcIW/0
p3NTicGM4NgRtrXKl4weaixFoamQWINFOTZcMeZrtVZCGIxno36O9G5x/aqq5adG
85ZrkFLKPMJ8LpNGc0cjY1hQDAo4+NyRBlCaBpDy0HkasnzMVQzNq4U0yUFlSVZL
tgKjQ20TCOMKpmSUEl3v7ePq/dmDfrvfXbZrL+dBA22kz8JzHOCC/Rzd+kBS+T4t
V6FLoM/O050exwMSrHaJD/u7b15XpCYEeOYT3VXQ7CpFE0GMvZAvvBUeYLXrPtsA
STChC4TefdZ9lWK8dxBpco/kqWTZgrezbZsn6mYRZfPjo60pMFrBapl0aafMadan
K2o1sEOp10fRLNharty8UD/kfC2pjZPHMrYiiglMrLdyYRRJpP68COvYUEg90pag
wzqv74ffEew7wjToz6UWNHWK/a40TW6UcOgsoaqSBQXSbmxrEFNZjN0uTVTqndD3
25DNC6pnRkR6rVnOCzv1R131KKiU8hlmnaMLA3N9KUla4O8e7K7zgHUbO5RnrTYF
Y3sbJcsyT5aNkiJYNXbMa5r8EUSiqo9jFQ+UkLySD3O/p5Y3fbRdEV9D76vYsH3M
fKuGNLoikCU/d4/nlDG3m6LynDdtrhgczKZ3Mghr+F5lKY/rEmAbLchTzmpQxrva
a65V7XMY47dP/AN7PeUXYlvdoIKF90LRpG3N79ANHSQd4hmcLz/ZBs5I+tTd/JaJ
Wf70VS5/fsAaFIXexYRoHxQD1VSOmR4coCAjWWSGdo5oGnlfE1Hdk4LsVeX+1ymL
pFHFTNVEGJoqkSanNOKNUlFEWtUu1Mgo9p7RGbuqIgp7SpuesvLXSw0/dnJvyTxa
3GKEqJCUOaapDg9hfCZ+xxRqKqOfEAnPCVyjF+9SWg5v1SUPTMQ7VnqEbjAU2X6v
cPRCQlQJdeA1amh92p1Ed8c+nhkExN0PdyM31dVSwLuVa4qLDX6Qg7qS6F7x67tn
aZHvjct9yW/o0sXWj3H5bw2iln1zz/P8LpgWi2MeercxNY9+BDx4MGDBbFu4Zr/w
wtnqDlpmIOK6NJ4Rt5PSVJLjcU8adnZzVG77u1+7+l21KPQKt0ZCFWFYiE7ExG/h
wZCstOu1MMAF7wcwLWicYlnBgXgjmhNl7hwHHzC6/EyqkhsjGlhPHMA4x0K7kLe8
4MyaizjHPFAZU37NAF6T30vj/MLp7qL/ZmG0ZRFay6uJ45tTjGTFd3VMNP1P0c+Z
RdqW7HrkBX+ytnh+KMsi/SwMNqjvHvWNelqJGh2feM2YCp8ngy8LbLu+9iGuPax8
atFlphI+J8iUqfbMMXYjX7/ttHiH2xHOlX0UiUQKXv8H/KkWirgrqwnAr07sZzMC
h3bpPbe3glBwMZUj7HNvfnOenFx7HTiWaFr3qBRSasCPel9YWcEvyqE9AIgTCbpd
xhoNWJpuvh5p7D7vGBTSLa5edBfpEbWCxpmvn87oyPGVkMfCvYlychBHdOwpXgND
taxd9T2GCCI10KYa1N3S+ZCpLPd3gTyjWYVYtWro5CD36h5v3jGTmm/YwSBtcLPm
j0xP7WNHpwRu3izOwY1wJql7xwa7DesO2Dam1Zhr1X0qsWQsgnC7pUMfzQnjV30B
3L/35/KPE1h7LuZvcpgvc4DZe+qWbYET7ONlNNOOBNoBcVxPVWjEeBhaNIMmYReV
974uBN5sScJrR8Z4vbPIxbJ+Vd9AlLKyBJDZcYjmHtxnmFNzl1hJ85AGliIXaCKq
VQl+wiW3+bL1LfymZvZBOijMVJmGMeOWyWhjqPC818Xm4RDKjLa5fZV7PlR3qOm0
Xfhz6VQod2+hhv0+IuY2LQz2lDUtlDflBrYR05UJgp/pRJzOp25CCrSTHkTdCrnV
GJkXKJRjFeYB7HxvSGV90uMj+Azv+ES2glF7CGwln7/6G7c2Zy36x/7REtCBPuq1
Utg+IKG3Ife/8ftiWfDyrysGiypVcDuFlk9AYshRS8wldAvuwgZ+ihN4qW4olDSy
QAtcpg1PnhGcPJ04jMO6k/iQkCD1zJU+BUKevRefm1pSVlnzitTu7C6xICiqMyxg
3ylMT4h2K27FQpYgj/2Dh8qj0OoxOLIoRxID/Co/n0rkokl7LRGmzUVzIjgFSeoA
gA+zSkc2ZpF8d1cgTsTvex3sIBRhHC2/ZMaz9wdV34kQKxtGUlePrs/wgp3ETVJk
C8FUuJIYMQmviOM39tjS/bK0wsbSu7ZT/yp4ZQaPyc/preyAqtSfYH24GhrtPlNq
yIwnyLTaJbzbNXoHyEInjdfCQbx455d9ulW30GOTcHfTUkazxOhhpdW0X2L5CQFu
UCUXq8UgRF22pbwINYmaFU2g+1mgAnVnS6oP5uQo/76K2+u9SssACKgYEWvK/gY0
g1ije/zyfTObM5N9JMNbqjTMdA/kiXDUTaDaRf7asue58ftcMSe+nfTyoxtGBrEA
d/CRnrktv9G6/cw0+2PzzPMV0ErzS2K75qrYBJcBrKEt4YZLZVDVjkv4fIgiJ4SC
TEESuf06W6lij8rk96kCWaQbnKHToXjovJQv7cjHaa4IU5L4v7gHfbQsUhqQFi4S
ORLZg6JUy/tiS19o2Foxh+f8SDaMPQnGGnua9r1APAhojB0HwYBGI+2SoZ9CII12
bewqqolspFeKr6fbhOxUGcTdTtyrLbeJGBoAyh4EdHd65NdJb3gf01/Md3p2junb
9M9RLTFaZVGsZXdJ5cmgzxQUcJY9TMnaeldHt1cwuVuj1HJjZ5ikUrsOiduqrHcS
CFfx4frPMhpCrYQCJO7MsqI8mEguV0gFLuloe1BQ4fceeL2EnvliYjF4feqKfPPU
SBArovQsR6Qq9NqoQAPGld0vccAqCaIADpjyfk7qDdyEAbVVb1s7O6Z9duHkVhQ0
b5MxBpZLh5UTwVdMct0lyWkWFFFPRBSGOuOfRWOM2cakehilNv7QM7Q8JD5hHvYo
sGYJr+I/qD8NBjFBBviCv6ON2EQBoDGyu6r6F2FzhzQF7XTJSxGuXlRfkNeWMwNV
vawr5Plcx7rhCPGmaps2i+z0g6XPkKQ1954vW209DcsBNbCDOv2Cszpz9LJMmyRl
MfpmiTHQScnwWfis8ZIGsvnUVA4/eu+l58qe46JAV3ajrJqC1eX4zg3Wlh/nvUu5
DaWbVDTmZJ1X0S8sx1F4WdaBpvn96ma9r9XbbeS3abkMA01uU+lJOx3Vm0UDX75L
qgt2JPpUv33KXz178V/PvNV5AuGMadQfYuu0o2b3+xWLBDD4YD8c1UDCOTV7FUcZ
tOxTkIydV1YsI8YPmj3dTsgP+KJ5BV/EOuIvgOjsV0GTA3w05OcThOIboIQitUiz
ed9w5h8JdlX58UOyGQn7VZcMD7EK7g5vfB35ziqiOel2FZCw+5MDkbnZzJC0Dp7j
kYamr+cBxv1MQwfAeXHRUDbx97TU6XksLcuY19N8MqBy3qhJgcPpNdRL9aeaqaVv
/rwntCOxZLg+kobMLaF1Kc0M9s+booCjCeM+AQGVas/r1eyPJ29o/ZErK1BgE47V
KhBoGqT50GP/rlBMV2WmEZq22ch0pkwJ9fPDMjC4cX/6zSfhzlbxyYGJNPkRB2f1
kXW8zw/KoEIhfeqx/So/WPunW1Neny57i7gc9RVrjMzc3bhtSxP+HAVQui6GvFVN
lWUaPACgPD0Rs4BF/o4QJStlJHjNKWPGeTXwEbDhPjsAXHFuJN3OTOqbkvFW0Ppf
LkfdyuMs7jxuCYdpBhMxQ8v1yU2rgFKEOviJiqbvgGmoCYnwrqEVqhR1uuqbAnDC
F4rjqLlnVERRlWeB4QFQHosD74xVsVBPIgzuJJCVWecn+BZ0+iIyD9rXkLY2PEDr
gaGpDliUTT61wgIGmM9QoqNDAMJf7rIK76Byq9TnU12CTF39cupIrxywyBOquful
txOpdnU+vpYUb7SVRrj+ccit4SepgMCXeZXnJHuIr9etK7BaCl/5shlV7HD1fudm
RvXb5+AJT74kpYp2fWrIXrS/nUsDg2/F655BKZAHfW2hqHNA1gkL1gGDozVVBoyd
oKoPJYW0TIWRNLRI8EZUXUiuemREnf5+kFBQ+kMij+Cb3XRn3o2SYq+hrLhwO5Ap
rCod98x6N34DWsJPldVzhH3bQE9q58IO0Cwx7UsmWk3Z6UxWD0bkL7koLiyXJjbh
qTlMik4qa9ZVXpRkEwu59HbFXjzVnDFZxD6XyBQ+2Jxcgb5TXcoks24D6E6MEwfW
flry9IdROi12L29GycceEyUadfRRzRNNGeW4QlZn+JxiP0JiHuhLoSQzIfx6QAWf
MjveVOS4zZIBsqSeCLbq68HaUg3UZGk9AAcikh6fXyuOJVJcZeCwsbGZUU+KQVdn
GwRu09ncUE5Av9oF5eIhKIaYMRt0LBno/BzWt2GWCyWqsVVqcQ0nCby78zCuFViI
BWlbLtxXdSnDpyD7wDFmJqHMyJX1b9Os5qBBUqZebmJ1Yep0kH9weGa6TxkGhcQO
0pNBEouV6vYwrxCjevOCwCiu9YDI6/SeSvOKSrvDAdCAIi8+mEnkgy/Y9UaHKiD7
1/hAOEYAbJuMpynYig/A5m+GPBdPQLpy298q1BY0Ksb2Tp++ZlSDG2/yV7Rz5jbs
z6qd45I+0a1yIdlhzDDvMC8X3fSnKeEW9qtrRjX8wIx+RHM/ZWZbFbZwdYaSMSHl
N9CS4ww/rF+eyKi6IWdJeaCuUK8Y5xuDV2q3D5BqZBFFCmH1GnNByU8o8KHxQY6j
l3hs1g0KlCoV9zY3s0lohHTxQyyVxhskV6L4MCwAcfobxXRoh+OFbkiGEsY0c9Y6
OcYi2kUsTBvV93g2t18kiQD0RMtO1roYq3UIYHFDMiCe8xe+S4htwSYOMo1LBLhD
iA4J80u/pZwksKPbncuTHNKoNhUcxkk22w/f3eq/tFtESU1eIZ4DNVjoVcrqbf9e
Cfd7sLeH7r3g2TZEaawTRxlGmhtevWdvgE+kV4oUjJaawNHONgHZBx64vFRGyKOP
yLUvywOW9BRpOifIMmkhVMV1DSn9fS9TD1DMn99FrHH0UtVsI9L90Pjx/tsHM0RR
cXqgAUq3fs1RF2xFGNrQTSur7NmjkpNuCatM/fbeXgL48UYA4DW5CKS7IfeFd0s4
CsnE0m3atX0UTj1wB0nOPgEs3gaqW9fqIXGmrRrpuWO0c+TVgvzRJNoFuFa/+XwU
u/cvgBamxH+i4RFr2ddGRo9h6tym7DIkPQgx1cZ6UDufnIT2sSyL/Pdt5Qd1ocCf
+a42CQ6gOJokX6aaFsLopmSKyrt+7nU6Lm2cnsAr1oizh9XBwvLbFSUQJpm4L41q
yZBockBOj3oYpGeRBZIQUrQmh8pndKBCxtK5hyIu66VXkcg3TN7rJb8zN74W9YZL
ht/WJLJlOrOGV3CZiffzlfHABWxcNg8WOer3mKgWgLbAI7uvtznsuchWZAinGBcC
47TNru3SjdS8iV2BbtS0H5mTYT4OqQyJ6BD8dliz+oQERFi5vncwnBn4FYUISBjQ
7VNMU0t+4dwRCP+/5xMUvmi/q1iq/384NpwHslc71y/DB8m94r57brT4+LF9LuDW
Qt5hEomTkZuW0QZ1uCpMOJ+9RhrgWO1Ly0tUthjm9T2JP9yEGmvBerGhoQDgQOGF
ng697QGFoXA1BF3GU90RcNO/pwP7+bzQSG2f9tS4gFtczsJyuKV861OzWXta+ABH
hw2Z21IXCaTNZ6Aemud8Wt96oet2m4QTawJwNONJrgDmOcVn5hFb9naM4ASoGAnr
GbMYQJpMH71JlygChRJZuidObSEqoo3Qef3M7fnuj36Cf9QEa//BHvnkmLk9xa9P
wSQHmJhySZRK0PjQoie0lGNJV9ZYjqhMrbQ/Lpujh7EgqA2UN6h++nw1QvEL+TMO
N0vG0LvU3RbSARf4jJffAavbS7yg1UiLQPyzoaZcipHbq8/UZrH0qlORFbwfdDGi
RRjodnUhE4X2KwwgkKYcOi865t37NyCJL1u53eV41g0/Zn+rGQH1R9jFJHSVEfzY
UpUr956yVuyhlamMky4iKz+2lXmdnHGeX+OSM/GKDUyvv/G18YypQqHd97N56pq3
Y8dKOu8vBH3F0Z8iY20kgRobIX30QWgpVPdnOECyTOPN+rANjsFmu9xu3CzkUqk0
gmyqCJ20GKVo5oZEubkECjzFP4v8yQUKtZZ3l64nzKQwfIqDTc9Pa4/55dYnNqDG
suRaRDSsvWm5hCUEvKNQ+Lnpxy7HpEfU4M8KovO3qPDsKNHPbwEuiFvqggXr/mes
vZANNewIdtxo+Ym40OLrjoEq4w5AslL+/lgDXNT7iQgoK94uHr2dZBorVvcI4WlF
/BcsKe/tfyNGeqb1Oz1XW0z3jWUed+mihPHmr7JGTNWC/CNs80u8PlqjkEn6LwFN
fgaJ12f8k6elp2GeM1ypNZ2RUgjzO0DMdRsW7Nn8Ga/hEU6HhZRVVWECwaW03T8i
2mYiNPZueJFeOZ29xqMDPwDyjAPkKOWmB5KcWufkU15/Z2MGj9K1gYqTS67qJjiR
x0QEdVCpNbgdmSg4/J1N/+pGkB9CgFYmZq9SUIz1I/hAy+dx8LMTFEWDJSGmrJnV
Zs97u8i1NCGFAIceWcovxuwaWkB1Qzx4uOhihe3SVyJS8LIILyPpePp31H/Gtvdh
707l7cdX9VjZAk+Y7RURffstZZ0GWHx06zzyKPh6VvcH77AvMAjTEABl3qgQBisd
p6JeEKT/Nt9/CPx3UwZ4bEefjzYpMC0IYlXqa2zKLoLY8cVBg59w0qlWR8+1kQBP
INlJwAG194GvlhuvtPPVq7iSYVr8iJ6iwwxQNojinPBH8rwKsQUCENhUiCGGqGhL
TbTbHas4Ru+eUxiFahCKbJW4YvC9rh3xl1AUPtrJ7HNXc3jc9cTPF2qR3Gd9ITam
qPWKzXV/doZkquOND+PDMdGY/l6FPURSvffi2GgixP8/N+rcCWYBq+OuLzlvHCNJ
GWTwc+NOnM0A81zd0ZgJtumUK0tQtnRbYQrfna4BHDEdhfQalpDZbac8N42FETSg
JQEbZJdzJIvTO13RuhLgCr3P6y3JEFx7vyUOg8ojRbuQugxkqzfQmUyJ3svR+ofn
YRXpac/PjkCe2QltWhw2f5O+90ZHq8qT7kfLV5zJZe1JsijGhsbh9RODqmMqlayh
QPDhenv83xhIAYT23URgYKGm4RdxgPD9BW7+b6WBKVTtYI2EldVKsN7p0jlg0rN9
PnwVv2FD0EzwaGdIvx66/ea9H0iuVDxeLnWvlskR8n/qx21mq8ocqMUOu95OYolm
xVtKpyDdG2CtD0D6NA7UdsruLrtUKENszPc9U2QGjbWuuXgAkanxiQ0fuiswAEQi
PTxc8yrOYHSsRsWbQ4kINdaKPoOSbaDFoBi6g8ks0ZUvMHtIGizGRckBPNAIPsbh
+0fEcH107xYqJKiw2VuifqJtGIAkJKAS8KYDioOOEdYb4mboOOI3o3GzVnAJ9YcZ
0O+NzgRY+G/GP0ehxS7XLduXtQ+2HHpy8W17G8TajRIfGK9lgwcCVAuFyPLNRau+
bO8iMtsZzdneuN2PMI7L5LBEZiAX+QrwQP+hmOnb6TPpFRe6R76fUCJIxQ1CMa+5
6Nd7FORR/Q2Uygp/pwpzHH6+G8IZl4KoBVszVqz5rJEnZwxBsNskqF2hSGrJsxvY
WqBQxIiYpdX+cJxH/faa4X/kKDIFnlL+7LzAqfODOUcktg1KYHGI6GgcrtSzL+92
Si4/JvVEi0pWCUTVZ68OejoM041kweKWaVIq/bYIH3SxtkcbhyIRACxjQT45scLi
b6QqFBYgyugtklzM8DC2slj1o+0u2D8WZM7yMue9uPY8utwGnH7Sq2wn6DOHAtNr
jtKy1oZ2T5LOArLTloGOjk2EH4ZA1M4jPIMeiwClUz7VEpJEHfnqYi18sgnzH1BE
+7jPOU82sRf8UrKfJqOFPWUXtdNc5t/yMdINDdUwx9MuZXQkdscxufMkjOSBlGoA
KvhCUhhdb4dZizrU99h6aRYZuhpFc24pnBVd5Na0FBtLvR4xApN/cNpfGkZdqt7B
XiFpU1shp/MPB4xzn1Cr7z5OBhy7FJupaxV6LWp4cfnKopK2XmOMEb6CdSCJhMoL
h7eWvOE7XR9r/VvyuYkT4OkTwlJKqynDzVmdlC0X7EmrlDCRFvV7cMhkYUyS57bv
H9tHRLgS3RUh31O/dlKTFfrUssHECQ87hgOsy47hE6TcxDS7FTxO6MmJamJd+7hA
dtlyZMvUZCAxmtRFM/ViC4NUXZltz7CMne9gsCjPkO5ZryeZHRNtjYhAbqT0sLG3
1qcjRpR2vrRMQH8C0gYFMaMToojh3rtQczWPZA+VVAHBGQL6WvF6U5spkUFyY+XC
tMrMZDq77p3GLRMsy/opeNtYWB4fVrdUmYSe4SDiOIV+K+dYs5lYWnR7HWyW0qlJ
UdzA4cudDmxx5FQlnTIyPDJ+chrl918gJR8I7avrkJ/fIP61lPBR1RZFPA1D0bRJ
aZ6xWTJ+hpGcWMsbrAB7b4MPsZJwoX++T1kKk8BdCLbqhO8bKJe2DW69m8BVDwaI
s7CcevI8ZJHbC3ds8Kp/JuBlbypfCqWJ8qc0IXrp+pN6hm3tupupy7a1Z6eIwc/D
mZWB/26Kp2gA/B3/abZcENOnMJIxxv05UZuOP47MyW3AzHZdFt9lFQd4nKvvcOBh
lZYHbRvE4GSTma45PMcODBzgDUIQ01qbti2qcu7ld2Np4Z6+zo4pgOb5yi+ryXZK
eC3fCbfa0W7YDDI1ulu1TSUO4IFrVxv4336JoYn0oDmas7zO+8uKwztpBChUJAh8
enmhMn5/m/9o2ETvfjMM47H4qAVgtnwBSaRtpLgdVObixuet/j10tnCQ7lZOcw5A
SyOn8JmUxbskHjOek5b1xSDMKqwyLz/9mVWMukVOHZHvotDc364PowrXcepAu9R3
djjMUwIg4pkrmBAkWRKFBR5z2X9PscVt8dAeylLQsmgbiXfVNs7plK/y3qdlWWNp
9hwL21Itzr5ulHVrhArfV1bQTDaM2//Y8Lbo4ef7WYTtI4MpnQW4Btp7ql59yjbe
WHp8T0+z/HjsbTL0aRt6GR/3Cy7+gfBWi01YjjMPSyqF9C1J89gWcc8CzGFcEYYr
mUJNHOXB/34QoQaxEbFvGyxswVsxpyO2Rmb10N7XyU1qQJwZ+TeL27xYQoIg8GRL
aQCLYMe3EHrKIFI/DzZo+Ljez5y7pQMEX3w6HAmUlzTxnT3tFs+8ttPBDJV/lQln
jcmtcIDtcB+tCSzGse7PBJcNWW5zfrJgZCaCjMilt4In71JBSi+Rg5oyCTF+SkfK
n1d2KqyQxpFbSLjfoImV3BRb37iUSe+kroVItlrsvSexdysoW+Jkmx4ZPPq9qX7m
Eb9k2osLbHuVlZVOObJ8w2fSNZV4n8zfE9GDMzYJs0xZor6Nli0u6teOtePVyVmy
bC/60SKBGTZQY1GXuCgyYcEdlX6Xfhwx5BTJ50nGdkoZZnCb3vOSAX0hlxnsz18K
EDluwjH//HuthLuw6eQ2E92HRqyNjy7JrsIiuU/iA+bwWBPs4yy387Xg0In3nIcH
z6WyaymAVzaDaG3SNU/3NLEf/n6laKn8yRQfvAuIZasJAeRHdJOC9rfRk4bYm1oZ
+1FCOikfhWB09d6LBcM6IqTFoHruD6fMrfNGoylB8WYFQWwps76m3yEcP/70xiUM
UenJAZKCvxzc3fiDL7F7gTe6AykGNY6mnjS/vxlrnHupM1zbRPRkNQNjj2ooehs1
LUQrvvCjTuu2osgK0Lu//nvYC36VWwOMZmn1p2S0va85eaUa0QUzImvRr+Jpif2Q
bNFoy0lg0zHKDWPtstfrXkZBdMuzhDS/Sc/u6pug1pL3SPX/WYiZ7Zxp9Zur7sly
xUxSnp/cssxV3KgYfpLHdnRfRl6X4HTA81jtb1GmDJuSlqTrWCumuWrnJ8HiYrmF
rr9OO7SOusyjQoD/R7sDiBq5LOaVwa3bATzRdVvocM8DR138AJLN4aQJMnKPwx9y
Hc+VipIijY1q3H+jn10fkwKeAs8llU57jgFG20HWQDPNDoVFkyxk8TdzkyyP8YRX
unGWQEPQTjKqK4mbuQkiq/ZuLFQ/7pR1W8CewiWr1q5zJKpCls6D2MvAfVa7FWlL
zyOaQeAafdJMuL4xmJS4NilyTJCay577t7pOWxIohEXvXghH3FFVpMRoVaoHjtFi
Y4RoV8C68xD0F6ftuGGMXEXIRxX0YPSUC4z787Jz0zt00/QSkjEJyurZzM77le3n
c8giZrfjByca0ZDLV0TaEpVF5J2itcggnwOifq0CVa9SFjl7Q2iY4vpjABguYhUX
AyTjJznUiqmuVCnEVY1vgin+ToSCYHNrA1YsGn547i+xjOWUy7OX2ylQURQN3HMV
hSYOhAWOdnS4a8XGNJA/0PydvUSXCOfR3zO08hf4yUWPg+nEcVBIEQKiT7uRn+Hg
cgX2Xb4KBGBI66gKJsU7tERit0xKRtt1+iBrjsGeCDunzXu7WuOBgwuV+JRVDL06
6BJSHr+F+sbQWwO4ToptpgQAMfi7QqvvQjKinXawybZg/bB/bZDBET58J+i67fly
UT02SN7o6D1yvyd3dK1H+9AH9rcMMMY+Uz4vR1xhVTzr35VB8ayVjHTrWiabcRzF
/gIqQv8xQCF9s4dwAkcqUIut6PMC4knblkeRsVRsmoZP98YBu4DDBh6lwUoauZHE
JgWPIwWawovLsiZivGACRPxR5+gk+sXyH88PTMyRTn/fzcVPaiZuctnInk7XjHPp
jJ2vUyePRw5Um41b1WUAqsEXkG1+hGYxGDj4a9LCnXN4ELpr1UI3JQAOVSz+Bgoz
3AyNTiYM2qpUlf4OvDVzcYNEmGiP2IzJECdqswHNipElrfh3cK8+QwVx6l5DttQh
2VA1s1/BaaKLYSH6TthxYP0HCSCfMg8bB7yiQ1vGyMDqqHXxkxMQn2euA4T56VS/
cxClbZTKjw3N8gMwYN/FhXMUOk/Zv8XHxhrBn8VNGfukUFoegbKpDIAt+qx3wqwv
8u2u5EEFk06yAmi2l3otTvpn02ZpJAL5g2aVWsITpnqGgRjUgCUtLiSk8l4IBRB0
H0N4jYjIAxDiTOj9Ylka+0cFUhthlYV1DhmTR+CMvo2xDDhX8kqvvWZKfHQ9Ihag
r5HCsJ4Sr4RfWf9Pki5K4tANv48daxNf0nyGCbnOh3ObgEhenH1ev/7woLcEz1WN
yP/6ogeDyJjFoPp3IgvyWPyY5XLcrYbSY5iecYRfdykYX4YCuSPMMb0QxWOAH3re
D0GRulcCm++8E+z9HLL78ggX8D06o+aBcDOs+QwKx67F4spm+XyIEl6KbarM4ipR
nA3ZwlgizwdfcUAoJePuCZgPNgpFmiND4udWNgg4w0qgI7iPQajm5B8DZLwJpWSs
vr/88hcXYiN2b81mTwSI6qJRy1n9teCwmXvxVM+Av/ai9iN4yQno51DkyLmK05kE
w2jIGcyw1hZ4GwQYSB+ce3AIARdUxbo/7Iqx6B2jyIeqXynydI0g3H+7+ByOr7Xt
01C5bnpU6Z/ac4xhsypCfFH5e3Y+zQzIeWXEZHdxpzEtQ7YS8KPD/pNiXObox99N
+28lkQgqJpZKsf4ZE4InyV2f2h1fkNVov+ubgR+xZvsrqPWvXZr5PqKzMWk+AzKJ
T0uihVMfkKhWX/Nn4STFCWt86xOQ5Dns3xfUOLdxvuKXfxnDTbi6J8Ry0c1q7RZa
14zYbpZ9RTXKVMXbDupso9FL2cc7wrvcEEwHQJIzdX6MFixC8sH+VhJ75r+GWu3E
2t0LGMVM706+VC76Vh/T5LnkKBBcB2Z4b399DN5FhlAEcreCtsrt9qFDD7QQdqo2
rn4UguqRNBh3IvnFKFnB0H6TwlPJMaglgZlJjhIKVZBe7tx62WUlZr+pHD4gjxZ7
aZgf5nL5xkMYV8W4wDM4ZqDGXhG6WIT5yEPhHnJeaycfjxSDYc0aVjAvtuCGUT1r
T6FPDjO9oJiYyh7SBUhT7vCnTbTWTO+Y/ZWYdu1Y8ub0D1ej3yl4P7RqVbpW8+Mb
3L9mvlejauMSm9XWSm91/N4XdTJfGcVHKUHSL6H/UWPbQhJzxRPzAv5YsqO8k427
RYjialK+2AE6SyHh9mOKLSpqIBqIWnaydGisBcx4KnemSlDOMCqFnl7/5ybRlVZa
OoRRkePYkXMYYC5EmXEZDV00BcGSInH8a9GUaNaYeY6Moyz48DQYs63bMdypRSfj
eIOLiQmRLSIKa1oU79okLV+tO7/BbnNCnZx3fAF97ULjHgdLnJOIgBm//XBOf9O9
kUAOMpY+8zs1Cc3a2+xkcH2ehucbnLfltoxGiBrSd1jBGuHCkn2nhDUsxFr8yXm4
AcQCj5FvuEaP2szpX+4biJ9K6t3OFqaSvfKTwIEobr/MACnScUytabT7h9JKCesr
5iNIoIX3FdDO6kMJyS17A/U6A0sKEnt+nB4+gpwDjIAMVdpfl/wJjU4mK92MSWcU
xfc3DPU0NAOODYzYlPLgwVeoN1JI5iddYLms9PKc5g9z69+M32Y5nJxTIW7z8kaa
Fnmo2o+jr8n1NO+xKOxvoDcBAZQfioPO4YpRytxf6Q+qclCNVWgrg3/5ZFXOZNpE
etW88LE8tnNh05Q+Ltj30Nj04TLDavzyp19IWVb9H7NlpIXSwCCXind+RHU0gWsx
0ox8HfBU/P3gqvDbGdeGtrV0uhrF945yQ8//O3rqzByn11cv/lMLdvmTL36dJ/SI
xZpaJn/6C4YmmQNM0w1GpNwGo9cA6ojnuc0njB9uGm76N+ANG6SVYAWZd/xK+CG5
y7CWju0s1Kq299FLk4IsK708AOQaeD+SSmqzpVJoPM0P3bU2oqTLUpfbMrKN1++z
jPLawQevx2DqZyvRBYdPyc6X2yap70oa32XyUs3Z/cIDOR5Dd6qbk7HwItziSzNF
tLQx5diGngcCyWPz4GUMHIrUp1n12qk+lYcKiBROPhlSHyHMsPZopoNM+hbah0Pa
4vDTeOETYiA+bK3W3lJIVr6Q4gzntXl2d8wI9GCRtg3CmS4t9Kw/nELaVbvvJ7+t
RfvwgI0lu/+AgwyRuhra3n6TMKBas2/Sw2g4gcWyWj85BEIo27NcKaTVkArYT1xq
eofcn+MwOirPe4M8IdTnZb61IZ5dXF5bfnO8mxtroGQN23EjMPGNwqAn+Y+1CKEo
gBk4SsUQwUobDRTe7Ofoh923vIntKJTGtzaB4jweM85sCWTHSXq1FbnjzgHg3obB
fKA21UQ3lLhAzCPOWVu4ebPqaUx2d4ZARWim7YnwV++6W3KgUGJdJb+fRRFPnyrY
FFWqaJU/OBNmF5oWMsyuRvPwvpko9DqSgo0T1/WZO/mRErNPEEjlAAugtsxuHilz
xR8fU1Lf782gvxS8s5S2lkaj8ow2Hjnow3/TFR2Stv6KuF41bLXkv3iRbryMxTm8
H+/aeKmemnMkhvpPNSxJ9pXoLWi8Gz+lTSzppHXyLZ+cxwmPz6bzopcwa62oBW5C
/cin83UAV4f/dzX7h4yECztom85TtDRgwZyQ8BLqGqwx/BCqG3al8l5tZn9S0haZ
GI4etHnQOJsO8/ClWTtl3Lzch9NiFsc8CZhJisjheFzOLuABB0Zwkk8kJ9Py8iwt
EH5rUa/HJdsaEUVASviAhjfU+GjVtwq8SKyNY9HkQizI7PtRPQQzh7AQ3qjYTIFk
KPFob3llgJxgpfbmglA1nVR2dZbP3gHW92NZILQfWJAOzHTYBBz8xw/BWPE6H1Ip
NNmc3pY4CyFx9kW2W+JszuJ7NBMmpiv05kaejVNxNfVcNTSa4SlQpfMu5jjqVqNE
IdeEGGc/Q5NTnu4hNDXj9rzh/6G+7YeS4xtsEzkNq5+bDI9cvELF4RVOIfj+FMc9
4XyzItsbTNlh0+CdOKLI6SNP6vz3RVVjZDNjH+D6IHUPK5ItfLGvN8TtXuaH+Zhn
/bcZqJOn0ySW81UqxihEzjpECKwOULHW2A1QAId68R8DIzt1/8Y0a2BhPFhLZZyP
6d8Kb3AhyVK1eJ+3bh8TdKLTkKEQNvBZOzSO2YPeGKvM7IPMmphtYItg/t+TY9tZ
AM7tvAeVNfiV3/+5k3OeK4p63oIzbYsDy7yJRIc8xs7NO1PBiotOarDWK56HFf4T
coTlburajqhxjifxnlguS1AoTGR/puJhg5FX+LvCcc8Zwa2lNzC0WbDzk9j0xJns
p+a3WzIGLcNEc6NXWNem6gx2HI/iysPHoSUE9EiZ/TFGkt+/MZGT7/mosCyNMtC3
Z7Ywg46A7pa88hrX555ZePhp+6FMPk12XRb2oRUIq3UzC3uOdZNRMKn1wCvwhGDG
/nI4Sg1iPWXSh61PBvSCUjDHO2jzeerI7EQUf1iI68JxDTXj+AZUqAO4dd+L0FCH
4EtVdfJPsrR0mJxG8dMygMmSD74Nu2fvWpAKNxaJNzYkBCTpmI6oPrUfqzULL64C
CEMEx0WF9GqrsK1gyZ+EOU1ecyL4W+IRUBJvvPWEpZzNyK1U2KCPCm4m6Iks5Z09
lcK25dBXjh7rLWfWOa8AWHT3Et9geD8VzIeUrfeIHBekM97q1Md0wrm4ugW5MnEv
ftK9rka+cVnXqGvlFNOpmJPPro4ZZjtWyydxlLPP9uLY1VFUxv79LTqmICel3d0w
sYmsEik2TgeUP+0PCqP2PDoF0gpbZ7X0nWR7n3f5Rv3dPMobWDydOOVfcsC5MHNy
2I1Pvehn3XO0KO5IeE3J9XBJknxJMjN0j7IBbQ6dRCtu2T2Ti/s6yRBFRxKKRd1V
WN+fxbLwmh0z1IqgsNvsVkJwUgcG4lLZNPtqaSDYjwOGFPVt9YVubJI/HFOTAyQ2
Ufwkrh0tj2k8+mvYsA8s0tMl+m3Kjas1gtPdYrvZwR95OtZkxq44snPVvybh5FHw
HTIO44cajyJmrBy2m9nkLMasNvppZ7eavxr9W5vuUYid6KaBPGW/dF9rq1Kn6RrQ
/9OWcbY8kCRxA38aO0GajiNTB9U1rOksRW1PzjFrEGiX+dwK0bBgi2Zef1UwWoWX
b3H/rjrXYf4fpTCp+3yGoAYvbs6AL/+8AUoOZs0Q0H22WCglTDsN9+BJNCpFUVaG
2WbhlmGKnzN1YIF2FvkdnQ6FU5HpIMstPDGZj5BCj6WZaauIshr/O9R9p7qgzG8R
xOZwmUeA17cY3VNeFDaGmwhhjwzIQgSU3OH8gIBuD1YeQsPvsY6VESxCrmSsXI8g
i4hxZH3eCsRFwmdQml+MV72C05p7xLg7wp8fjloXT0ZPcsNPIZtvC0Ju5whkKUnB
r1tiil4MQxr4c7j0Q/uQEz89ARcdgt8qSk3pZDpcAhAbMbXpoGhYd6TEgqJMPJ5x
5mqZHCMxeajv0jqvPladVYtkLHfZ5LiON5ZpKgXSQnitAGzdbbxbRqvBEN/hfXI2
224T0IYf3O9yK7+gE9TWkSrlQEt2jahEcsdHT5nQJttTXkCmJlTR8P1Sa2fF604z
v0dTAI+3pG1yEjN0DzJ3kvqASWzs7My4VcKCmoKa40l8E1qfMm6mE921EGZyLK+n
8cHzdn0O7KUpb52suIs2DY69hroeDlKRh5YT6zXBkfjOY6Y35t8svZBExHBj4M/d
FZQiW9OLykn8c1n81QX8ThtspVJgc+N3QvPGhHU7hhKtbtwQYGOBtwaCS7CRCBTE
CY0pIr8x59Tq5My3wbtACfs4q1nV/DTDY1wbJqQWIxx8XgmQiZaMYXkGof/37nVx
GpSyYL+1SlX3JJgBSgbcCMw0xGr6UunfyQYnBt+jfufs2s+qA05Im50nEeyAaynL
t5YeZKMvFJnMmvMM6kBj95Z9VkJXYYrVNJ8CLTkb/YeYI2P4PwG1KPuaGG0IClCO
wh7jQCcS7SM3rgTbGhD3SLUXyG/AD7EzTYa/4+BPKwYW152MRPaQRlAaD+M+nRTl
yTb/tuhoLIJ3O0EqoM5wSQEOJFG2baeRMftz6KdFTCTKiY3A7hYonZLNWbZKO4pC
5PWsMTYXaQ2yew4pt0X3T52MpkYCGV8BDYgpJcpBkRK3s36lXfY7Yr0OQzoeH4gP
BBV5rtmQvvX76ei64jA2VuZckMgUgVLhrB5JpRcnbCIv7yrS7yxFuVppIjxAY5Fj
g+pD9viUgI0kRW68vf4gBSgJz39RCHt2jD/6zjXbkQSMyjuPb7QYZk9dkd0Mrqdv
F9iWHPNkoBnQHtCKmPB2hL4MMIa+kd9eH7Zn2qmSeRCr/e6eoqgy276t3fphjXRt
5mbK62A9njuLRezmZ0XGyZxhRZEezXZFZb7LWUiJHzt0RA+Li/hU2BS3F/ZLoYDn
ZWtQaKW79CD+zvSkjJVAlwV2AypEYvRZnBbLytcWfPsmASqQaBQ8WaAvX9R1R5Hc
OBvj2YPN28jTV3pxhjqxr3JJxoTTMsInTzJnmBMZentQgfuC9kDHvOZwRQZxFXrp
z8SoRlyCJrtAkSkZ+NTVKU6rfnsWASVKOfas3jpbDnMZQRLFJUkP8RsqZuTqKHSJ
wyKwBxSGZi473ZsHCUKxCWo1IJ7HwvXSfZ/0vccjdY4AGjFHbcuxNss2E7UClD1v
HfMGxRAX/S7uooHxKnpwtx9sCqpCR/Jg4iyEss/5d7CUzLSvNfAP8H9jheAKClcL
r7uSJ0vIn4YdS3vHj1tszay0aCCCNMH3hNs2WyLPl6N8eU0UgNAl5ReCY9hcJevU
eRG+CLLxBiPpkS6C+DII4BTkz5PNo56533L/U1+Kv2P6KWaLNm8vX/0JXWHYA3hE
OssFuK0R4MJOh/qAcvkJQO2YOjvp8Q6mPcM9/q6jiCDw5rgTt6oIYIRgNeI9DzO+
5oS99LqRMD7HQl3p8nLT+eDe5228EcwhzE51tq67zltzMb4eVINJKaXMccAa06lR
/5Dqp76CMVhVx8goocTG0ocOWsQuLvaohH0ONkr9D8Qgnk040DdbQE6xvySaWF07
AL0W8za9+8zkChcBL1PIIwAGRbJL7zKuOt3iRa0YbO/0ESdtlJpm1OctP1KZCZTh
5eTtJy0HHzLDAN1aCdRZkiDNx+rtFM4PDZhM0lqII02+p+jqmEdTmly3xLAUBreX
5bvIo8HvSTYpIU5PktzUVL7cIrCrBAeCwOpAZKT7e1jV5ta4ldMJqOUu4NB4f8wW
Wz8EoYsMOkBoJqHb2Vtb9I3FdURYpMqyJiuQaXgmvXypt0VZ5TUCnAFv7cT4Q1iC
Rpk4NMgvAkIS2/FqcKDl1YTOs1eVJWsR+tWmYLdIChcG3UsuO1C9xfL5e7y8AtTX
u7oqq28GjDQjstnSDgUGCXcKMw1cZwt2018NznfCQkGQQyYNZU4ZoQz6GOT/NVem
3wSGcG65SetXd4rvAbLooufZe/pzLHD9B+V+BWqDhj0znIBX57tBAj4BGJrEJS9E
g8FQnJTtPeD1K9Y0k17maJXx4UasFD0ymBoeSkeH5MOYT1Ass/ir6QWHEwPtek/Y
XMj2tZtFspXptSQ4nvyfIrI+3AhQvot6Mu40makw9LctT+hOB1cXTjh1yGfTeSY7
MPdSnXrqdaUN5ryNjpvvFc9n3pF3sN93s9GRMnX9zPey9wm6tPWzMSwVeLRCxshU
ONancT5mWYh+8LoqjCYNxQIbd1mWvwl+gHkfbcIzeg4wQPH9CK0IuITKi6Z07O1X
nZzr/CdRA4b5u0/ZwL/VojXrI+l5c76odDi5lGgcRNqD1z//knFtdWSQFs4VzQ5I
2hXsEtfg26LAnQKC8PaJIoThh310k1LQqwY8ZQeLxcmFuMujLOF8gfu+j0U9FArf
0VY6+7HPY5P0qoliGDz50+T+E3stnU/QPNO4JckagEWFlWhv1Lh3TOEtUO4HoohS
DpXHKXDr3J7HsoSANuJxDbgQcn71Gifz8e3XWdeXwyw1j0xiDA4QLxqDQN4m49G1
xSkQut/gTJrfl9CHehopsWlget6jLqt8kno0sTjew93yDEyZ0xkapyiBNDkb4Iiz
V1kvXmBTRRFnUYwQtKElGTqsfG2bHLvllWm42rGY9iDjy6fEViNdkwaFWt2QqKK+
uI9IpP/ygVsk8+neHRML1qfLl2aV2JAhW0h9+Ae0Vb6xnQurE13b2a36ZIvom9Hm
7RSct7TwBdYzXaqG9O8DapfD9t8/d7u32NM1cE/fRxw3hLoZh74FQk/MyxgRg2uh
RD5/y7869uiwm6SYqN+hY8nCm0BPqcUWJjMRSwAles/FFXfMNbsfLmua7qWZqbff
6cUIpfzsK+UM0DvfeJni6apmXddvBcUh2h03fVYN+pA2HrIMqm2CtjtEEicLLzuh
n8bvKOdpRreP/UMGCzOkrODdYrYuKOAZchgrIUJfATz8WeqZcFcn2j5aEyvk8Fiz
tTqcLsQBeoxhrRnxvqjjcWauOMnCBR3K4FU3P7zaB9NfdPuaqnQT2MmfaxCfUEj2
MSb9KdkAVdb6GmgkkOhBn2A/mSkc9/hKA/pO5D260VpVzaDEGBjDbUUiMudUmIql
ymm2Bs9GMfJEJ8N0FQhcm31PdwVH4WctJgd1ewplsejPsQjFZbxPWVlq0w66wkaj
qnrevDbxlHp/jiAbHnH6udfAvq6bdmi4OBh1QU7itMS8RA09YzU5dwDR2zVkrUlJ
Y4lfZixiiJTzG1MiftegA+HpN7foYDv8zw3XRab92LG7EpXvw4bws4eXDQ5FZRyj
HDF0Q3KJ3uj2z2CzPk6GJNVPSPvmuxf5T6qYELqeMg3hveCfxOC9GqKYrNhyTh+K
fdZjkC1JDLkFEHLVOy886atKgnk+2e8S6YGqs5eU7FgbW6QnwWp0FsgxulSqCmXB
p13QHeB9JDBshohbjkillzkuLiJ/fkuUVHQlgv8SXMkaOlwY/0qar04HXpMy59ii
RI+0nE7U7q5BJdatG3kCAmglAc4aui42K0g0TWRu2axHLZKV8wl/CnNYr8by6n56
Nlp2rOJqvYe6d5bZifOa9hzfbsomS0UCNalhd5Tw3XHpjPt+en/hcPlPPMXrFUFp
RJVQYlZ2Ft1irCGWiFptawPIrmCKqc780DYNPV/yplwCMkzIutQI94+CDI8mcS4g
0eP9ZiNhMdNPXDz3pCEVegjyIphhoLwOYk9IG+EvHbhV2wa2pxwg7gpBPVOPqRrF
M5rs0EqpaZ9rrUGLlEw7CnOtqfpGjyEobVdHWayL6M0YWsAcCtBrA9lqkfJ7Qd2X
qk7dLUSWUKAYP/1Oinrjgwo0b1GHyVXTiqmBVfHA37jIbqeLDHJrH068M8SHwDio
Ry7d1Xzhz64wwKRXIXaSLy1kmi1Wz7M9bpl6pdoUS93/RJ6M+9/ZUXHroQha4n5R
Dk8IGQ5ZHdepIPNeNMRSp6ZmSJQgSjx3JjLN9l7379Um5xxMNhvUWteQBv0qXbPi
u2FmPKNDPKfl+Vufnduifif6RWyjH/WAOwhzwtOlbu3YkAnUZZyiX8PaqpJImDk2
iak0FKyh+I6mROkN+XoPM8v6fbh8LdwYFsMvjBEaCh5WtyeNpYnUn3CrI5/PYpry
ccIvFt/fbhTSt0rIgtjAFJdvfR22o3nGu8p8GEG5KqXzkB4NllaPjJPaaoL1TtTH
ei0XpiQLoiNsUv6iwsvRC3LskDMApEvvmRKFciMbyrhcrUj07Ua1fHzVxJRTIFyG
RW2LDYSU7wz9cu1b4ctUjW7BPKlBnWQoDY38N0SBDU4UF6KbdEzCsJbx7Z+yyyre
H1xamwEF+6zkkBNLkE0MZknw75Kj5Ji0m4ExZwT++97QHZnVtfME3msnpyCwHocb
hkmxI+ADU/lp45CgZVC6s8M//J3bTmIFV0yp8AQAtWS5X7+fiGd7nR+KZ27W0E9q
9t7p7t8OSUvalgqbVP7Uj4ddiVzTLdhRKaPfoNbE1h6W6/SIr/Lj79gXd/nmGiHC
ES3nuM1Sng9PLoOU78+eTfsW/7kjkUJxIjQYpHYMxnE/Efk8h56czEk0tmIujq4B
t18ed2BizOa47lgN/PVMdCWfhNFSBL1NfTFzIfDswpmmiFmbLQGqLQRpRnzuSg8O
BMGscaZCt57byk7f/DQsd84NNYsYFUgIJPyLfaMr/N2qmaVPJ/6+5/wNp7r2N3XS
StHgNMLxOlA5VTw8XT6/0+iqe0QH4K0NdfwlKaWlp6SFaFlw+d4J1v1pFWHOQPiu
arwgyQASpkhGlL0fh8d/YvJFd5g/B55Xv4rI5Az49IZ1YiuEEhvQMA5KTHDKVXZk
W4L7k+GxzfUTL6BDONpSlMiSP4RcMHb2EDTGH/1h6IiE0zXJqnKAqWi3/JRgynA+
N05/FFp5L5T23jlgqiSq2odXdbsHdia53tVF4Rq4xz/yD8+1sZqInN7XVrPVtYTC
Q/pNCg84jCspLa51q+v0pPtVvbDRHDZXrGqYHvt4IX2totAzv2YYN6l1KsDPK63M
5scYddYYiTtOJMahrKCCJJApWH1f4nzCmZdyy4UIFf0A86bZfk9SVd19zLRrfmAd
LzW6VkjDgY7xXTMS4WzoY5uGRo3BD915IHNXqYqlBPxJnkycfxl4rUjYuABH2c04
uZDribOatNMWvwvIqckCaCsfBjnF+55zAM8BJvJVy3NJfoAIfBlC7VrzHO2bqd0M
oxtL3PVLeDCAHeRrPBZmM0yfrHN2rHT7KYJGRQ5b8gnpZG/UkA4GfQfVE/8o8Hj2
54j5md18PF4jQ91UskTncoqQN63V17dRlO0F+5OOTqdJmjVSCloZoWkbj6hiYM4D
ZsnE+OvMR8U0lp0sh8ODCFZb5LU3IOR5kmjDx7Di515Rs5O7LExfWX2eeB5xtwcp
2p6i0/cdi5PnVDqrvzE9IQvhYTGEf/xZ2YA04uba+Dxeq8kICcUnkmR5Q8xqXQu1
r7mWJPQaBdV5aEYvY7VovupnwbLBB6A8astcJDHZ5nb5+nfjo9W2bFuNsVGxpYfN
W408KESNVuMCQwTizkDs3MWqB9VLGStdzfiDfhuR347q1GniAX9xdLOk2yZ1o6SW
E66PLY2thErdD+8Wl8kJS4o8qjsWyke8cckPOu6RKYGpx7RjA2e9EnWkzqXLWEPD
SJBxT3QQlyGOpRQZGQM4NgDM5zf8hh2ut2YK3IbSntK+BUdcZmEzYojG3SKVuY3K
fKjfK1k6AZlyO+h7nOnMtb9ANU4Q6qLpaWHxFrwkHLtFuafaqA1fY3NE95luxbw7
OIo5WeGwBBm7BJGDnQVPBjgdKyncV9wkYGYEnISmgONMr2m8fSpXfYb3WgCpitqR
CQiAkHv3KD8KNS4PP7ePiKSoDY2xmulWztE73EqETCY2AEFpD++JzmgmFuvkUMSh
bGT6952LrEqPo3gftofsf0aLbI+R0sACZPSOjQNzBJwoa2ExuwlBC4XIisQdL7v7
w+IwqgN5qNgHjf4fZaiEyo5pnUctxFQQayBqT/QeWlL6wH/VxV2XcJpcjH+rcC1S
Y7zHYNKQzFaQdJ361ZJmcbnMUnz3xCdQHSUEAF7gjfG4r0wenv04CUOq6RkoykfG
W+VkfOO5RoXGRshXl5Xnoi9fmuDyW72AhbNIH2YDStwGn00C6yUq7lrySiPmArLM
kTQz2Gs0frwzIWKs1b9kx9/vKgj78Z14EJ7DbnHakMl0hbf0u6TjS7P9ZPd8fNco
wujgsB3Ps45zG+ercU3eFJcDNA6WHl3iepu+zq19Y2Uhk6/1XHivxps0AjoqT9BG
NAe5sW8tnMsqclBF9RT+fx6w6hVWERpPUB6ubKVX0JcCWH56mdjpvnKOMk7K31Pq
12sK7EmkIIn86ql5YPgNvCcqAEVd15fOQy7xOaOYk330S4Uw5cjuGXTIBY1cafOY
ftwkQ18tq9Y1ixsL5Q2Khle/D2zst0t16Iw7y9N9iBzG2w/ra55l/KZW1IJHmsAo
JyF5yHECODkyO0G8Qc+aeVjPrNeZKVPsBpcW/iGTiAJzQ2s7DC3f6o1LtS2dSbyc
nIZEr9eseiQhsftO+rOsukehAh18b1dzHk74+SkokQUVfw6bE2iwYR3se0vcLFs8
doD5BGrSXY+171lo7v0sKB888LPzrl47U85jLuMqac8wZSeMUMOFQMDWfbQI4FRg
Ya7HS4ZFnEC6SbNN2CodSlxI0hNG/GTMBDkQk8IGf2YdjMouW7rz3nHJMmTZMcwb
jp2MkBWycwUpbUDIDcSGramlbsO6PGDLvVk2r3uw2BQJHNuKipTCxW1RAg0PC2+h
dJM9TBaXdDnl9GirulVoPKfpO7Kl15VIWrt40CBrS1doFHvKHjt1vS8DGfgpAsgk
xo+8/qGmcPczVA/WLwNCAMHFf8PzDfxMAtwOzB6gIrDDxgYso5fwsALLdy8p/o0c
bRBYoD0O5zhR1mLmhOfccMwlStFgrBzyNIli6riTA5xLL3MMgtkb5YXb+o1s2MUi
xZBFD6skP2s57xHJLp4OmjlBxD+wf3q9X9ytKOTw7eluao6s3UmadiH2g49xUOzX
kt4/xIk5DmzgvUnDIQkKqIQN7ghz0gcHPmoghE5LITscQ65cNxU8NR2umVaQkmu4
TzBaAt2uyeSNMT5Z92rCGPD9X8CnBd3qMcGCzn70awatiIDgxHypdjX/bcYobztl
yMgYYVMEawc7nTnslS/jM/gfCnYidan0K+V6BTn7gH7ffnr/3jT26/2VdvqUdy8X
O1z7iVYtojzyrELMzWwAxQ97Xi4f0u4B/gYxPuhkFGwPckKOq7cmHhBAecTr58Yc
dSVjjgDbESG56EPprzPAyhfjcNcigFSDWvHTdbNUmkpF7rAqr8lTIX+iEuZye9rw
F1eie2zUU5/bMQdBvtwk5HXHiCQm3sOWKaCFX4EYQYZUIHQqIxi3FyshsfRY8qNt
a92dryLrslThnIKiFch+QGM0pWTkX8tpxxmJK8er3gdYoepf7L+qicrxdfTbxDWM
jnugvLjjJIDvTTnItSHonAR7F+nN4PRDzlkKDxZPNJ51nFfAV8A/U4kDo7y3QOT/
ZmjO8qxUh+NOBCRxr3crpPP7xdX1JQu/1MuF4yMqHBn7EcltKn+k2UHASYk56iA1
424DWuDMKSf0Vd2qDa/L68Iv0UAVqZqbBP6NkIWXHusI3FUUTsZM9gCevnw0qf1w
qkz13Zk06iTCw2RpjJ29v+mgxPnDucZsF2H43kjYUlz78h0iRQO8LBENlZzeJ92a
o9PoyXDTtZR8/Dk1LA1L0wZchAH+ENlbhf59q2kqu8R9BfSvgPFJQ7mVmcFBQPjJ
zbtTMAguZfSj3x/jejR6Ki1qMEOLXd/YMGKFfRsugVewhbaYozzZ3uuZeG5FwpiH
6lISUx90amdn5nn1JmiSffhr+niZ66GKlX9PlhDIVw2wpOtX2GqL76eaJreDUaq0
hV2yBFas2VLO712vNAI6uG+6i87x8h/i9g3wtDxxQ6avbsdUISlSNNFL7lw1c/E9
/yhQcyxh+37ZBip2VZmgNYt4nWcmaU1Jg//N6fVVUXVdbFXt6rMtsBfw9zUf3pC7
WOiiHZKRmYz918qspHh93GxROiUTSrAES6hl2p0nPsFskZmY5E2+eZ+vxo5e7X96
0Kvn73dJNcpE6WoD7tBvD9DxbnpGC0zReY9ppCgSOnztw9/yKZenEkgz6L001LVx
dGeg7FE9jd99957rbPCkjTR1TtDK4+vBQ+7SZWqC/PMDd8/Gv9Qlm4FnZN5xAnvs
js3RLKtUPOiU3qhEVY9/ZuxGMQULrrqaywIlV7NgpSHme6Zn7rKOa/ncD/I6eWwl
ZRLQkT9vueRvpsbMm/raG7Fn5OMzPVnGcafCFvb4ay1SmDfkTvywBcyDbJOYys4g
wur9/UXtiVDwPcYbFk/fZoj92PovQnyM4td16qjp6xGQZg8euYvYI8JE5hwvbGUF
sXNByv7dTJGnTPRxu05Nt+u2L8jhki4laY6HUrNJiNhTf6KBtF/0++EnTwo1h4D/
tPP97wkNXBRzOSKHDmWD1aIXa75Q7SyWjf+dHKYnZ+SrkyKVMGQ9OUpfnA+8sfTL
WuxsO9+ia31paBdUJFy0+IZkEB+EepbiplyghPRuVD8vHXOpD0t8JhkYM5L7V/73
lTvGsObiNUmsHqNfSYPfWCyhoh0HdAGNcKNByRKalmKeqJVDwhN2qQXdWf3KzdvB
0eyD3URat/Z6yvm5iUSXoynB/DffKTBLMA4RV8UrPQGYXyQ464Ro6l1QaukV+60Y
YPmp8OOYz2Cp8FMednWldjSAc36jtsN4dAGfPA61yL/tlS9e1I2KcA/InlGJfI7n
m7zUssKqoV3pR+osRAIQ+ntDwlHYSmqYYijVaGCE3HTXDU4px5/9/f9Obof1F/+S
srNzJqrvBdoX2QgnKQaAccnffa1+0UPOsqTmCdTbP3mx6pPIc4rIBlgA/5IZ/qKr
SQa8P7ZzDoJxpAbmZPVd7RkVCBkFScKTnqpvprTdwieP2GD6ddLmitE1/kvpu7sC
QTCch81O13EUuaS64JUgOEpPHsrMGCPgvXIOIY0rw5hV1iloOjE4hTSddKuAO4+R
DDcng2Qqf5xJsuvuPK1mny9MPmQAhdwUMnGfnxpo2jrwX0nOXAdDH5K/Hy13yodo
URevBV564lPk9XYcp9/JkGyuMJkE75rzr+ZB6B7t2KZPQDakFJjkYpFzGibTMWW4
gXnIPmJEqGpwAE9t9Pits+zNr84fc82DqFcSBho2+/Pyv0qfEaRFkeurpTRASLZg
Snsi+xxQaTiemmvPifAtE4VdXS2h6mUYCJZTzdzt7Gvb86hWxFIJn8QPZI7zr3mk
GNDCRuHGpFTdCOJuyK+3bnmspjyS0hvTBUqk4Vt/OjpY35TpUwhmP60OcvuAlnHB
+GQwuLwD9EXZDeqpUqe6/AmNPazWWV2URwY3lS/E4aBLEPMsMVa0pkM8YQ6dbzjk
mii/Q3celYhSOSZi2AiqH9i+ukUhMpGIgZ84MpEvIwRdZX4Nw/pbHNOY1bS50zrK
mC7rkg6T/RVm1P5o2uKTVClYWdExi0yto52Ay70cuMuR5kfAUzPycY0VTCWOTc7B
zF3g+4rbYewFM37+GtM1giz8eEPLPcJiWbCch8MNjRx9aXt5jtwuOC9WoPgZKCEZ
MdiMyxMvLxSQN2SiRVf0YwhGcHNxzjHcRPrwg3gaiMpMfZKFgdp5cQu13Q3yB2Wq
snRH3RwXSs8dsyX7MU+Cid3mZzLpSBxmnzZQW0mF72LDbYLT6eFaNgOYwqRcXeTE
mymfqWB5SdOqAXK0LS0Vh0gn4F8lSQhUTd/z8T2gcerRpCh8IAC6oVIFnsYGqWwt
1COZFb45g0cvKbH3YNwGpD1qsgpAw9rL3r8h2McMVB0JRFQ/USxLM95/t7idmrBd
/MhVcHVYXCJnIYAbEXZNaU9FHNbQtKDTMognzi4WS1+YkV+51eFAlnV/5bKcRTqm
x8hV7aZBniO9aESHXnqHijrq4w+zDzeRYKpT4+RVgyfMITDcs8q27TMXpeLAnaY+
3oI8NfS7V8XBhYSbUbqF7vFd4e3OQY2+jN8qmrPPfPYg9LrqjoGS/MGqsFdfVLpK
8XTCR3L+CxpSMEpCzbaQh9SI5ZjTd7hF/6bWJloLuR5CxWoPfdYc2WL1eEdbgocc
2TBza4k2hSt7W4M5Q1qxhW7hjeI6PfPSkkI/wEQErcFBxtn6s0mLpa/hPNjDtH6+
IZqMCkgGUFJ7aKriIwdLjnj7Zq15cSDngFD2BbyuDkaX4H+IWfTU0F6TBzQ4hDMw
sLF4hlW5ZsrbYelmMVK69yFqVuru7NkZZuzTvexyCS4775Ay7kRNj7suR0lJrkVU
akTGfcBL25pnbaMH0ANwbvAK8f7mGn77Yn+Lh6cYlYgIuFjqRfqXoeeC0e9trcg0
cIex5QvnrLgw4ju3RdlJfW9oCDzkCAO3q7l7kIdHxJvjmdvLxUr6aNYWrli4pf/t
tvAaJDjYbIu8tpzsRlgpq9vfuckz8nbJZ5OUSt38rK1WnC4DItcFdyAtB0djwrBs
slrfwgQsue96k+ScRMxIwnQ0GB9Raun4GCqo66spwLfCTgAcCpQOinwqPpkNd9w4
cEfc9boM/MsGQQsDxSn2+eOSj6bYLojV7jM4XOigIvsdkNQ5cLM9Ez9lfrGfKgoL
xK4XDBucS7YxsOyPYj/BMO7Ncuz80UUd1DqSDKmKAgiCN6eAwYP81FKT7EIdOedz
/nh+z4XgwDn5s7EnSXPV722QueIWNK6S6T4vkuO+q6VNLVwCoEPIsVge+jL8os9Q
5TxwITI1bj098dFVcI17lzVWqTQgy63StgSL15Q5fl3Axa2Y/9qT5qsNIuy3ottT
O8a4XPvowEYe1MF7cFoi2+g+arfasfSDhk6pkKYo0hDIYm4n55U7Dp4LKlf7BHcG
e4qY20M0+krcWgAW9wxWtCN/YFkJazDRoVf0zb0HtG6Tej7n4noaEb1HyjeKaeKE
o4Yy6nEHZz6TWuvrSgPbq16Z7yvIpeCcAzfeZBX07X5gHyHeDkk0NyREJleCiRrS
/hjy79OSFU6yCh5TkQWZErjsx3IKIUfTKSbsO8dLv6dUenv83lZQAcxEv4GndxB/
33YAhrqVmBp6ItbqU6ITIoacr+N1fL39dtPSxyxKc2EAT4dfboxWBG/BMMDg/0d1
lnULDheEOfgSkkDPSDl/jWLrY5/1gBhiYRd+d3OAWFnawdNB/kWY2zD4CoPLGkti
jhp9zm91WJafbc93214TpRpJFkYitri+K3K1FeTAjtnXETP+tiYDuOOOeKT5ydgf
tGDNo90O0CVLCoR5iXMdLGHw0yw4JDzNTQMAEbU0QVwLgq9CN6zGzoE3e0EtNNST
9pkYkTxyTNxO4GS4+VJyOGGgonZmoubnxGE678G1O4KOitrkMrOd/3oaX7WYhvlc
pptDT9RQPt5XLMXE/fukKFUfpyx1sZNubZmzw9LvrYsvL7mz7AL+PVbrZ4JErgNm
fXzlTgYSwd3J+D5QBnXHkp7VTR4b5yhZJe+pbqGGYHCsJXrkbOapiWHvgeGage7/
6bN8HaR7jjqe7hN++/bajbJE6PDRwUPGru95a3DZsmB2VQ4Rsw/3Ll3ynK0PT1hX
LLi1151HILgB9JLw2BeDthX1eiSPmlDFlw3x+uOW5hoQ2BgN0FNQQx7DLluxMdqi
q7+NNCd5NiBSP5Bk2TNmUlO9Wjn7idSs20YgA/6crnemDK6sTLWoFOS8dObit2ok
jHXE1SBlokT+HmO1TE0PzM9XMrjDVhxc4UhKfJ9MIIx7mUubUzcuttAaPjcpLb17
1l9r/Am9X5RY3nq0bbWmS6OfST2hD9wNRl2r+YecPe+VHs3VcakdF3FnvuSvCd1Y
Wc5M0Jkqj0bS9Tdpfu3d8FR2K5kRnilglZUwy1uhFFGM0wkYOW/ZrBkKNFbhseZP
K94KqRC82aCTLPVYyFJRFdddbN6569AbkKehShHI/k6JBuKQo+CPIV74/qRwBCpf
98NdP7zIwRGsyOl8C/R/PIz/W7KO6khb+JotKfEk6Iy+tRXxsXSGZKshROv7YCu6
Uait+KrpKTidV3q2vX+VwL+A8TOUKzPnx6vyePQvUbdaiCWyTSU64e2B21cHYZwV
gCXiINjjiaHN8c/jWtr0JM3kEO3JsCn71LKhnLV6UtYeGGs03EvM/gNCCYzu19wk
+1RZ6eLUJyYRxl1BR1bU31ar9ek+mJighAHloBrNI3Nx10CCm/TcWle4TTmYj35/
aPWqvMxnrwLNJWHu7+ywFhOjTIx2ZgpwSibtl8msApVt2GebI1HhbfSdB4p98iBT
6XPmaodxtHGgYN+pEgAdALiTYj1e3ve3esFxXAX4N0AUptljcY6dVA313wcgllaU
WYYzqydzsNq1QiBT1ho3K08eWx3n0yrD7Y2VG1bhndiGW001ZWyvvCb7crY0U212
xDTh2H44/HzMWFDzvCMToHIlOQ0HDMLV6D+aMaX3K9lrH071BynSS7FaEwC4B8k6
x3fCS0d2RVfcODEqCxlzet3UCL89RPi33S3O63K5USEXdAtOsABR29VYe+wQLucU
R0TvSavMW0sY/MED3WDErP/tWvXKLP0+5R9QaCul1L/GCxEa6wfcfntrc9tZ7v1I
MbGvOrm0mPL5ujVOoqEVijKxht3wEQM8DRJO7cWdaX1tnffYsCzuiIF/PsJ2eapB
R/VwITTbYlSc7I3GKtnyaiJlsxpaGH2Xe5J/Gc2wE+EYQSD6KF9W9UV9mihWCYKV
gLlpu/rROm5I2tHq7kV+ojt0xq/7xLTHBZACpTjB67vop3VhomrdMI6KuUUENut4
1Nw9/vyF4mCn8gU9KRDHzRFptar+dXZXzuWW0jN8NDuKv6OLCq4AQm32SbNupD2a
rg13tMYlnvnwZWxI8hKbDGfTn4Iz5THKMIMP6dmxoTOywsH+JKbB/yOhg4qsNcDE
RUmZV/sBKYimrAOqQnGN7kVGni2eP4PEzLQklKWufFaKAVJBinP65J1rf3D5rbv6
eBgpczIlokrUF5Q/Cj/x+oPWp67g2ryttlZD0S/d1BIv0kSXgrhZRB2Uh1lrqlNu
apLsZlEnUXxKbpag/TnYARxfCPx2/A1jQW3AZBFy07/09NdsQQP13AlukgEVDHaS
mPcv04sC4HXsiz5YQOj5JWYBY72cgE5A7QHqHvaiKEXrv153hP2aYUqa66NwJCa5
T0nxCosnYGDIW24sUCfXaZKKe7UP0kN2TdwuGEQxj1wEKaM2c9R38GXD/WGs3Dgn
OHgdhJ13l7nARjm/Hj6E1z63EtXdUjmV0KH4qW4j3R9euBVClWzBd6VM6hPZccby
5JSrypyJxfyeRNjH1NMwqnFTRkABlMWI4MoxOrbyFmOWkNAMrKFOdDxJEHhXByRP
DHiC9fjm0elJhnXV38z0UFsTk9R6YWoolBhVfWVG/MI6du8NtL1x99eiZuvc9Lnw
bAqeXjlXV7ipFo1guREDfJzxUMz30RKVDDaEdrX9LgwckBlnBs8CSjjfqx8BV9mt
C0xSOOL26MZqY0D0Ij8PynPktJW9rv5kNSMiCKCRJ2fyRkB9ceJa61kmXUa7lwmj
CRYx+eNCWsAz+SjmuZEL34JgkLnspEPg7M3RnmF8HeXcvssvwSim7EUpSao/bKd5
fEbatxNQXu8PVdtvbrvoNnzXvgXrNXHOIxH4TylUHUlJ7a+TQr3UXVTPf0DMAjUN
bTlrShA5HQSF2FpZr27ewVvGR8idmC0ciGXKixGW8Q17NCCl4dHQoF3b4rEgP1Qr
G521skiasek3j+802HFL1yFJc4ZsVkPyQ1m8bKGAaI6PEjd6gAO7bcp3b8Sbbypn
ALwAeRfvZwtl0pMz5M+H53fYq+FhMxCjn1hGNAwGT0Sdk/ym7xmWQ6BCUSpLtd4G
fjNi1WCHz/MUohNIFesgsWVnTU6rAj5cVKPc0FVeQDFCbB/AOiAl1W12o4EuGT3f
uA+J8whQ5MVkU4mRkQ+SKwo6TOhvu8buKkd1YxyVtmC8v2/Y0PjOl7xpUZg+AK8q
Y3nqVe2re1rlalQJw9FIdzWtGRVVAkeZJV89tX4KeqfBn6fmWYoSzPXsVVrS9Wmv
b/xLbrxGnIxBRdzb217by+7kp81qjp1HASx6vapq/XMAT7ZtXpFJdK1jKg+nb8N4
oCNfQCX/EFZibAqRzqTRC8b+0vRjlVVoVgSYWlF1LBfQt75XV0v+vZDwclBpHDP4
Y6yEJi1T4hg4d7+WvPU7g+2spYXUt9RKd9iUPuwsW+ZIVEiuxchr/MwNcEFzCORF
0lTYzC/uxOrtrOG4N6tAmUx+ZAe5BQL3ZB7i0C+R4IJ6LAB2/V9TLK79aDdybFVE
J9iS5QIk1jiYYJ4yMTdXoz/l+LIJ23/z1B4GRqaQwWY0x+HMijnk/ZPm4aLptIFF
dcwjoq4wU9IbXGQPNBtABMOuJhs5MtzbIBgsWL38PGdc4m8FNruji7vj/0PCqcbW
Rr4CZxurFnY7Ri8Lg5FxDybsZGniBA5sUSmIO3PiXpqVwbg5uhpfv6x7lnsmjM5d
cNvkxJI/6SdNOaBoqYCd+pQjw+837OGzgFXt9Sx072ga3Xn85rKdLuYwG8qNANFq
WRxMQUlchjdpKTh5kQLgkhw/UADa6W4cUdoD9Dv6wnTLecTA2Pp5+MYkmqGAAMWw
PvBcx7isKXSYZGaOueE+ne7cqcg18VNVT/3/sM6fnmykOs0fFJiVHTRz6MSEr28Y
FDyVYDV5kTXkeFPNyZfnBztCWjW/RYNablaJBW6XmLr3wEn8FqakqSlJj+NA4vVb
mnXfuY9KhA0jqfmBBGk4KX+lu+tvjOOZrPEA4sw62dKpTJrW+8cvqmkH/SqA/9hL
ForLsfgr9OLjLNQAbWHvwM+x9o45QC7XCMlyRNl+CTn7PWSwa78JHAmvQksHwjGP
vA89skbpWaFdsDVvx3wcKm5RQhQIksqE0jwI18mqoTwPIdU+VJX03YiutBcUHRZY
8/PZzMLa2XKoH9eNXMSIY7sCIyXeGZbGcunYZ0yUbUhypcRa3RRZ/pcDmgB++t58
W6fCj/5v6SSupPejFaRuuobg+hwfyAnjk93DsXOurDqX2mTkGArznHbIbOI+jCG3
VIdyzDKb4lieJc8tiFr56k18ksDIQIQGiucBCclu+t7W+iESYFj4u0eXY3s9BzTj
2akbh/v77fLPFvMDfFNoZB5EMIBId1fJJIF/qh5bsV63pXry5BZQmnzb40HM622u
1H6wy+l/lNRHSO7saXNIVsVWS72PC2bBAPwZzPtoWLQXHvZlhrGUnGD+s93B++VY
MDmi8b7ANb3xNjUZ90r10ySVPYIUpYF+k+KOwzkagCoH9lOx3drLyl55MNG02+/c
SBOYiB7okfjFOYRdE112D7UG8i93EAV5mN7I2Sh1UiT98RoJCSO9sP7mth/4+7j4
+DwFDMIsmXwrRmPRcSgTUiy2R/a1h3XXJJkVd6AOKdVbbDrKXjUxzJreQhqS+a87
pifK2I/dpMvBt5Ac/txia+V0Z1fh5N6p/gUD8vj/8tV4PzvuqPE45dtV/h1aeUnf
LPga0zUVoymsBd6UQMQQjQ+Enm4mjRSCGNrKjx2uEKfYJMHtpaAF3or6TL+1y23G
ZDwZUF5gN6p51I0ZOm/T9T4D+274L3oPNOyRq0IPc8tFpSmXP0+s9pc3+u80GfKk
EM5noZzTXFC4v9vtTIB92grGtFzaiurjDarkEfuEwxa6xx1wLuhBl6HT9tvKI33T
S+BaihitoZ3dODGYr0bb8QrRYt3LFrMg1kEdA1S+0nUnWktya7m0RL8LyTZkwge+
NmRzX0JFU74O4Zps0PiDmDvEhByTJSspcWZ70dtzFmteNa+9zWYmkIhxuLvtvQM3
Pw2SeDaHVx+13+PuFS9o2ADQmUqz/ynE7P8bNq7DPJTqfv73ewAGPsyTT4ffbuSJ
sXWM8UPFRFuwAtdJAT3vwu7/FeHtptX+b158O1TZqjLLB4ct3BYfIEV9ZvY5RWjI
W5YGn5zxzV1HaCjRVvp3pAUA8iobK05s1bW49o2rqkW8Al2IV+Gb8kptf+tYiZC5
SCMFK1AdpxCxjENvz0UT2pZSGldDz2eh2TSI9m2iOBB8epyxne4wpMRsGC4OsUQm
OdCNK5CsiOrJRcHR3CGULwiwWVgPTkoYFeVYLJ1r2Ac3nvqYzD1+taZ2gkZjQW8u
udnPQsR5N6h6rsuiOTcwe2J31XRMUducYL3/MLOb0yagpAA5noyHeAHiK5RcnK3/
T7MF9UD0zdLFrnqizuffAJ59DdYP+H0homMHUcdCrD3hdsJ7GRCSA30PXF8sSa9Q
W0VBziez79ckXG5j8R18+uXEsb1xhxS2OvtyzkbnisMEq0Tns3nWB1VIlN/99N2O
0CXIOiTNF0jhtO1DiUZ7U1rTMIB9xv4Ba+/x70e7L55Z5LRdNTyDLbyfDrvO4rMg
W4lCLI5jVNonUUSPvtgfvNXckJdeZU5ON1d9/u9/2VYGepF5DGNfEUaCUDgCga37
mJRpLj4oIyZqvCqxn4z74HmEpruEfgs8LmyKgRSzPQ7OoFsP6L0ED3CBVtgR+B42
yvXDPqajz1Ai3R+6x4gDKLlTtpS5k8dQ2F+26IP2pV5GpLTQcY9/fipLcj0W2kjA
WuoGvPk4KY6kAIV5zyac67ekpjUp28ynO8VvXQYNP2vpSnbHQpum6/E1fjYtGYxS
RDZoAhOOhbQVxogHQ+M+iBx3o/yxSnGqD5DxydBjJBLGLl/Fk4OmLwETHuTBghQm
bFs4po77EmR7xP+s1aM5C2U65Fw3ZMge7Xmvc/5+OTejWwwuC3ud6QGdJ1hZdyR/
8TqWrJMmL86qt/rDoyFDrD4Sj41dHFJGKYlkcIzMIjHgU0qh1zzs+LRIhqvQTRq6
MGhkeA7fg7GkcvyXcE92wH0mVzZdGJXm8nFLCBG2u4/RoQ71enpbK0tgTuazC0MV
n+sYlre4vtuftGPzBgx2+H4da6plebIsi8WJN629E8KSGJVh6Ore+WDw/iHHqWQE
/LecyZO20ay2TxeF+m123YRUgd+pudr39BlLrFqn64RlFuMkKM3SfxWsnjzOoasw
x2ekOlIqV/b7GOHCgvL3rwB1Qov/y+xP+3L0IkZa47Dno9gJc/g1Vkrn24MvQkJ9
KVdhiKXRvWtvdvxPCBJD70796Pgk6GHZjIHEamz42Is/I+w6zmQIB+BUTxKqeFiJ
MXzDVdVzJnmrG8kw/6pSWwsgm5KXTsSJ+wyHyViVn75G52midW3nwHeZa+0q3BHN
qBUCBcEpnopHOteBSdPaeHOSpIrI7JggZHdBqx8hIP+edlvJdJP92u0tmXNbPnue
ldPS8TzhWtH+Y8xffcI+FbIXdbK45JOB4ybzGoAjMl6EZuML3tJTs/FScGHZ17/f
5MzwXDhOb0U+OuuN2Pbv3T1036MMkkNq1FpoL5/f19jIRvvCjN+uGIT5W7tr7SYi
bvH1d8doECCWsVXJRCyListq98vukmrhlxpRMngKRwWmoqXM/Dageiw+2+xHF/zu
jxgNVNcb66SAYgVWWiowxEXstGU4MBCuqvSQRB4t+0L4nFwJTwd7CWhb2eLbqPnY
iolzvj51S+TrNAift/+g/pijNS4snoLFOchfnkiTnmbYqX/vJc1rrvQ/Z8EjSkGf
HSKoCNxwZQDO1D8huXxzE/xAoOoETUnCg8JpfiR8dGZcFK2LoGsnK3/+DfxDMaom
cQAR8sNpl++HmLbibUmuM0L8H21uKB6soDPN0Jyc5udsL7GcDqMPAZMAAIgRizBd
7ehvuXA4265zH+LvGe2R0BOeweibPTRF3sjWSSXMc4OByO0o5DZLeGQZUSxKvrMv
Z51NWKvZEGfbqb+gTRCPJ03tgTb48LiiKWZML8a6We9T4YCprql92uwvmLuwH8mu
WTAfIkAz8W91J7IUUm/3Rax6qQy6vRWf51hZjk2eqAqkgK9LSMwdau7NZnuNLDJ3
XveSZFvcQcgAI8QeTpQ2ctC8tf/Z14rT/DtDNr/+94SP2s+zvgfpH3R4oWkjGju8
C+qauCiYYyKPCDa9gzME52I11zUPJxRkd8TkUg+vg++EisUbiSdX/WRDMQ5kkc3r
LMY+pZKQR+QMbVlgqKjR+k4uTrv7rOi5KR/Qh/E+f09WbowfiBKrJaYqiwk0GfpC
YZIjhoZDPlLsNH3L2MlsgTF1qjpyX9kvagY4xjZ06C7UKuIwIpGsNf66AGRL9m9/
6RYZ0ThMaP7UezLpFL9NVVGoF4xeFVSwPgwGfVOmXaaXrJgwii2hggf1T5p5ydtJ
gcrhuw2km4UUQEWqjxf/aw4ByrHcVqVOlXZ9k7YxLQCijEjNWo1VyDdCTLLO19d7
CZjTFWbfZx0dozzSvkesP/vyqubKrtUON+VOJHIRJhkpBKMuMJmFHyLo3nCgHS9c
HI6YLm2ZEfzRg5TArU536RsK5fbxaWuWLctunZYOEr7zvGf1HDPWlxP9ri0vvv+g
BhPyGBmtF5aufAqkPDNwSnoMt2HirTt0uVOlsuGVnfs94Tb+/DJYUqDkPcpt50ch
kmSUPidvAPfvZ59ep0TF0Y3KQ5eQ7A/oIXW+4YE929zmCelNmeXwaRX4TPd0A5jH
JRY3KhQjhfc7T1C02TfMo9BkpXtGcF7SqpAclXGSdtgXyJsvnHLH/3vhFJ6Z4MIu
PSeni+pQjDGV62Edang5OjGxJVBWVQ0AUP5/DMMdbd0iqyCdLKQzy+Nnj6hecNAh
zYSRalxYKQ7PTab2r/DZNadMsH/SSPeqgK4yhT/t+CfTTJtXCyKgyPhez5/PpNlR
oaaB90d2ejBWhHS0aeX3mDYqUNHjvRxgmdJHTecCePAgvbJfj30f5VgQeEMUWLGR
FkSCGu5VibzT583eInZ/NoqXrxVz6DLLEGb6ZiwumMtaPcBhP7xQxLE7GZxC/xB2
kKw6jx8MNY6SxImSScj46nuPUxa2EZMN1KyeA2kPylnuFF4y3O25ZOuvtpbewk/9
EKchaXMTIBY+ckfmUoAeYNKl7FsmLFAi9clbVx5arxQskjiLBhN5wq1H7fTLja7B
pPflCTmzdfArqBODfP/6feZ15JtL0DNn/D3IgDctS8mYN1TX1jGpkQXx7XAQt1zb
MZFSQDNIotL488jTd3F8PQy6RHW5johKVQOnoLw3lXbDcoOloEDuBhLBk68h3Ubr
BnTCNogt0W5wwkJjV3kU/aAaaHnAHp4PrNwMU5m2ItxIrzpTgTbHCBTu6o3D+GHJ
uy+aomenX+39nrDjnrvFnaJyEWUvSj6r0surbP7dShSAjcLzjcb+nQevcGb/eNpS
DIYjA1jofFChFi4Mv0lqgTq9skKJxvnRb/ObCcrObXjFTSQJIO9CP5XCMN5w9ihF
0L5dNC4aK7PE6N+J7tC8zho+U8I6PyiZ15m86ko12znmIfzTGJO9fUOmIKyUuJ87
60i7WNHKy/IGLxhG7O+Yn/rgkKQLBLVLSLnXowG5pIxydJlZoXWJqHvbx7rZr4rh
F2BR66575pT4X2Ksj7xlqQNbSYVCI+lJ42Yl+STU5A1LX8a1k3SjZRaOC/eWD4V+
EG09wt17fFYeEzOpiMdqHxm3GULVPsHYgLgoBz8Z2lqyKFAXx3U47SfG4kDO8vOA
UB+C1CleuNpHCmCIxDv+WrtUg/JaGHO8UT/Ej5GrcKQYYSYFkLO1bWMPZ/yRcjSG
oGDQCBOGg9XIg2NyhWIquUUJgQLUlJk6/ik3dRlCyrShZrjtn/4MIbcgICRVcFGr
3YsSfbXmssvQYO49X4V0T5jItI6kHrDl3vS57jksQDXUyw3sDredzcZ3nvoh+KK+
GQxpm/XGEYfElhTRqgcLORJhOQWUJPlGsxSDWAC9ZCGOlAxJr1ehtgMI8ZAsK9Gt
jeP9sBEEO0oRp6m5tXeDYRIYhG9kHdFWWwuIBDTOZjnxOs7RVZQ8BHCF8d+UUSuL
yqfuNTlvYsp40drsPNKQMT6X428viS7jCWHxOLcxQLsaIKd4L2t1DIx6R+c+FHTy
mS1Q5iH79wXSxmvWBfG73MuADKSt+bG4m3AZkBeQgcXT2sHTAcJH4f7H0ZTBnaz/
v8rjHBz79wgeKbArd8X8y+9JA7p+bDsVAmK6A2fj9P+C0sVinyiKUIaH+C/f00WY
cqPFJmOm9iMwiXfBsyrTivkB94SwjPorhYoDFGhp++psE1w4Pcgn6o7z+IkNhikM
Ma5o4LCT5C3Tx5jSgZxyhkt0cTfSjyu2d1ITIQVKb71nsjBWYr10fkVYGAisyyAT
pYwwHRYlBYalu1GNFZHsRzwScwMQbAQL4uj5kASBlQOjFyUhmOR6o1BlxWSRRhLb
33sqMqIXs/IT4qvbPK5e3StaI8Sjf9iU+LoaP6iCE4wKS3VZmJuwbmQ8tsE/GDVt
AI3ug53N+blMH2ZiJ3vkqrMdTsJZittXCkA6PlMEKnD2IElBsYesb7jq4Txe8cYY
fUtBLtf5og0AUtyTxsXZUKRPKIFOZqril457u6aJIboQX4px2IEeZS5/rIm4x3To
RzOCdbYMmoo+vUbs30GVihH3jyMnHqjW/Y1NRGe6d2n5xXefuqiowOoPeJ9Fe2IS
1GzhW+r3Ks1/u0Q41jWftM0Qm8N1AHiMMOlLvfMD7ol1gXjqo43WSfVWLgZn1DHe
zYf2zz9ywAlZr01bx4v6ib2qVRHt/Wxpe9k0nGQT8DHt4WC3q3IQvgZ+B94FK7qQ
6NLpp8Y+hEsxGCYVmjx2z4PaXEL46htToCQ7e8N3aiZpQ4cvpvabod2aGzFWTcLl
kX5k6+JtO2zT5QzYnGae6uaH+6IEV/9oA3p5F2s+3mZ737k2bfQKKfc/Q/iOfGi5
/I9FvNp4Ee7QxpPXi5h9VP+CWM1ISjOeMlL6+CdKpA6E9yusitKyHEqyGVZ/MQIV
EoOmkwFzh7dU1IvdkWqq1PKy6zO2CTieRmRS4qYBgDMDwPy4EGEhFaOzF/HRKG77
PDij+158pSUJKc0X/mHK/actPvzcdtcrg3PY9OKhnSQ7PEgOyyqvjgbNraaXqErm
3X6Yj0SbtoH1uR2wq0IITPfIgC59zfoz+UCUgZJPZys+wroiwRMIW9OVZOdRPS6x
sZEe16ub8Q5uwotURJx4J2rfPjSmweU+nC3UkP6HwvhdW6n8Z7dqMO77Ku+zRcJM
/qQQQSMXFiq0DUCbXLOc0NHgSNEQ0IqewrQYQbFaYEr09JC9YocEQQx9V5QNKsSv
VYsueu0BOCNn8ql5+M8i6LRBKWmiiRZGwLDHOnU75EQnmQI2fZ0uaLWCcZrFZH5K
Lp7MS1VVd/vo5A1P4yDHPt6Yo/ETdQcCez9vBlGyt7LIUxWovjh7yTiFJuwE8cPE
v9sspeqW22wSjS9ckorAT4TcwzvWVojBzN+ToWWecTEOZtiU7NGUSIKQ9PLsRGNE
AyfrlZEU1rryLTNoAAGp4nn3S5PLhKW2lajrJ5X/CxZCdKYRxgF8Qw2h7D3N0BFC
v1mcz84rJj0hsSZmpSNbRqmZwAknGQzMU8Jd8Fr87X5Y7E6IfvDdYTxDIWMo/Fmb
FdtI3x7ZndTCv9RkUl9BSqc51vS14peDce/OPdcEncviqLlwTdhE03YV0+GfexhR
LbPUy8RMWEqMrrVa+t2+3IQnTeUWpdgTfnTCwoNBkT5YNQPzAe6xwpw+hL/HZyNa
BcCRf0t7Ico3wcGUpNProbWZ0J6iHb61dW2toraEoW/D/Y1344iMc1Uo2Da/h9w5
YFE9TqFC7oFQm7L6fr6M44D5hsoG2/fWRGnJIV1hQyAar5r0zBy4MhZsFKFkIUlV
tpQvR2NRn4WwF8tXdeyBCh9s42h40feUU1uV/EmOle4BhZ5zA4KbVvf20Y0gS44K
A4pIlD76NbCibbzYxGtHVSGYCIRKZqqyikhowVUeh0x6G0PtpNeTsRbM012QwHXv
ZzyfoG6gbqWW1EvWm2PbCw1xCYNErw6DC+zK5gwSToVtsLFoNPjtNBErLgowGVW0
q6rqEw7NTPGiiDqZAySKBN6k+KIjbTxUQ2Q0vT2TRFVbKGwpCE01ScpY9rmI6vwu
r5MBBPklWbjmywaMnU+80bKQcScSYR04qvmdGzWq3REORyoYuMHTiTWddgEFIJ/b
9BjCj75/3R6VbJASAngwSdOMdZefhyhspQ+HGAzzKHaOiCuFKB17p1aK9wb2wtYP
wKMfAWZ0V9dZMksZuEXbGkhvq/AdMJq02MCMJ2l8vL6QeKv5JcTC2x5TMesF9jEt
RiRWeWQkRRyLgRU0gC91PDGhdTNu7U1FIIuJzAU9mJfCQNAcPMoQrMVlXCHkqKxR
J7XIezU+sdFPYam0JA1RAJXbKxJwQUyh2/4800NFMkYTMUa4V4DzDdXCHF/ZxHT1
yVgixqNVokDmpO9NNT52MOaRqPIcBN6UCWNF4ZC6D4I4PKHhPRKBHPmkV+00WKTn
knetqtlKX/orzGATvSAE77FeSxHs3GXfp8mK5P1jrH2AiX6ysV/VoEB0uylJUKeX
RXpYbW5C0ywbcS/Sy7QY1kTWJ+9ojyYQiA/9QrJv1QReS09G4mZqHSC2nnGl8dIZ
4Umun+xFv67W+MzGGKlGgrQKf1VyV4bhEH4DrnSZhaLX7uaBzYVbNCjzl7Yr1Hym
dt8ertwiQCPDLvhAwuO4Lg+u3gFWUWc/rwfcwYHN1gF4Xw0rMtpBuSFylsmtgX8Z
gq2mJnpUc2ASC/87Q8dmh2oLQiGIrs+DWwF2pzMCIJ2X1VS4lN7QUSr2D3/4ZS2u
8GatwLFygUdgr67FwNNne70QUASEZU7pkZ0QdEWdeGd/iyskicruXZhxhsHAW414
3RwzL66Pn0VW8FTvGr6VLBFHWnthIZIvi7OQkmh7hxvp6YvGN76GoPDd+fcy3JX8
vc9PG48GkDYE9N0bnQPbXQuKhiy8Zpz4yanGsFInbtAc9DojXsqPjuRfpbn1K/M2
NEvuFnOb6M40WrlJ/ZmxXKzzrj1un8G7xjoOPkqnD7jtlZVfNr5o2dT+LQkL/xsU
GI/9TDedWfH+05YVXDF4jfz2t3j8MKLX5MsbHhbAUvP9PJegs/mpmtxYvUiQ8b00
WWhw/r1YZG4sSKsepN/QdBTVQMfGw+A8U97oDD2JlbZbrPd+sKcGFz/KJVi+ojht
ThxG+7ZNo6Kp+EMUeUsKguMRaHyfymHM0BxT+U7eEkcIm96eKO6xXc54Vq8stwfG
2Yk1Q5O6Q/9X2GRJQlqYL4a+lzHAyUrz1zhzJ4zMAz+tD8VWvuArTKhUglkijVS1
aEjbpK9DZ0cBsGRQmgQiuXQdGnBITL5UJ9jXaTZEGhlWRvaPWW2EuV/uL9YbFcmh
cegX/67WhqMrFfENEOBC0buDHb+WttDbDxxc1F7B8lHswBnGYyMS+PfmKKJsBCTK
ZlWKIxxuV97K03iq+mu55BieCnPsYwXf0dCqQmif+Lr+hIKi7hjMZlD4RIM/iHnl
/TK2Rmt1J2KeQcyac2f0slgp40k3tFOxk9Ri36ORBn9JPozzcnPNoYyS8ZD5YxhF
1yillEziH4Asj7G8Sp65MbzGPl5HDeQuBCOAo90+/ksk5tjlB8oSCSETh6g2nsRh
yp+zeXzQxXIZ7jLQOvM+AEUl2zrEpf/I5EvDW3M/jSyzTXBCwjHQFyY8W+Qi7xi9
n3FETw2cVqHQNj9hsESObO12y+B/RZRQkPdKistGlMot17yv/HXqwUjzslTXWmuK
3+g9QaEcNUQVKE227hh1mgZeKbjhMipV1nLs3jqWtz0u/RI/fLmmirDrZIQzaTzM
F8jsUrDNSOEPUSMZBjNKY9/tj91gNI43Yxbvh5ajIyeXucmNqv8jpUfvZ4JPmfPp
yJgqEK+IFCDaEsZHWruZuvXJVl1rBAT6B1dcbsB3IYq/iD54Qs1GzNuV0/NAvQsC
jDnzsR0bxEfqCo3uP2Vt22B1os280O2zxYqsBh+NIoHD3qzpXZJXbBKWKjTslI8s
Ekm7KFjy7UxbBmDQFQJNr/WJv+ulFeq7qJyEvGSyWO+w0kDR6JMDkMPytGd1bOW0
CptoERebMJEQr9teaiap7WpjoqQnLPWSxPWfISymdwTIv+8ZslESbRFi1FtxoVxA
kWaUmYClTMR0vEZJflhfoyXpCDLnoBceY9MH7kKvu3jccZlLSpwyzSUeYmQs/yHm
tB7p5EtKpiP1bEhAmMzZGda/rVCeYz+eE9ktXNamyil3HD6vHe7QMVDagPu+h0iy
kt5e+mDK4hZDfPHA5Lrn6z9K+YuAvCLcnR6nduo1uaqjsiiuJYMZupVmtJvh8CSG
hIDLgOD8GdSlXw1Ht5e+zI+hkipXDR6Ehb04S7TnTMiM9dyUPdhPpBUzJF9fvi1h
sHLgmkSOThQCoKhvy6TbkilI/sH3RPrDzGzE7i0C7ylUoGn0HjGhE4yBVcWGXnAa
5u4vJ8CFlbor8r6WIg0KioChdmheF5ghoEU3+jGxsMP4zKeBSj9oU41P8Nzzqou8
fwuHNF2++EhE/4VsYTPpxif4jUSro9zw1dIbye52PgwZ0bEwYMTEOe+7mAqQGQK2
hPmGqtdS060DyLb7YM44KSngGj0Phc9rGXrLRh8r0NpK+hVkeptzUL50wbaAU0nU
aunCDhfzfOksJ0r1Nq60Nf1+vfZeNd++BXknygrup0HkoW4g1lKRU9splZGy49u0
P+SQJlMBdmQutJ9MUgWbmcUlq03n4YFjIiw6o8b4Zs7SCR5TaZCTt8cKEAP0mcnJ
5UgjM77vmlNQUB9aNXjS564EYKvSZZBTm4089dee3uvG6z/Jm0JfZM1gI8a40x3E
fVN1PjBq0yErOb2ZqNarygc25Vx+mVyZToOamzFUca2lLErX9nPWtUj4Qy/WWnqb
uyibMZuhOqWn/JA9VO/UJe9pfvSaKPX+22/Jj7Y6LV9blimcENwlrVUUQKE2OB59
VmHhkrB4duKfDi8fcEHptCAPRVWFVKURWRVMvhjIdh3w65PObiJnyIFTz3zPsTCw
33kQe0mx7dw2O0rResk18JrWextryTCul30HX/ToyGwLu/TwuqBkvCWbbYTfFmPa
bJmEtxr+ae8E/9Ns496N8XILWfM/ajuRXTbkVo34Vn4JucoNocQglcRcFixuPwKn
hapUv3kJ4QmZo+YVdHmtDIVUzslka9QzJq/rTIfjogkyMMC37hBnsa2CwcuCEjha
I7vxZqGy/v8lzIxkM9MoH9Jo4jE4Obobozw9JYp6/cDwuGQtB3Jbkfp013XUnkXH
beP+qH1qNf5Y3VbOHbOqLNnw/29kKfjN6/1LAP+s7xVaOtPQ6YCizryJENVIAmuX
plGvrvlP8iM3UGMUCX3edZThaVLnpJi933cP8Bl1+qpwh/JumoXM5uFIUC3Kxei1
FFx/e6Us0opTQ676fgcI1vIyNmELvaGU1XU7qIoppv+jfGGrMvJJ0XB7Dze8nW/j
8spTTu1Li5YailRxG6mfOFdKiWHER1OjEw3WVXcZl3cPFAAXuccwkZIEOa+MGMCJ
MRyY++MVAj4gYrP32GqYTDa/qWTZVIMVuJELVzo1+u4YGkN4ISkm1zv76AxvFy4S
gVXlEAisig2AALnPEYUlzzEhKWDmCOAP2N61IoHqgRTWjik/vIB3IDDu9eYevs/Y
HptZmyaUTfW1AqEeHYOFYZG/3D5lH5kISU9AJbhhmB/0lVRK8AurDjNa/5eVYjde
JfiGQ4rROxshoZHDgEadv4eM2PtZYLSnouJCAJ4xIKyqkMb+ppGROlfuJz1am6DO
oLnEnTU8GDMq5+cm5sb4FXm1xoS96etQzyP3Ws1sftwnVazsCVea8sBHQgokX2K9
4jhsIG+jhtzg4BOCK1YDAC3HfLVrqpINR98hs3FIbrVbGazm9uFHMHgPpFrSvIud
ClJ1wb+yQCsQ7kyksMZN27DD1ly9Z//gBnPCTrdiI/bwxHU44DUYDZzpq5199mhS
QzqhlRIMIeH9K/0/ShrxC+QntbGKyY9XyYYZ/HIKJAhaCRObkTNAJOYB/pU4a08q
lG0g2zAESSwlsw/RhbDdqCcnjxuQnl0mgOF43obPJFa4REwJKz1G7myncH/MWLPy
6JpQVZzoDQm9tOdLMo1qXUEjry38om9YRoCxty2QI0WhLPV42mwWcxPpdvsai+hE
imrf3kQhYbs80jPKQrwqoNfFyemShDWQ8THmLWaSgLEC7JD3jS/Uox5xOhCn6x0Q
/yogpNWyWDbxSsUOsRBXsCHkavIQNvt1sU6WlxzqPR4HrJ/pFDOb7uwwhp1R3ZqW
F/VCnIrkBNYkd4+b4lCpavuA4GBeGfB/UFotrop0ddzGR7RPcAiLMuX1OydpOyzZ
VD/LGwFFqBSrb/NRvRtOx7IOaal0B5NnKYyYzdwXS12GSYWPBuyw5Exz7hwDfmM4
D1EF9Wt8halhk4WYWNsxLDil+HSXvJ6/DZp5LSA4agkjgoCf1Wju+F/kfTgc73GT
L7lAEpBzx6vuRGeyqxbOIl1/bdC/5SslGd/UJGwQsmivPi6aQ0rGTVcjf83Qu91X
6R1ymdLEb35KxhCElHk7QGSX8yjHitEqvkOFS+t8U4ni8WOfnSrXE7x9bZJI5okc
SDhnFtsj38gwQoCSC+XiuaYn99uUPVqjPuf0e746o97sKTBIiO7ZkygIycBFvM4v
V1PqJPl8yG+Mb2L9lAEuHPG9zbHy+N3rY8FlLziXJnnxfQTb7r04aBxPJISKCevS
FbGrpZI0hgeplqrGDNVElGBdmB2YfBUPFHiet7ZyHnVdRQ1tkuE64P3y6S/e6bOF
YYey5XrD/tLPOxHlJtjiFZJ8ZHXGKSnCuYQt+dIglnKEQ+xuSKeY3nJ6crUcPnGx
mpF370K2KH7m+tcirAx2wMZSVVzT48UCD13Pvl4YzzBgq5sXYQtW4WyGyWXGcrCD
/WR+MElmLpQqkic3orOYH/FWCfsL0YLbM8vR/jJ9IxOh7ezVVBd/2ozI2V/Hg7CS
/S1u7YdesNDpa8JVnhwZeSmkI6KM5rPjFkF+wk8EoVRGwBXW3xl9Uhj1kQ5hODPz
pB4HtZiGSuO0Erku5RUb9TTAuBfJ3aaOW5bitYRlx+seezqOLm9rbh00cIYBK/En
ZPBzb+VU+Fk9hoGwmC40seBOiWbsDnw2h7g6CQedfJjrnoFNYzd5m2VPnrRljPck
b1w5z2SNbZlJ6mgJ6vOvlyqsAl8H5AsWbWbi/repSf9Vt7mH+1Xifq1aVpl/eF3Z
NRYFekX5sCOaIx1sh7EYdWsAlYcAtCzISeo+sDayMiznGjOhUyDRK7EjE+d3hBJZ
iO83/uKhzDX/qslREVBgC8C7UNG85dA2Q4WNEUAI+DkeOfSN6J2StlUU/3N76Exc
2LgAjo++d13VNrEK5B9qa3OEh3s0/x3qbko8bONXQqCixBrPCfv7ZQQc14F+h1iI
qC++o81zuzdy71tQb+3D+ZREENdPIXZvkUVqd1a4rB5DDUJkQ3wYPz78HgF4yD4J
nDGzL0BxaglcfZRaKtYXvnGiP7S4cFMYQIgh7DTjZXK1l5gR7/7As2NFi7zOz9/u
jEtVfwQ7A/4OI+Dm/xDKf6PTAtylPPRWvBqaUiO6+GtthvcujWyec2aYAHV7sRaY
S7IV1R/WTVcPK+5ICW00efPdk66HIFTrkN2FWz8XE+veDQNXHQsA+QkTaD26+KG6
eSAblZVQuGbKO8AqxgA+0nVz4XeLvKeBPOgq9wLM7fNaMyF1lMOyjF69WiNXa7+K
pByzwsZRtClhmbWNblzfoyqWRuF3H3uk81sqXmVhSneR3WDxz2WfJLBxrusD4Cey
G5vOuXAOtfe3ftKy7P5PSa9XwFNCmfrnvynG6ebsfqSj2iz6e49NMcQFOj1jjbdH
wUJkenv6x+b0aj8wqi6qH8he1uvTAng/t4IxOKCtaevfm1Uy3CdZwoMwTPxo1xM7
rumuoGPtTSy3nVgYYhJpGcor37k83BA7D+2Y7urtRYKptDP0kWEmdk+XhAKTyuyn
+pIWyiHvul/d8sQOKTniIvJdXunGEr46cgn9mtJXZ6bWa6SntXAxQNiZxRaz+4A+
t+hvM67KhUiA+PqPiBc+jqLI2Jgk6Hiy21sod/vavbF7p+kCvXbIDz4kQecHJJcH
mtvqRtwUxXaHUzOlESzSsGjpy1AmlB6LMz/81n6q64W4DkfHJt1HRLzCu5PfUKOz
9UcVrTYoyvTu/fQf8cVvnQBlnAOMsSgDS5jXkkKIfHbOAInp9lCS3Z5zhESJySZB
D6cgVwUDMHAH7uQY2gxOGjGBPM/ahiCHXMz7Wa3P8Z9WcYGyL6krSCgC0HZJNhdA
qrJgTAsZwEw+YwfpA6U8FS30byrQMKjJ7EykmxaYzvBDEYXVXUyIunolSgkkS7X/
MGRQt8hGlzr8BiS+V0TXjiTi9nt/+3JTyxVqlphpw3ZntWZ3ZE0ksSsP8R6bt6zs
ZJ3T7bsN9F9ZYT6uCiRGC15NeSzj+FcLcPNrsZm0CboffUJsOE7LkFkZ1sKnrk6T
SFuyVlB3KY8P6zp68NZPM7qenKnItFJ4JNiUks5PYz64wMgarkHF904sk5b+AD7j
1NAy3hM7YIfmrUp9iXM4PRTXZnpIFNpP+UvPdZMWAJ+l4Q03AuiQCb7DJEBtFVZp
SCAbZKcnwmjjF19OCeuZa1ZUgzuZh07FROlAVVHaZtTuPw1wvU774MKgiLCdfgST
nfjPQnlfitKOeFnMjHURS/tRM4M5j/SOa8rPvshVyq6MTG0wZUrIix/Sny7r6EUE
FNuqktXWHfZwbGzKW8rP+96twonjjvXfVln5/+7Cl3agPWBQa9Hw6Re/kXlZzcJq
MtFiSlxSl7Km56TPfuPpaBJXIOfUXdZx4GLZ3BS8Y1HVZNZC7AreOoA7nShsEgfk
fDxyJbU/XQ8HnCVg96PctK/FOkCfX1KQiDO5VruauTAuJdgkr16KlJUFYSQt2lRi
717XGaedeAgqPU8xq+S1kZwqmIYgmgBayjEBIoYySbecjtXbnUs94r8YanPpdJlZ
RYaRD4i8DCx6DpaAAPWV1SbqyavWLiV/TxzaIGL4dL+BciODsSi9NEXBVBpVWEcY
VNSb1tml9G0KpvrKqI7DF2/Os50S+11Gt3KANI+LdnopXTtxHLIgJCiq7uppfh4I
az/CND1ekPiLtjZGv+HwctU6wtHWY29tKkoW0MzRJ+hSxPM1FFnDPfV9DzOQ2MrQ
LJve7mL//2qcYvdZn2trM9XZMnamKliZkvXVWeLlJzrXUER0lUEqEZAvMUCMxqvj
3MPFEsiBIFcWvoOp2HzxoDmRmbQmX5DAvTly8eRja7CIKZi4Pc9KBogKHPFHPcPq
EC1Yg5zMHMGNKC4u8NRJlIUFdRPQNvrorDLcOJVpRe61zfHJtC7wdBnuXcB1KH4u
+6RHRuicWS+WCptme2OUMjqqcksId8paf0sj89fw9kHnWjS5bKV+6lEc0gGJNHx5
GZpaYwlvslIV7q5ZLJBjM++IFL62h4wbppMT8XW5kUFglT/vGYt9KSFxi6T30oMt
wFshhF6UCe5H0zvhOgsOGkRKrd38na2jilHhjh54AREhtFfTe8d2ldpCLCUYXX31
FLLxswgOart/ggEH7OM4C7Co3FgilV6VCJcVnfYN2FVlGb5nD8sz1Q4SCcqjVqcW
pehrgWI6+xiecylG/rx7GRZ/BlqcsC+8Y1oI0eXhSTq+dBcOU+ANX7pvMTQUelB8
voXF072YK4UkFPeORA3IRj1ijag9eYrGZyO0fq2qahGnhiBU4Tyks3qboxd3SWfp
YnApwSYYmF+1bBWjAy8kS2adGw/3gPzPRL693sjfNfzUdfHTq62txlymdJNisAtc
olMDVP40wSzAbsx8gIXZB6PV21NwgS1+ceYEU3kRMFwTmOqwC9EJCWJWFb1MSfu5
MKznNzo/PGOOCEbmkZ6CSDNM/qOFITIrn9b/bRuXWBSSMF5vJheAmQSirg0B+T5f
UtL7IGWRGipK3o01n09XiJgewjCpeEZQCsMqXiAJNYV9K4S7cyHXOhU/SOn7u3G6
6irH4NZPX14XebnnjfmzPOiQdJanquayNxqfXm8o2NoFwBUFmnVpzUtiBdaNdMTq
ehRrTWiCY9+iJ6oDIfrMbzPWFbaEVGJ8zEVuy8/c4FvIa6Wx3CELOFEJmdJJi01R
fZ+ypd6JRxt+Ii5Ohhuuq5FAlWWXeEvmuA8QuQqox6q6Ve4l1aqwhJ8EFRIYI9XH
D7HfMWan+Tcg5dCOwqHUjkN4m6rzNMdLjy/wQ11KxAti8HHJiTjU/RFTVKAzKRA5
ApVEpX1KtxJ5zgE0pgAyOYFLlddV86+C/Q9Jd/WNYq1BN5b5xpjuxtZMH20tzdM8
qnWh2Qym9FtpHsx++YbNfgdg7IxSTjKD/NZGPbgUms+m3pSUUZmg8KixfMAdHaWD
zWz/pFuwHMRcsfYl0Mr9h5xK7/REfJXaea18c+q/iCswEwDRKtkid2vcmPHlT9im
UgrV47qKWoA307Ki+enqFdiPTVhEBsMPGYANEREs18lDdTUpWZ89AuLJEMwsn4G+
2Rlwwo/em6WU0wntf6V+Ge6yKZr4YnisTrr8c2EIjks7TGMqoia/Fu359YT0r5sQ
8/JH/Q1OqSVPdx5iN21kgl/z7kNxeoTnMdywMhvFaLXLD6Ps9FKMxBzr+tspGVBz
PCLFgl06fYXhSYlRFwQJ/5YOyidl27/U9nOkSEolHP0MjIdvb86WyxLbj0RJVx4o
Lk6ynLpujOgBkZeVR1Ezac0AJ2juaazfAdlan8P9kk7N0aHnKdUnCbrrkYC1IEob
w1Jb2c+PzH8rJE/dbbDSa4hHDycj7PjFU6ETQJYsuSos5IflQ/TQcejAA6L88WrB
bI1rrKshRy5dxpIMV97WUkPAPKJN+Hqt2LebJpZ4LiHpOFJoBLxtVmW8fdgyxUNW
xQA2L9abMFuiZxsTNa4Cm3YJizfyGGHKUfHIeBzXCxrC2OnGGVBRcrWOeOcywTPU
cQuZf1ftq4S7AWTF5F0IuTAMXL7+k4YloWufkZvZKkSlB1wcxb5sLWL9/MFQX52F
UeW+GeymWz7T5ka0AajOykOTr+lUk8XlWB3pCrs/KzqRmWqkG/EOBOqdI6X93kir
qYDOS/qC775izk1xCLuh0qKGUyDL4EDHZFKT3wwzvKqE5SQXE88EhOjpEuuR6DeA
opyMGsBc+d6JUbDae/CfRbyJfOrQ+0ljigQewI6cXYg4quvaKaD1UBB8eak+bETX
OFMZIXWzUBUyT37eOcZrHYuRz0AIQJk127A+ii/dm5Sj8NktTq4BXpjMoRyWtcbP
LPQZs1y0OqrbmKS10Xh5paz5A6pCwykpXGcWa3+ES0hxjNfSxt5FYjjoG7K4e2z3
ElEeCY3OdP06KTVJeGyLHz+1+hcyQvddWPly8E2cqE+kUGCYn6jnrzNA+ZntAI7D
0kFeWLn6xwuMec6zsnN6AZFtmFHUiazE8SZ61+zR5x4JSAqxt5b6xEE0nlRuxXhO
JJ1MSjSyOdtb2i26gAQiuGG0dDqhZEDvFHPY0GacdyUAfLRHKiCIg99gc9UuZGzW
T5XcPlodNM3rrygrhqWqAU1sDh82Oe5iNKBOGVLAs5srs4bJKKtZQEmUJKLELda3
dwz3Cztrq1allqshriiexNLTEOtogQH5AuXzk4/nPX4f85ILR06v+n/IOf5lDjmJ
3jWy/KDctTktOruzBBBA4dtb/Nmpk4P77e/h/CZ/Yv8I0FggeOod9wRTnKE9MhiY
am9QMOPTPVJ5v6dSboxXZXg7owGYLhAtvO6+ASrbFvPSiEL/Cwt9zKIkib4bGgmm
5xHzprQzeQXOyH6WKUv4RAOkw69EjJMNrHV0+mZHldrG/fNO1k6U2kjAcJbuyzQx
+ZytTy4xFvs3NFyOZAgMxUbq6cbTJx5hwU2VffxaPFh6HhSK/oQAmwVNmVJl7+OD
ZpVZ5HEK29Mp7JFmGZLRFusQUgxiVDdrQL3Ov0qO+xUQWq6WZr8ea7Vv3877QgC8
22PWeQLwvSrUIrUKW9VOXhU+Q53QwcgRCsDek8tun3SU8Wp0tGDGYkn22DNGilW8
kyLnACKwR/wtNa9hER4Og+Awj6RaMglm/2zhd2+37Ku/rosq/rmhvUfqf+J7NMge
r9rs9swv/Njlj8CSkpdYxk84jPnKNK7Nq6Z+HyNgq1UPfadux6DWczM5zK1GRPKC
PqaBOgzMylfpzs2fK7y6npe0tHk1UeOEloodb31qNXuCq21Q6ibSmZ/L/JHw5l7s
tagqagh4KoUv1U0tcsTkGMBJR/0Lzr7dIi0/BLcbpkaWKKcf0CyO3GwAJBPtJhL/
ibckWuAmQFZcRecWQCQwAYgg/qgoHzz2NAb4KYzWqYyw6HnspRC5h7LxIL/v4de5
KSiZDBctsjYsJP043ZchiFqryvwkqHaxzWTfXK05Y5tqnShIZLevCb3K+mRed+yx
tC5LRBDwam60aVOc+UFnP9o5s3YFKPSzOFbrr1GrYsloPEpF0wzldVw3pET5vMKF
VMwjb5UgZIlP6VMEFhCQ2mayBhmLUgQrORbwjIxU+cUc8OjkcNOZNsU2v/a0WZLa
TnLDQzAOWypztfInApxjt5wuYmR2fb807V9E/FHWJ1rWLSfwSxfCjzsq81I0JIt/
SV2FmCodgewpleFjjmJ4voV8ltxh1VOGPO4V942XP0ew8aVbasgWh+QU/Vdn6STb
0DZ3PKnc/qrH8RSZil3X+Dh83Lf26me3Zck8V8eLbmqn0BXgu1fpRCIM76sPRYLv
RZxSFa8KcvH7/tz6PtRR8vK5araPZLsF/MA8FgtaULTMALZ9fvbnAKgPgoDdjAsZ
yJ5OYwg4MewZ27677T8Lzp+AGNk99xTuM3EHcMl65179uDPtFVQRyw4ljvFK626q
NSzIEFHSLwV9WAelnsUgh0wGw48aX8VpOmsu/lSJA+94n556GpQmyu5xlRNx9BWR
3oamKnqDOYgtynCSt1cpgAUh80t9qFSm+oK3x0n//Vi98IWFZyzNXfJla1aP4t+F
HH4LmjlWmHSsXaPJqmefmrr7Xiuvj8vOLbYRwmGhQtCAlRJFqvFJmEMshYpLsg2e
66VIiiJCcjPzXCQkyx6E78LIAaknC2V34TiT9/jS4l2dKg1MQ3jIZTj109FX3CRa
9g1IWp4DqFxd4t1ZDzAj0EXVrYe9o0F2rm292iixDLL95OxVccQ1AUErYyO7FEAi
taUToilpXW1IDy6b0a1yCRCp3BVJTHKf+twJxbw7pIBT4CgOh0RjBQuocy8raFRG
nyo71Qa9Lfs9+38W+T45Jgtq5eWmfDlp5AG+Y1ePQNR8+dkUEN4zaCfyJcrUJxAM
eXaQ83L7/diZKRL6Qy62O8Ps/cvlvdxiPJmzR3jVUdVd/74/ind+B2E2RgunFx4Q
T70Ri0BD979K1caxJnXXEu1710hFodEVBPDlFyTNrjEtjc8//t2kfUdjnF/K3UMi
WyFXXJZPs4Mm0V0KVRJcAIeIUq/LHMOkz7qCArGhtwkC9hlVg1Fndm0vyVWSCLnP
+l5pTGuEhThZxdF1/gMvSgtZ1E6nr6Xg63BKEtvF2YeoYJXCDYKPPbjPA5q8t+F9
OKZ3+St0WFdR+Cwsp+DESox4G93/qL7RcAbr65GtiAjdei4D3EsPRaVS+/uNS1ib
BaWPuYQkj7OPtEL6++aRWdevLaz2EhWgUZzdJWboRvZl20WUoGNMZWjZEhCmdk0w
yiZdpwKt0e6hpEY44ndSxrGiOr9bhG83+jQ57zbqT6vJTWxVnfx+iqvw27bkXXoz
/DxAUWTnkBjUid6Hoz9HQ4VXs16y0uwlj8/v3Cy6m5It71+IhJ3fV/O3fluLB2nK
TU5xoZsYGuHLUD7WpiBbCpMQGYlpHwPKRnKTVOWMXJlULs0zcDlJDAeHE85et0I5
frcFoU6lp+31YgCl2Ma23TkvVCjPy34HEd7Iruf4sAfcd/YZpTP16NgvZtjFCImS
eLqoXzbr8W4dh0mWk8qR+URrvD5yP1JF3+/nwszmmL63Ju9tz4Y/uGn+dKlsam0d
q5qrmN6oYqKhUZisS+P2xsFnyoDhFI5q62b2eo2EcD8Hil7lP8si6ALUkeNpHmIk
uIU8MWTRZv0ATKQavhXLgLRhIUp17hQFhASlzSLSqH9zOgFHDIiEWL+Vr9mOzuv0
wSg8t8JFWXgu/qOJbQhDqiHnRRioxL+jEegMfCR/r1nUUKephqdR8gOK49EH8m+7
0Wk6T+XEK+aIxq+pHQj5aFwH/n+ji6yalN0XsFFMHKmIly+Ypr544+2VFaE/Pfey
cHFL4Uw1jW3ToP6hV1ns8qMH4O1oOhGfJ8moW2Hmy5mmyPxhH1cAPJU633Tmxhs9
6GHK8+H4VmHbc8KGaUJcdQixjVdwbQqzMlhttZomsXroVjyza5DQV81kxn2yBhX/
ouqHzRMrE3yZ31J3/h2Ax5I8Od+/mCTjJ/xtuSXsGpabWePwSlzbXyXge84n958U
M/iwg3oAuHVWtEW/ML/a9e6jqgjDbXke4vsJLFq6nYDVUYQ3BjWx/f7FAVKyh3VM
rZaoHBXBE9JR8w7J25lG86HZ6KO2Py7xoAwQg+uKD2M46dlpPImRWXEACgbi1cXa
gbD1Y+Io2UGcB2Dmx+KOguO4ndNLJzPrRtdZTlbQvH3hCVQSBqeWy36refgEIDKF
q3U1NHGg13jrzK3WnNfVRSFs3HqKhlEsVgw9rYzdACx1mjfhtKdA+JtmPbvqe6so
1fwkqR1eeofiQDUInUNA6CWgfLMBA8q9foo7plr4DpTA7v8Li5Xto+x73vkz92C6
VxSVv55eSALwh2cSmpcSxx48aSUCTBkeC0tvyXkDL/0CvJbn5hN4JSWABITidpXY
PKwy5c8mBETg+xp4DtWJN9hDV/2j2T3kLyHMobpLOj5yrVwW6I5qQFolYsr+/5PQ
qqDBPHwVxghU3uEPM0ws2UOuJDyFjXScyP/pbY60I3r9nh8ABEVbxTuUb9RIDADw
fkXmtcGIMorzVur8v9A9CKbmN3TrZvae4zOlUVYItHiXAJ0uveInyl9Pn0c2hk/m
3OiCmihkmH+RMkDTgV3F6YbO84CL15wo36sTNaZ4E+IEKAE1H8f5hOY5Y0N6f9yt
q1KS+MzJt/G4VS3QMRAdFAlA0qls7tLKvSg8++pcKNNSN8+yxjnzlGxIlcfUs1iW
JcV5Q7EeAVnUPinW3j/Ni6OWXcdxh40RWmz36b3raEN7q0P9ctZU+bKiaC43odvy
Ig+DdLW5lZeiAAsd25TMVNMpH/9w1hwxDVxW41yccJAb4yA7r+MZTErf1g4p3IJa
2ZLlg0y+wE65b2AvD0hHe6ocUzOxZ+fFPGgXJ8H0yYjHdNGy0O1fM5LwhCJW1Cvn
K6DzLSlGl+Ucsgmrn9djTskP7/g2oHAiwPMwqs/CnueGqOJtmAJSyTdsw08QWZtD
2PicNdZWHgFPWObY5OqvMUYdhDoHlykpRezeLEzJgthsfecEFla1+YpIiZQlb9ft
i7skSO58WatkV9JXVEhGdcRcw4y4VwH02bkbEY+YC/iEmZ7kSvAnXlVvvhYKcGzR
IJi4W2q4cGdSld7e7lUo1/rdwu0WSfe9x0m5+9/4r9dcm8PwpXOgktdImcGbSrfv
RwkRL1NlSbnDJqOsGeio8D7KOj/cho/dim9TYf8veubOXPWFeiWQYtIqeSs1sAwl
cE7cuau3JtxMxeUIBpMWUYigtBu3WJqzWzmeVxEhw3FkmSeWcycqUhd3VOQ1U7mq
asudKBI18jLJdL4Mh120ahtLAoFZD1DQmGT/mEknfBg/by6R9SKAS0cTnD0Lkigq
nNFodDao7AASD9VRoUQiqRTug1X94AZNZNGYTiyXCTAoMfjnA6qW6kATYNcr653M
voqa3yesKNNwjJDmOAnK7lWE8l8QQ9pcZD56G4sLf6zilC3BIT0/T7HHuafijamv
lIhRt0BLe0mfyuH4NKOH2v4XNMhtNlC+nm7F+mgjhP0mc17LJQbS8pmUuc/1C3+k
q45uxBd+lfniO2U/LoRcQ0WfMvkqMQa3xMSUqkIYR4Jp/MxByHWPhr2awNB6IFag
pOUIWpE1mj58IfJIC0iHtAAPhbPI0nx5sHLxsFD56aKULonhG+Wh8I5CCYPaT7pM
DXcLBK6iqEvs/fQPxBM0yVjnBqE7Jut6nlG7iPcD6CgvcXbqdaN9Hef208YqmOub
vh9df6L1ePBya92VkS+Mc6E0vGzUEnedIbSuMwYAJscLWEB9Qd6NUx5Mrm525C1F
GvYt+F8m+05zVilY0agiHwyheJnJQt6bwhzoRRDLErpPP8UDyq/vGG1zXqzYaA80
sC3G5iN8avcsTZ8C0zTOoT72cC+NE1u1/paAQenZQuWuGwIUubhoxpBmDXv40N4e
5khIj6HVuMcLUj+FIjZSvDvkVpyNYP0YkH3H4f7X+MVfQ//MTe7ofV+5104MjKBS
wziHUZT2dyqTKINuH/L0m77jHepN/to4kmYK2ut7Uq8FUWu8ufaQ8zMnFke+TKvO
ZcwVpy/zE0o8c4p+/QHRfp2TMQEejLmQVm5j+49oaO+D9HMashYPlRKNUfIHnj2z
HsMDLw8s7kUwaI/l9Aci+I8lC81jZpNMbObwWuI0OYm6OlY28J/bY0EX356WmQiP
2rts1z6wlEb82X7HTOVl/INsQJzWtWb9bNEi8UxRJ6bOKUMyu28F6py5VYmx2hY8
pj8gcMMvtP+YENAKjxLlXGViOTonma4IerZrXYTwR81VjK+70bFGAGGBkEcm+F6F
QLsFpsdqWv46ENI9akU6h6tDAYJQnH2bh6rGmJQ5ki/BEIQczUB5ry4oAp1JOcql
H5RHsgv3PkfkLd5kyOfsbwkWrKYyNGBECmVju/teVMCKyZ1pp8nAfnJupOI7Phrq
Otnwn0LZuhLQxmoInrwOZ2iZAgSiKGXA+C7AYUTvGeXRv/pqjlPNietk4yAMfVj8
vftvUFTk9xBk8ZMhxGwSux5bmQ08bHY6L619sQzSA+kg9J9i0Ize6cJULB6RMwXV
/hWUS5dgyn9ee/hNM+N6vwKqgmBWRchtfEm6O/yFgB1a14j1mZsc7lzGhCaX891d
2SunI/H+N7s0Rv0rmj1frd6IewDjAwYjDEF6YybbPp3SQ7kiBkeVyQcvgjo5LsbI
3hvtQquum+EdzBB2ya4zOODgcTUl9b9CsoegJdFz6tqqJx2djeT8kgq+TDXTPSp5
JGoFfg61W9imosrIoXze5eB7mer6BSXLUmh4RMepltgTS3DBxb9QXJqMmSMJ2Ev1
YftfOIDONhDQiy/0nJmEOqS6uxIpcZGJhnN7w4Rd/E67gF34krO/vSHBIsjkT5Fh
2WjnzwL2yLzwAV3X/EYGX5yXf1sGDsBjShY+bvklVrolsT4t5k5IKCpEQYWO4oWR
HEiuyZjHwFa4U42d43tafFBW6RhbhgTXf+HCMB/r4scov8hugQjZmEDEXzCKGaYW
DlB/iTAINomYwMFWVSOTYLi+UL1g1zYexYXnsWa5vyAfLJ/aoDfSkadSrM7SHtah
sYYqq3R9az93ErY1OwGh8g1KcuVlM28vVNY/Hl9GQPW9Km252i14NoPfwcM9/Dvp
oWCk5+lnEqV2I+PN85T64/bT99iAG+sc+0IxxSW1IXmDa8stTgvh+c5wNa87r/pI
ibdBGxcygCkIEQoBEeC27NQIdIIFru3s3m7l+P8VkPwTArp45NPQvdvhg+t4Lt2E
2L7b6+7VNMd+kjA7+DxDFNLvoEap9EKYFqRxq3nq2h3dCKGJ3vWxUm5RfeKnjxvZ
nWPpsPabQcM2y2tckc/XA+yZ9M7iJGBq3iISQnKKXhF3t9KgSRyUp4hI9w8fE99L
S6LOiYwHjXpmkRLPGZEqjnPHGP4Hp+qes5gMADeT7xhrr1OAUKj7Qbc8jKt6d6qw
qVevF3jN/IOmr6JL4SvUpCjj1qlRQQtSauWneC14qhu3x+kzKFTLMfpaeWk610l8
5zItEwQvy6N/Rk9PhwocYMol9JavAArk6yHgP9HlfzgCtN3nSDV48ANKbvUHYjPH
lTo9lvqes/V+DlzqjV2S3n+vZWgysTOas+yCWeSyesOSYt2Ub7mjCqcEPM90Rm62
5o1nxyl0UhTv8DwtycJ2d6r6cUZ5MV3gUh9fL3m6rUaj/qoW09EI+pS7OvF/EK1k
F58CzLkcozfkYT7Mm9hg0S49sse3WYkxoZ+lRZCryofqMaa03E340/dJaDoj/WnD
K5uJE/SOQuIlct0noQbjo0UoY9sGYIiN3IJnFi2icFJlq3KPjkF3ohhPKxRT7B5R
rNo0cGhuksig5k+EqtnoAqWFyz9N822XRlSmUygtHj6jwtT/go2vxGEst/A9BQqy
9yzq7XjbxgDLpyFqrqtkLcNvcff4DnWS/47zXOQfKgicg6po8Witd55PDsS5K6rv
EAm8+DN9PwSuX+jpK3DyTod9IEE3+WGjJ2Eeeu78XFB+OPFj1lCGPKaCg+wOngtK
lI6uP61K9VeiX1OgbB/clWwxVyxka9IC6TVTcs1K/0mZbYM6RIhzZhMZNEo5Bm+u
QI8alRg3acHQOK7d6pH6nX/+3S07aEwny/Eq1liD7YPOeafo9jxjYtLyoJZM3FRb
Fr4jwE6p1j9tbSLtyuSYU+1LrLwrkokfE9zG2Ups9qhqnq3rOlyiK7ZVnCe3+Yh/
GR5YGraIUEGhn7IjctIKfixhxvwM2T5KAKnMY6WvBHxc8HJY//6KzQOAASDyl/nL
G33yZm8UNDWd4kc296Z6Cef1Jd6NMfghPEDnmGMwA9qzumxpQaGIHZuIIec3D6+i
kso0QFnwvO0e6Jkrsok8bczSAzwKm6/Z0dVgyCDP7gMphscU/W4KlD+DT2CnVWmf
Q/jY/j2AgxxvEQJqQWRVjDVfYV5tb/Cr/Di4FRJv9Kyq6CVSJl10cxstuKNyreY5
WdExpDLVRyU68PXRskeIjr1HVmVbo/lOSpqnb9gksltznfYzbo+D8BqVHJtPJhA1
Z0kBFhDMK/CVJjDfS0jVKfAe5bWuynO7qVhwAsuvaRrmAGEB/xx4XKKfdWlfpGB8
vNZSdSEt8evJ7AS+nV3K6APog63o6QyW1lJ8O8R0s1Nys4PY8mjD62e0tRFFV20E
Iayle7322ApKLPLYvLnezoVgVmBAAR2i6mw4eGkZo/P99VcvgJvezy2Cay8Yvy26
05kaTJCspMXQmwN4WHbmclCBYxqk2sr8dKwZ96a9Ih+Ljgvy0v+A+bIAgHB/a/1j
BIcQ4Dae6jIV6XvPMw27DFZlhJl0CaHmZXovwQhpiaCCoLcX775dsKTHBavV2Zos
6gF0WVeQ0We4So19inBKXXmVT792Wre8zso7lV+4x8fW5TF5ItN1GT7GrnEJS4Xq
lOH28e2Aoq3fW9EHVLDUIB0RUXn7z9e33v2LkrkB3ZrB5J8KyjhDliZPd7f0pKlO
+/xYmfEKIAQypShPn6HiOPS65xZRPneRFHVyjYw4p8oUpnIyb4n8dmdHXCeLuYRy
3if5dgJ09U/Ho0IBgLBabnLXT6SIpb1hQD0RwJO5Mm/Q8UeBGhyLOfOEWlhPa9Qu
D9b6NwvsTikRoVP33j22nGPQ1weuX+SRqV/+rJUBRbnoRUq39mPngDqP1cZ/nr4T
bMFAMFNvzr5ct14Xvt4xFMnlG/enIPNU6UiuFc8D3ZiR3CirEyJsfF8uj2o5Brce
pAWyMMXrT3GFusK6SWwJUs05dJGz347Ep/2b8uG/cS0KiZtoxvF78islImjVchLf
nehqo9QzDLkOO3AdBee9E0jjCt0PB6cO0p5wyt4zE07d/oqArkvCptIh806eMy+8
RAmSHjVvBwNjcEGOvL+p0t0XQ5+G8SWqaHi2y3JvGcZazQZ3u64j3SK8fTi5gHGx
L1dqndgCzgGex4wm/JR1O/RAcbM+4OHwTYiRwaBantn3rP35bs8tK3l5X5AOUb+P
kKQhevcWKTY93dMuaidJ5GdnO8JVM/FOC41+6ig9GgJewHHwgt3LZGucAu+46Gw3
4N5PRwzoDhO9MDVBe6appMi0Dqb1wDL41Xfi+3Q6Uorh6qsYsqNQ4aMsnhzSdlXX
VwilUR/gawrvCfRCcBobFYuTiRtavfRk0QSMKdskM+hHlsbLP3YoPQwly5tq4838
LnPPVBFrvHAji6WyphxhJPsBuvP82N9BzmdN2dFsAlI4Fbf3MjpOyBoSD2yMQJkz
cWrgvuF79GJ/wDNRQQXaC2elmJ8kwoerdiW0/nAwbz+Ys9G1EEvBspmobhP+DY/Q
MVPD1WsBoxwp/AyWg5nQ64jfJy+5ij0ZUkG3LC6JH7NHZbd9TkUcz00nB5vvWDZd
+YbbROHUPyprVRSyifZzgAJgqLBCptTGpauqpZ26E3q6jUt9/p0+T1/xozpUdclw
d+ZxMDhP+uPfs5nx47q4PvL+FTC02pzEAHRgKESMbc4XlmWlhxqSEu+v62cUfUrg
LCg/EK56uCDtIQoSPTB1YKiozcRa52KF74GpkPa6VKw6YrTukDec8ATYAyDjRlOf
VQ98lq7s0wS7nPu3VoLVyPWgvhCamvM3dbQqQYCE7gvghM0lXATUcnErAtmG3Bu0
DeghC/EodMeLtfOMbS7E5uacLqxGK6yiVXRY8RwU9hwbH8R6EDj545kt1TDlfj2W
XoEYSmVfycpJ9oRWnHPxf9baE+FnzsoIu5b5sqfSrssw2pSWtk6YhmY3D7aU7hNm
ZzQDlFjZBrTicq087QtH6aGSuqMt0BTOyABN8dBvkCTRHMOS+Tt400Sctq2P8Kmq
wCHyFJruwsNz/O26zBK4UxS0bZ2Jqn0uMzQdoSom6YQSNbMYqPuVNgr+xunqyJHy
daSa/alDCh7Rq4m5oKNHPiDhCYb0hUHW4MA8ViQ7JpE9RX7sqxRalPWJf6r9lebu
r+8VpWxXtZX04JgmxYUNqgb8j3d1SFpmk31+rE9+Rv46QAmYm0KxQJkJytM5+9Ve
ya7yWpCn6IOudhtKfhag6z7mWszfel8baMdYnXRZuJd+aq426FFx7Jl80aLJoNlr
0ZOyeF3VTQ1leHJC4NswC0KDbpNcs7HX31NLAJPFIfjBpKP/KtAoaINkVAHScnMg
iEDAWm8gy/bb/EEr+ViT9pJ7EPxW+K+akuaZaldYxp9qZVBnQvV+e9NwVt3WUA1B
0BRIlhtyuuygUSdwEocsdM06VrrN6UQnItsDimKBeb1/kgS7rwwrmGjKEpXV6Bxn
95heFFViAwLguhGkn6wFuYqJLxbDI48i/DBKWBr2auOuRixWojqgHwFz7CYvy8gp
ShsP5ZPw8wLskGoo6yA6zboP3/JBA0hznZi8D4omduwYZaDu571DOMERthN0aIp2
2gQCZAOkW7PcxYAlc1+VKae3/6M/RLBsdvL8acLlfOTrDwk6nm93FrAdzpv47Lbm
q7CDFyEzSHxDznWIg8AoRSaY2ZY9LL6KweOww+zV7eXhe8C0PFMYUbmbibByjXx6
s3aUAfSopHJWpnfQGKorAK4BBtewSD3j0c5FLoto+uZwNa1JS49KBrH2jvLDsUiV
4HmvdKtqFaFP19YzivBc5r5i/aSjGzJ7/m6ArLEjXiI9gtEAQ5pVzj7TJVJBG17t
fU6jyLOyGDbgjWAm7U/e743qqwFjAPCUDRHLmPL1iGB/+YeMUJgTaZ29vLiFChYc
sE0lmGzjrBo/flUsmw3ZI8FRASA4XhPmDHeoJtHUqIQfe75n6oMAJHvQzm6UOnR9
o9o6ZrFkUKP++mHKsQAHoCnAFoZKXOJ9QH3P0gLkLWYINT/tH61gTqpmyOl6qj3T
Gt5E5zH4adb049/SXNsvaBB2vXzmW8oHO8toK6/okhSNUoX4Npidk+HYT4YIRDLa
jBaQv2cTYSJSnFJwi7cTpdC+C3HbQhSPyyNEDHXUIxDrr9lVEfjR7hx4WCN0uED8
BsnCc8B6wpjbbkQhyMb0xhG+JUneQGHMCI4bgbR5mYTMX8OVWsHGWSXRySzQ3y8O
Rue+e+tVa2q9Zed7VfMyJxyOW5GKB68o4OYkU6NKcuzBjzS2hiY2duDk0HFlAWho
n7x4fwUkt2o2/RNtDllVgq60ldflHpAzButA2u/Lq0wmVBmKlZU8JwzIiPClVrnH
Y5DNOrVPBZ1DFuow3Ka4G9bDOyPlRJZrufMldDDUuRBH10h6Ni/ULEBfHZfG24Lh
FuOvdJTuzYqCZWPHXFNWkYuqGAQhYNeuYsZpYwnSpxfqqmBTgbk6bS+XVZ3hWOs+
ZGCjMrMu9/reAk0thsOjQbkmw4Gt45YvlnET1xeXjHHh6UgAt9G0Cva4RL86rer/
SN7CQCQFhXtCe4YgPJVoKjJJhagnY+UUUDRljOBlsoASc9SUIS1+cKOLYR82Oq6A
aDDOjYx7SsbFjgHC3aRwvU7nwbt325e+A3ZOSurYZH+SxZ5XU5X/c4GMEcfu+JBH
HW5ZVdFHWpMms4pFgu+haPFhLY5lmnCwSHJsAGPFJD1A7WND4FrBAV54CsA6eMvg
M3OAm0qC1LXSXbcjfZ/yY2yMY0QognRCx+6ZDGUmHrGNtfqyFEnOGIy3KyFvZUef
OSvsrSrov6tUhlocamv2fgbxHG5z31wMuNcTOL+wUpcS9tczfdXeTbxTSkGoZqV4
y0VrAB2O07wMUuNFGV5H59+9b0zCpAZ5+oE+vP8r2QxeWR9Nm1CD+ZH7TCIANQS9
YShKEaJNx7tj/2GrbQhhziP8xnBnFVWFCMpO6MZhIDvpTBxm3X8W50//JoGbARhX
wblRw9ymZ1ltfibR3zrXuOsQGeDNqHD0WlKeYKqOz4DOTKn50PyBJxtbHaDB1v4E
R0QC97hgh1BsR/ScKE24QuuWkjypSyFfrSmWMEe4hAxDye9Y+TssRfpnSH1zfdQw
qNnHHThmjpRlKaLFpWF2er8rSCZ2q3FW4I4AT8Slotb4quD/tP5SrbzWIN/Qay+R
jNdTvo+32ad0K//cyOVs7YNHTuo92BYgxnX5OQwYuhOzDV7US6MK8dVifijTDKTj
Z5mxJTrOWaNMLMN0Uxl8dqdR7fAph/OLgtspxGLIkHPR5NdochTO/plZNN2I458D
b/IewfOcyLzHH2nfTvoscXErzyBnpIvB3/Ajc3JNWbGhSAgox2c+Y0SpBy2mw8Fr
1aMtYNSxpfA3tJvHVmyTkSmt/sH2bg1S4KKTdNReCobRzrK2wUo/W15HO3tBDsZb
YTIH8lXoqJb9dGyeDbE1Rq1eQASqAIjqSLIWhusGl1xrhUnXTwpMIO8rCn7oaVvV
LINftd60zKeW5mP8ZHKP38EBee8hClHJ78AijLkqZu8WaVkxwT2oxTH9UvQn2Fqy
nyDsxi+HxXI2gNYiMPMDpjlwiZE7F39UKwFx/D0+aKO5vOR2L9DouCxkEYB/L45s
8+LLfmzGdmEwJ/6BzlaCQjv6pAlzPtxPghdSS1oW3RSupFi55yyXwf7IU7gQILsu
4k+gFCRqlSL0FUWT+Tpt3tSwrNQs+CdNA2j1qb1B2jaVxH8YI0q5MmqioiNSJGt9
nvQyG15H0H/HItOg31xSYjg2ByFIK1aH27rOut38T3+5SLMyuhUz+Uji5BHf2n8E
Wk06Schf/YsvnOKTZ51U9MHtr/c23G70u6h6Omk8ff0AO5OAssZ3AGEr6kmtBSq5
jrq0waZtWS5GEA6URSVfxHgs9Ewf/A+rmXI4r4NOoe2btuAymM1lv798pMRfK8Rt
AW5R45hr1YQEOIuRjYb79dOzVrT7OFAQjn2vXUCQncuNHf+3Q9gj/ZXB1BDstMoo
NAumP/PeSYoZHXQ3k8omXMo9pe80TbHCpAKOnbQ5+F7wTRTlbg5d9piTuF3tFp3h
h72w3Is24RQ62Obht+wM4Z/ytJlasFigJDphrHmS2k5/DIblaN0Oth85+RzsOMsb
O1ZEJwPwuFJ9Kt/o7MYUbFuUremde/RGU/d0sV7km2MMJ1BUGKOkt0qw0e/FsNaa
YbLtgJm4LzdUisX+tmq98pk47aTJsqnnLz0Knu0O1lETGWbLVhQ9dxFTkcLPUNvA
2Z06L5V6b0JlmF/Dp+ZCqU2l9gJknKsR8H/+xsW3da0vHklsMy6qwWwY760s9myh
uBCWGwbGWqaUnZrh9bQBi5g0rkwUdJZ2emkwf73FIxVrFMLA0lxjCdb1qiT5uguY
SVExNkBkoPVZ900D5Y4Qf3ZLkPs5BIKqQhDs4EC42PPgYlAdgevNDAzPa9a8D4ui
hl58HOiICbCF1+IP/rv+70PuvgsgBHQ6Bj2NJ2prH3j2zGSWAhysUPMY1w2RDUt5
CZOcUokhoWBxLV64oIxm09YczHfya/NuR6R6wseFxw6Ouk6CFSy0gc6mQDby3kJd
Itj/i7a2ZPGYhvzYrIESOVRZtnnA4fOdqmXHZ3WAd16KGAjPNAiTQ+/ErMoX1HVK
36wM4ENzWWjmiUj8qN+pN8kJk36tgN+mJ0zxlqOj7hv+nF2SqLukQ4zEZeYQdlvS
SjXL3gicDb9f4GJ+zFe8hk6iM5t38NHznOeBdEeSB+qfb1kLbLcQFkfVVCoeKMCB
kVvJOxeiGPtBaiC25Y13zw+fpsdiJ24/HsV1c7qifFIdHxKQbcxe2HqLegFzFNk/
QpcSpVgvuz9by/AVtJ2SQyCQjX7ILEnAjs/fFmrTEvzSFuHAZpLUt9EMvgCN8Rxl
2QqUicsCoVZT/lwz1w+43AiwRDtGbpzWqMB94p3NqjPsfiWXxkrnrZf3fiXFQE0G
YnzMDrefPxv9ZdXIPIgkKIEvtL6MkpPIOHj1irAjBE4856uTYYAZKgcn0xlV92nX
gBKvHSSneWx7S5uoSP5uMgVQETF202tiKZ+pCzAJyQSlFEmB9Cnd7Kssh0x29sR9
ivAOsve5MvKJ1mxx6GTsRvgTGHj2LGNO57+fZn5QDxRQzTsKxiHTSyz7OC4bYzEW
r1CMraTjm5bvMBpWoHPrWA8VKrBTZpBB+1TqsJ2TRJyhgabdvSwDz0fYFt7u9UZ2
PQCExzpoNCotbxZiqSK9SZOoUqOXKDSZm94jQeprgc/LzKGKj2O0UFyDO2dWBufH
UOt6cgRmvMS6rP1Re2S+/IKOeppVP3TDeKNTeLYA+bQnmcbWQ08ijrr8NaBB/BjM
dWi0U1DXglMx69tBuAw++pIzs8iC+OMY80W7RSjjNHI6dm5fmgf4ycg63oRpA0I8
LT5UAIkGylTHDzD76vHN9xsgpaUy1B4zpdNxlRwaVfTgtnrgiaiyZZB1GA9WkrGz
irubdtc+UXcrIwLERQDFe/OKb948dRWwijs0OL/iyX3rvp/dBEDWkQ+miDcz3mze
W2LX2yT0YVI2+GjTOmzRBnCxTvip3X+6KRrlzbzqzNQPc11ngY/Wgf2iw+kycqXS
Svugg0mU1n9+2lODqoO1Oyp5GpfrB+CBmpCLznyoOeFXDai7tWm8FtB/GLiX72I0
e5z638vU3vRcxm5rCIti0uKsXmWg3eabpc5bOrJ4ESHfzAui696l7AeH1od+tKB6
MMQ/Ihl1+hlDoyuQDuewc7G/M8eXPa+R8ckxSEtZpwo6clkyvXc7g3/FWi4nLr9N
RFgO7+AzYks4a8BwwwqOCW1Dg+vsGC+WrW4RW8hpK/HN3ObXcbY5wxPev5HIvxPk
Jma8mp82JFfUlXGrwBVZP2YxsbKCDc4RQxPzJ1ND27FNt+i1gbyNgk5etyZTCwIy
AczSRAMebsKwCoUQGPVp4b/KPbuTLPwwuQZdNznFexGIWpSS/RspwgYgAjYp/z0m
zlbDUtZd4P+HaEV2LPV+NmhjECJTzBY66L8ypX6c+PX/5W9rpP0XTp0mqcHHk2IX
a/w+6lHYwDLNSZ+NCibP5/0JbNgQuTClCgmOroxM9zCNG5RNkX7QimVAwpkhsfFa
YW1aNmZZCby5MPDc0JWRWG8cNASASvCzYfEWa9nyCtlW/a7b/Q6GsviaKRSy+5u5
cKuSJRdWET7g2gfNhEtFZwlMEN0ZpohOzOmGAs0BR8hvdO7HZDp4qvYG36wy+lcH
p64yHq5wp3pMUJ8FQOIEPuKn8j6dyGQz9j2ji5U3N8eYPNSgsdZi3QGId/4OrIcU
Uj8BGmXRjzZo6eVDqIeOnkheD0YXafMF96WpnIUD0RMAAHWmrmxnAQTpeoOwYhkK
P/df2y5YZC21X78bRuJZXhsUTDhvPW6HR9lexvQnggnNKMlfj//bUxng74kCla5f
ca9/YArgoJzPRmTI5dqqCiSX6AizSrDUaT2pgqI/pH+YvtGGMHlF42uO/rdYA4ig
n88VFxIicgqumk2N8XByMewUXJ3EQuOj34F1B1L+zqQMjgEp8NRwHT6h+e+6tYtK
2wNYPxsmNiL1hkSE6c32S2gujIbUBuBoJkvpq3iKdy8r0MM3YbW5zlSmcXO6wlkZ
cKPESwbUynOBTO0PIPc1OPYoJPx/rmHK4SEjaaV/7fijeRS+YQi/lwS1pH4GG3uB
TZXoh102YLvSdEOTP4+6EFpje77PjCeYhPgJ1FqW7Y/ETAOCmY9lK7+d2EpdqeSc
xOQ1q1em/iHmVgHpOArGLgmrPbhZYd0Cvh/x+PusJ28FtvuXEuudyOJGO/ScmDuq
n5dsCsz4hevfaWlUOzVOtWzA+FJPzVL9rkxSOJdQQTuWayBX2A9B+LHV7uO5RfJ2
hjv0M2HmZJsp+tL84ML6DRm4dgJE2UbSIIUkbx6EENOR6QE5H7kRM2t0UhSF++fL
TEiy46x35gNjU+lUhnhaIMVZE6Fw2S+UzY0JwG3Aggt9FYFOSleMaS7xG46tFRBR
JOyjJ1ePKTTcn6EMP3Bk1LVNnMKo9XPbby8tr8gbpq7wmzcKotzc1BPQ1dZxIm96
KVVEdPrlJADVtLesbRMEXPSePL0fCLPXaE3CB/3SZ0iXhnHVvCnwAtVwU9RQeCHo
4qNiwgW9e7OCKF/uJdX1q0JjsNlEyU+I/tyuCQDfLUvduTVm4mWdS3JDtoAr+ORF
7hSXWe9lHAA1fQB2d0VU8lhlkrXatYZbrMZc6cNQ05jbl6p6HvwutfPzemC5a+2v
zO5fKdzBwU+vGpMKQufLnvCBsNqxhje5Subok5a5CDVF1vagva+G3DdD1z25MGES
0WNLrP1Gx25l/O5QVDyVaYBjs+qR9BuNjpL3sGanuczzmli4RYE8oOYU1Q8gf/nR
xhqAtS4PtSBVmxVThbA/Rm5nbh/u4UidpRPAtE4KHRUfXeSUGJDK9lRKev+Xmy/m
Y1IU1C1QiCcY0kQnrR/Crwmj6ofabCnA0IOBcNziyZGTX3KICvlislu9XjQuwRSj
ecTNi4ZdVcVnJSsxQj5WHB8Z4zrJBIGXarCyIoFnxKmTzFkZC/5KOx1Hc4rIp9xI
gDAi3xQkGkOprRGE0X4DYbzbF1nrEeS1FBf6S+THA0BC02VGBFgyLgvJTKSYvPWZ
FfPlm7B2KIRx+Bc1UUohZEBwe8SPkjlLoeYb83ZFqp2t3X6hkZyk1pFSn1MhGjne
CtlCXcfyQgpdTPI9k/DW/sP5/hxxJp2Pm02mpChDsPTIkClRsauC47HRHvsu5E21
ZfhN5tBzmpZ9IwhgbdNE2NLE0mtbgqI2q+laQXXqjFSmQvn1fkfLWCAnT4goy7rF
zrxcCgpJ1gAIl8+jEjlXtybH4huILDeiz5Z7hjlZcn+ghWH1VddjlYCzEcg2j7Pp
N0/Ii4C32TA4kgrNFsd3Y+7mrJM8C3VIuH/Ru24tlM+Z606cjD4XsaoyuW/5fsPq
i33Qv3XG0HxrjLeSyqJathzD1mcQiDb70uPlf3y/VkxBcdtZsvmSDOJoE0uo255S
WzsXIG4fkv8BMFe5rPtkZLOGtIE1PU5oHkOEDtXcoPGTJQlPFov0gLdGeBWXvOI7
QyzTkFmM0BdKa2zYdVwbrsr7A3azs0BxlUE9CSe0k8sQ/twSXR36DFPF/mpKeCWv
O5ihmHtcDC+i99AYlR/h/12dSkhDmo0Cq4d1inWwkH4ueZuow953EnuTHnOmVszf
qYia3GmDHtYBUytcdI3dgWf4tImT3vxuWKu19vKrrKrhFP8BA4crV8r06J2O6tLw
IUL1Xeg5aS3lxmWohrLP1MVmTHa1Tp7XFPvTZN6jFiy3HUD9Eoeh0txF8x/BpkFi
iCblUNG5YXqxYOZiG3GNaU/Ru1SHs0X8FP3Ma0cTnLhupiZ60KFCEBt7YqTxk2KQ
s7+2iBYfWYdyMhoZHEqTQb3VgGmSKwV8HSLHV2W00A2UZDlgGceMU/A0YuUKKzbg
T98itGiql0iSZt5KgDLBMzX5Id/mJoWORvKUQKX2aysxBJIl5Cz51fPLYMkp2tEc
BzAaXWUfa0JnFQiUux4DuuQlC08opxlQGx33p7DXT65o7OgztwZeZxQ5pDxmoGaz
83mKqVKiOvsIpXJon8Bpu3n4i0VsxZtg/g+u8ZTsFbV//a08PG2/JbTP54Dce/md
ngiL1Wjpty4mYdzxWwSn4cDKDFVq34IYigSXXbKJhDKKnwkURJqk5eKGcF/Z6D92
4TQDqX7sASB3Qv4XiXSctSbB1V5+WZHyXy+mqB3GO+7u1D89dgfEx1pFFLUyTVji
oOtecSuXXxGNk8tdGuH+jW1hW7ZFzI/kAHAa9rXWmvhfByoB/l5CE3Ace++3hccZ
jVdmOdEWl83Fem1duM4jI3IIgHGfYkeH5nKIeYNwZegVfxBPskPbTNEDSmHpzi1+
EO4QSxc5sTugTGn3TKXYocyCDSoLDygODwbWz7pMszdleWWFhfqtMxTD/2TZmUhk
CgT2VtrX3DXXIA7uEtEWMMLSCndw+lwgkOVWZbU593xHX0mjc5CM4NMhwQ8rknhZ
kfGQiHDwZ8gv1PBcvcT3qUyZPw5y9iZ0IurQNYrpRJ3xrdwwfqno5wag67psgv4w
HDw2MNEKRaZh7OzZZSbwR8InPm9MTHSGmvNm/qwWhsOTlJmkpTrRulVqo0sJlXR2
sJx0Ao7UAV6Yx3QQFN0+aatsp1rn4NR+XBci7q4x+yf3MNrA1PfPUBWUHdzbS5NJ
Qq1d/OpgWP40ZkB70ODuxgiF2mYBqL+coYHcWLuOSGlFbXHf1xFlhA//TeUq0xt1
LmcET2Td9kafKUTxIXCVijbgBtWFDtwdlOpfFcGf7W2MwpkkUGSi0KtNhBhtomPm
0kcm/fqtD8hkYAh54OWkzF2ywFQVQFG8TYAcVYRA3c3VdrVidq2Fzo5qq1n1Rmd3
/EQsFCdx8jFPqFJ80WjmyGdGpAxdETB9v02at5T4aU4QrdzVy0EPpBLinPhZmuW3
24Uo0OmpQuF5dO2ZPOdyIb9f0RPbP1zVKkNKFY2jhNQYK01mLbbg3YAEUgNNZrPX
21dtVErrT4YiPVZQU8cD9kMOIo9LdjA2FQYXwwR+9nu53aXX5DmgjlaDH4iCrsUG
EvYFuP2vDUd9fTX5qVztW0ZCu0Mr8vlMCwOg1nVJqLRDwqkVbdpPWuqpJHEWYjiT
5/7e5c3M1iqMo5y2LFV9bWQpyhOQc9IFUi0XBVBaHwKLXxTDegtxva8kleLkLZ6h
a50TqjUkjTgbvQxv44qGSdPg0bE6MWisfbD2fHpn5SXil1TW1rbMXbWsEUESAR/n
yTZYundme2YeThfG+6Nc/CHN31zbeAircJmdEYYydD0PLwo7xYIUBmtdhg1WJf50
OI4LEC7tHbkC8NjohzP9rOh7hM3+14YCXI5OF12YpDSq7nvdSppn6RM1/tDvVED8
43d0mNTn2NzanUfB8ds3nQdEG1GbCcyO2UC+PBa0BY6edb9bFpRNzQD+4z51k5oE
NFrxq/YFXXXuM2Xh2Kv0CzfpmKya9GUvvO+118a413YKyhRmf7Omc2T1yx8/+YVC
CHubsWqTEpzMmlyJ5wnzF+DBiYBfsDikRNFkx1nQtaZJZn3qvLUSzXxCgFB8YOMT
UP2Cb+IRgB7YFiGAFvWlQzk3eTkx2YpEQ3u6CcFm7FcrlG//okS8tPpfSO2hIIwl
g4BlvKx9prFjWZxKpxbzOKnTcztiqKuQ+xZ1fFtUQOxeqaqj3VopGP0gBX+dYpmz
VyR2GmdACt8o1bpVs5msrkUGSc76EUEcjfacwJTwZM9F62GwX9nfdlEuH4tPwcMj
/XCDkem9ioDNOP+G7FJucYf85cYJTQGZqD9rSdekrnZDsTfRHUzZQ2jlDResmsIp
Y8V7kUKs8yw0Lan8jBbVcEQprdePUh24YJNgicuEpS3999j+qDpkka3Uh6OI221E
5DFQ68Bbphmwjga1qvLLGsnfaf83n5HdYVmmoWtd4t2HPoFXfBvSfmE+kFIlBmzz
On7cDDPrQGDdSg+mJUWD98WA4KdOSAWtMoFb9jjLyxIclv4CYrfQNXuRm0ON+NmC
Q+uMzM/gHCQTmwe3gExOa4/k0wxF+sm0SSy1xuX+Gk/YXOsLQTV3msD2B17Bkjf/
8D9974rV4ty8CliXdEtlkMbuOvnlq7krS1j/KP/a19TQVbost/iqtANL8GedVqY8
kSH8TWAOS7mSok+Kb/2vE/sCJ2fR+r1+aTGSz2ibmvkMjK2k6pAqGPokQuoRAaBF
3UOVnSXquDa/+6JxKXqnj14mPIQruJG/Cnyj3dbUhcgUCpmI8g9HPlxTrTpvQdTn
l9BQuC56Gc1uA/Gr96ULOD0XxpsnM3nzwjn83pZ3bSm7wlJ26MONhmXpHC7HYpgv
UYpg/tgjkPscVsbc3BgLV+43gVBBFIelSixkhcvam9m6c7FrSeyItaNT3Gl2JJMy
ATOVk/kkHkgf/CxMP/LhEwFXgqqbQDk4IOEPzV7ln2NLKy7MwvPT6Nq0CN5PV8cM
WuRCKXUz5uL+poSlpxOkA3jHXiKSYetZjiEvjqIEQwhZ77gJndMgFJ9D+4SC4XMR
Cqt+RxtSE108d3w8N4/8QrW2KSXlegJZJy8ydFEDVpSHlQubomZ82gjVkiGwIg4w
WltyLFpK+xgvmlXc4wghB06cX/Q7FTILCUlCh8j/0ekmqvfMpBp9oSYD37PQwIS3
QDpr5GKR6faLVzRY/qpoJg1kun9VZhtFN02KqTN7nisOvIAfcRsH8rMpZOEeJ0Ci
HSAC6gni40T1WCeBDvNsoYMHA5LEX/WpbjNQyecqJdjSRqUfdMJDXPoi9jCjyf64
LzVArPsTP+z1ynp5tTBQuSK4AWAZLYy1VjPYNFZHdpft1HqPGMeYESc5sc/y7k6Z
WG3J2ZrFImX8lDna7I3sBtIsOHtAH3CuLf+ymqOdagrvCWGjg5RGLDnZge3D4OjL
1H5pV8CRf/LP7YdDetlHlHb1eoaHPAD81WUjtaENgpY7rad7zBXUeclVbtTIppGb
siddb9V13nB9j6qp1A+RAilc6MT9G/U2H16oS+QWCvlU2DMH96IiwM7KnlmfG3R5
T9iJcR0TdEtrW7lhiZrP3xL+4lVCihzKYeNcjI7exX+l0/zTso0s/zZOH6SRP3Gy
xi6NOGjRwqGnWTyxnUs+5kJuUcgMUbdlaihwRjhaDeOBaDpOMctUgQkfb+IzBXft
40UaDJ+TkStqHK+5Kca/BBlR7CwEJ0hKKSGgwNkb6cHSnBcQCdGZkhsuYxzrWiAi
ApjgyDpmQase8YnMkCj4TUW0/oMEq8RiFjzTJqk/er3Q3tW8BDnjU5qNTglapA3L
OLTKPNTfJARMphyvNqeHRu1Y/llg/sx7pe9g7MOkQT6IqJzAjRctEDxXIzrVB1Rs
QeEboKhZT6u+RLSt5rW6Ljefxxjj9rRDhkaCKpLJ0nZoCxlmlQ2JLMkKoLAoc79k
dX0CfW/2Bhhs5WJ1ReGxTq1V5CneLeB2QrUs4uxYwY9qM/HsucOJKE5sOMWBC6+e
gLWr2MzBTors4xelbxm6b8fhn44qBw+st+BTsveWsxn897nsxTa3iY8ao/DiLt2i
vb3HJ/jHZfnJQ1RYDvSGoNfCbhsXZPQ/iTIMWVM/OsduCQND2UV9Amjegv8/71C9
IZvM1PAUlYQp5E3gLWAsvZvTBneMOlI+zWFxzLn3T44xwmrtcUL8xXVZzey6UIGR
4Z41eKbj+qCr4BYGPSwBP4GTlwj5Yzli+BG8ij3lau4tHk/Kaa4zo+2FLV4Arv4v
J5UYE2Hh+kffrZBtA6vasnhewe3NozvSaj2uExWIwJ4Vk3yIf5I7qE3IQj2PhagG
QCBhWw7aSDxcD9d8gDi7iubejOVnwHHVsORwmsE8O50ScJ7eMb2FQBc9/XVkDF7L
Bhnl2mrDbTe0eQP28KMFUGd4LpTNTfAvg9jMG8OBj/prz/DMXzDMAswY+qa30sKq
nBPK/2+9iXHdiwtPOE06sUuwKUlAu/lfh8nQglsg0Jsq4tNO0B8GTeF6eXeyOxEG
BHMJz7NE7vl3TcoYLtW6Kh/6KGXH6tGK0sumTF5aL/paYDury39b6+AR779+VXD6
Q8B/1EormjH6VQ77GkecXpgBdOTdrbZnqLmShEWPaGnausxfHfC1eQpsu/c8wlRc
r18V3ojbxvkJ1PgRVHeAvbGkDqFGap+4cqZZLfPjU7Oz54BSXoQsIRKNkvhYBE/U
h+u8zo6ihFVDzSPjB6wkSAV81GPYqHugi7LC7bnft8dSxr6sfob3FXaV1Ij3SfC3
gcB1xvW5VnMYSiUf/+j67FGIQ91qX8DJljUv1wJb4jOizM1NZEsDVDr8lKHV0+DN
1SWUQf9VaYB5Ls5bCHFY6aFlZ3M0qBixvRiKgfOUzTq+cvAgLtw8/nIK51AfvEGL
51nuUJY5/IecPwGEI9dJU/sAumfrtoPvTxgvSQsmn6eWZmKVU9ZQzuVZUEJk8zlq
C0NSPT0XU00GVrlNfvyHElTeM642EIXO6ot2ARBi0lwgeLMqSIxdnbh+XhQPp7+C
E9kRl65hHQNGupvLMmxamxNqBiqewC6byQy/XgRmvhnjPMlXa7K7PjnAcXG2WDt2
yKgkmUjhbc8MyCwEavp1D0ueGBccEbQDnNbLwViuVn2KoasCFeQiwXclWb73YmC2
tqzLnE+Q+YAD5cx0Lt4szUCf/ehfZa+ug1FvEnZ76riACToVYrS65XiadJQL73r7
1v2yeVBsYK3fB6Iu5x11pEbtZ39ERIeiHySapNf4hA6GQYuATCziXR8sr5MgQgIW
w65U2UTN13+qrB0A4vk0LSQs4xHIH5IoigBA0U1ze7piaTANbm7ovbP3BzI1qHFu
qBYw7AUotlmhWtJUMuxjUF5fa5nsm+pGG5aOTmG2w1CNhXnZAy6blv04eMelOJpF
Hsp7kFjO9aS188Jbbij8ekXNZYDlupLh66jeOz2VseGQfNWTpiFzynI9UULRrM9s
dmAb01l5W2dq6m8kTnHsQycjmrT4+2aBf4vT8BOzIrEOf/bjM5mj9BSovcvaDtYp
UZZAvhrdDDG9Mie5PyeACdifiAR9LlZDSIZG637KpgGRUtvOBKjvWv3E66vpDKyF
PuAJKvcwu7UHzE2LPEXx180QXbtEbX64Vkpo3nxCvFoHzsWlOC+Abjm5DsoRmQpz
zPMwNLzZYcBcFNNo60JH4GaOUFUiRlvWLchcW9x3HTfD5R1FmKwZlix3BTeZVcFU
CcDwy0yewI2/rdKZ+Pu4zo1kX5FnAaPlGrAe0MMa5KhZDDUd9uD00CwyZ+T6/U75
ZdcgL24kK9VWo8hVfjsicqUI4JPlbLjyFnMrVaZD7boBNkDq2TF09v+mOGnwLvla
6nO2/IY7CrWO8hqGgAAfluvGb188HyT8Sf0+3bHlxQcphizhyTf4uVTiAAvKp4to
hV7xxE8C163/yGWkbyxL+NarLxK5U+arf/nf+oKiv/i2Qplrqs/Kw6PLnDMMpzD6
KSgiCB9kHAKZXjJKAz0suVSOasGqLyS59O2n2Hpg/OiCC5S1w84IhgVSpCtKbREt
YQaMayI30x7jL6nmihiK0jX+p4wI8ukVvRnhv4vaTSXlq8W3JXexfVRUHmyB4RSI
yxScyz1LZmrBYCNZzoy8HiyNfAhupY165o+JRyOBgri5bAeHZFBjlGKkYaaglSzb
Q4t7vC8GEMEjmiJrHKWg4FNWWW7OrKA2ozycnA0Sh2+mzMVik7u3wfSbWgpfPkDB
FHDuQQgp8/7kYjDiIpXVNKXjaWp5kAUXMhI6YBvzfPutft16+1qH44hJFxFj69MD
4LzF5NG2prukqYq2bg69KlBL85mlTqDD+vhOj0enuWxj7lZRWT45+60huzaV+5cT
Fty+juMDbMbHSl3e/fxl7XZymledXjunp31MJH36uunNxxC43pEUlVqXE7tIu0DL
AxmvRf6mMsVmU2/fyy/B0LF51WKWq7V4uiaKEQyyA57grW1wBxjRa8X6fii2GdUY
gl54ct65PBOKIyzb5QyivMrMVJzK1euseL9oOSQncPoihBjeFj98FQWXHBHHPjDZ
a3bhC0UWqsH8X2Oaa7QAKEZZfy9/3m6n2A87+hZamMTRWekyT7BkTOoStIr0Qyqz
r9zjAGpJ25ORKcKmdv565Y0YAieykD1yIuxACizzodcmiCD3QhSux6jYg+IcjwFn
2884byy7qDliYntz69tEEix0j60KYSKsFIBSKHc+689yd7iVewM2XrU3Dr8bBnf/
MbpIf9p9kLvEr0UViZSFVdYRPLHwRzviX5FQu/J4r4XTD3X9ZC9t9boav/HLuTmu
jfM1Tsu1VXUv+LsB0BLUdQqmlDnOdsnjvpXjCJmc9bT4mhwcJUA21H1sldQF5qNT
la9dT9e7KlbleEK572n06KuWg3v2VPTzkSu/nuNLy3w3oeRRZSew6lg4znYVu/rb
t5h4M5hOHC/GExLo44hZboUJT21Kf5bKXYjy0MeyImX7KZO0BqYTxQ8Eul8BGLLp
ixr7ZiuoCwhN4PxDyFUJ+AQtd20Vy89b4mdp0fjzgfhVbcQ1SDah15xehXetN6OW
kWn9q6VtdE+9kenR4yF0rIoh4fILPwaUmnCa5yvdvruryLNOCGTbyEia+OczEky2
zk5RZ4uVqonju09EguKVVvty/oKP9vYoHcUkAxZm98RjEYSZEVeIUZqQ7GyZC5kf
JMGkybub4guWtIf5KjJKMnyEhFcdfUasr+q5TMbtnhXiej9HwOBB+pfWBrUzrXJ/
v/sCrJ8OgZacvBufZZYLjKKHDudx7spjV4+JuEujfTYfJ66pM6PVGiPr6WQhgeVE
k98TlQgHRFZgsJHLsWq9/i31h/tganxSGaTaS1KldpAA/3VqFKkbBU1Rk+A8De9n
SDE/OX95k6f07lFH0BUJsFXmmeXl4+ZwupELSwSKMt47ueQd0VD32ng3E8YFXesz
kjqGKkDPOHZkyM6tYWbjz3zAZGy9WruqqlpXw6dFCOATrDI9fKPyG38QzGhZzLVV
S6WzDjbHSlJr+h7DEuT2TjvR0yPrpnOV+M9e8DX0YBFoYcwIc8RKflaT/zA+oHFz
AU8XqVM8jQZ3pcz0382EFvV50cnpFTEfHP5aVUEASwGwTEYYVpUwcoIsH1Tfv2tC
5AdYoc9Sf9vFAUCT7LZn+iTyoFPQHArswDDdobUEBt6ApQqAnKYSuMVmyjuIKm32
bMvbG1hDF7xRwn4+FzjViPnbPYQ9Hyd7WJSyzoDAZRx9AxeTcLv9N6YbX7tUfigp
qylRDrI1cd4VTi48MUaUunEU1H2eqcuMLjpyfXj5s1VMex2b5gRApEkKBehwGf4T
iWLdzba50kKxv3TBxrdvlGUpoM8o8lUBkQFFH+hB6h9XZDKuvJor4Gb9OBFg90hT
iGW7T88qlAYhRhwMwDBhKDzw+WpKGl44ykoTu/eYqBfVAgBbf62lqjJNd/9H+fQu
ySov2ab+9/1KB7XpHnNV0TxMa/joHofE+cglWvTr6R/6we4KCVsQgjNpCTzbaHvv
TFDTT3MTouVtUZTKhrh639EmdreFeOR4rwLTB5R5/PSKruOqVzMcYrQoIg0VvRXZ
mZyqYO0FvwbAFbusMdEyqucrN5/4IBNftt617WiDh15uK3GA2PSIs/nSdrAYr3kS
9wPAvGI5USton3iakPiyfOZfVAXSqxaBhxaRjltGzH9uilZwc1SrkGiO8ddcxFfK
xuNyvd+zpXYoRBm/RFcz9oMkRm0hG4CD87gdKMUBmafgyOr9A3iBtmEA0AP87BIJ
AkVd0le5bwS/Xn5K0sjudbBtd9+5ioWilcpEGlDYawKkR37uIKoYxq3N/N6RzCsD
OxAK0PucwPNn/LI9Fx29bGberD7W3bzEY1hvscaTwjqiedXIvWUjI3Ib6ciX2phK
Ok3noExLEPGuRNg39/VxLcAl9WosFkh3Ue0wXWxQ2njeBI3dgbidudB8WzZM280F
L92hJLa9fyhKD4COLa8N9mu3mlslzc/oO3nzKeDwL6llQMvnXgLDg+Ru6ddzMnno
mk8uE34ejYoUMKucAtEF89+prMnDhe4qJHr9pxTzskemRrAWF9oOsBx+4oxQxj8P
v543k73HQbfgpKNNPO+PzKVnp6j2/oSrV3XQE+pdZ+4TCO5Yc1l/hi8SV/0DglqR
lc+45IZoJ58hlfjkSJrgEz+v+eMMvpDoGWlByjkvEhxA91jTDkSTBrKXhXdQxxy0
9B8NjguiFbVxkk6jmEYBIxV0ydHaN4heohvjxHUJrVFQyT3y/pvySibaqIEzy4JY
O+TdNXCaaaLGAnv3TM6cUOANl3OADcgQ1T+0oztI8rW5rOc4eziY6sKoXOWehvRK
D4Wl7GUqn4H3l4LpoeMQ+vzb/heVAEJTWvcuyN6vBMUwZEAi9t0aj+XQk3sqjxqN
NYiqtXaV5YsHGqq2iooV2+s564uB6k95UeXO15UupP6WtICVW9VuPyJJULfWHaZR
CYf7l2GP7U5AXTrsk1vr7saEdWqsJcPjBytNPC//DZHsYJ+nrWoIVX2uv+K6jehe
HG/BBxWWyfO9YBN9XUogAu46dhGvCt7zGtPPti+OZfq1v+C8i1XWfpRJy2eH4Vxl
GWLiQpEpnLT5MI5DlIgESlRuOH+Vq5GIN+ZpX9zd9cEvRAkk1x7y143434aY5Kym
LcUbfqwexI2gNTbqOuwbAcmIW6tSVsgzoJdjzTPzPlpN1UpHZSUgZi3OpcK6E3s7
5jg/K3xPUfjIz1o6xXcCs1rHn0gW7pqdQG/N6APNG5OVsPvYcQNJDswFqY1pGVxn
zjhypnLYsW5XIp8jZTmgHaAE31umVxR0XrZRqvaDD4T0GDbj/3raBbt7wSvpQS5F
gLPbK64nq1QA89Rf5OE85FhSvpCF03clv2N7cmkd9ypgX49QLzaZJ/oOuiN7PDHb
iACQr88K8TmLImQab2yQ8NFTf3fLuvFjrK6/TpBvrUsMuZzFWONDsMiv4HeuJ4rh
Q4XQDwAe1I27o6pHIwtiGErgakRQvxK5Jf/X5ddgdXFAS8maQgjBxfj9C0cGDSF3
pXWtOhiaMc3N1lJOGKKKcyyVIo4xjFTiaCn7HpD7rjGqQlTlQB2Owl5ALGX1s0a2
nbKl5VEGHoq6EoSGlrHZGwleqweBD6HOpZZXdHDdjlrtbM4Ix4dNePyCBAz2SVND
akGMnmvssfrHivdO24ewzweKFG+UBb3yqsN8SeUapLqiP/O1Ly+vxTYjEBb1wO3h
AbxrYYwmG/cqvcSrObqSzDZn9ugoaU3WU9naVLz5W86sVUkoHLD6Vjp02skBKH0N
tvi96YWu3N8fgR2J+HK1MyM0pKuA6NOoUxbBzCNNm1z/4q+4Xku1xX9REk/WdypI
CC3g9IWtcmrvwfOgvZ8Z6qM5PAfHYA2sKBwOKoP1apjJuiYFga+wnUwi6hRSsNVO
AUecwWPYd+o4G1TzTfOSv9evN3bnIQtrKCa5gk7qvrixB/VRj38b/NsJx02Iy6JO
taeHd0NbnrWual9Z1nfFLQwGqvbwd4wP/YQQ016vXU89LyFtEl8BCAGj0g0G7Ymo
5IXNiEzzbHL2eBfhtph5OCWv5gn3za804dJbrMH17YiR4tN3oECpWBw1BiIQ7syG
lxtIKPPsuoTYOEbSPmgATwn2vIzZh/za8TJCu4nqPEqYu/W1OgR2uopQrzL5SL6h
WodgxvrM8Qtb5E7iXttydD8zO9vnxPbsaQMp56OycoctGup6/p4roTNAqFwtoxiU
cwOq5lObpKwAiv4IUnMrpdg/zzUaRem23WgWnyicYItb6mzKFKm2bEG51aERK2Lf
oREH73AX3eB9JHPKq36VEaOMfL0OBV7SYHJoqMuSXXOjKacbcvTQz5hitm2NIHfl
1q2D6YEcTscUJyK/Ty8uEef+e33an3ip0IB2jT9bHAsbxX+hktF392aYe8xZXU6Y
+76Jq5ItkpCbOPk6gIX21JX4F6Dc4uPiAZ/ynZ0uk2h2oMhpAnIxXko9+59mSQAu
cYMiFMHH4wMlveiZqMAclOZ3NqUYdI5XohPHG7l/1LTBhZm3RGSX6R/eo07N5F/B
b6t0qul/O/GC7RZM89xpLWaeQnru9b7cP0mRf22KCHypseWlOjMXjteIcL8y2GKv
5/12b6BbPycM9ti+LyUQP4FyO8BQGSv2zLe1qrajhRPOdq5ILhIn29uUeaaI2NAD
VwugNHxRL9exdOpFtBGsqeX+29IkiCa3vTtRsaMxBiXkvupUDOHviUxXKS7YHliG
EvscQtE4Yl4UKgyU4hkFLMAih9YNrk47ZVzLjf+Irpt/TZD1P+lBwzySV46epjqr
01Jdyp9Ge+knolO5gMnakWohRzAhsKkfqQRUTNibEzX5x8h0xpTYNDPbnCzcOYQb
7lS5PACnaTtzF3fV/VAXsgeuSlB0eupxEp+5cJRzlspHjFS8u5zqXeaCiOCAbgb6
zC16CQnO31LMcPpGXebFkrHkBEZ1yty9ei7fcEDLyVDMUO5PSpxYzAOJhlQKB48u
e+vA4zFJ7bqwGfVxA7xluStwLGBdMZWjkkdN2TDTmYvC4/RfN/iAXoGOlp8LWAb3
c+6oAmn32FbWSIaDqNIznG3kXN7mQDBeY1AE2pH1Jd2VC/gE7tl/Uysxtn6U1MQB
gjsTpvSTNjqAN7pnujE2fxjS0uTAZgfhNMaxSQV5rC++CoTIPPgy5OnvmDCYdXvr
V4Y8ioRmBel60pe9t1TW8hTOy6fdr8e8C4zP/f0cI684wKWGbPj/9qYLWn95W2FN
3g5a2wM8m12/PONdrzd5ovx9gbIagxgqZA/N+Dcp/zWfrVvfl69WAY3P2ZHk0Oja
b7N0G6dcP/euhLfmKKvjw0x/ZEmIZ2pWbbxji5Zgnyl/gD0oVsrM6BoEoex61sH8
yxntwbJdPnDiVICdgwY62xXtSjLwF4dSWDl5oIHQNB8yHPLHAQa7yb6ZnmBNyyW4
gov37U+wuiLles4gUYvVPrzP1QYKqgtO+U1mXAqaZt0OXOc9hSBz1DvuqV2jNO/G
bw6Ms+/sfC6BLuFggOOLPvXRWj8cn3ja9Ph4gbsYNEoB5kwyuzh4hZTUa92xduT3
IDzeI6Aiwuhl6GdHaY+5ITKdxTbMZbzcxCsReg4GYupgYXrDMSB/zCPuSQWKr5Wv
bLQwGWygms8nal0SpagV5sizmkE8pQLQRGP7cec+aQ+4ahMMM64R0oO39/bZvcut
smVDANipX2V9728B4b29VRXqKAKwLE+Stj9v+Bj7EDFTJc+JZuVArapCYwxydAFm
FRNqaYq2hq5+TaIt5VxlxUw8cKISzpMIbB7aqJVKXEXm5SmtuHDRdcV19g5CrPLd
F/NJBiGlvqR1qm6kLzDrOwcbqE5DDvQK6+hZZmNax9jxpseAfxTo/L0sKDJzsD8Q
v64XVv+2y84z34oqMQ8T+zWlshssjH09xONZ1DeWdekdTo+506Eg1aDQHp+aCebY
fZDH9j7FbKpzcKKx5tqPFod7pij6f+QtiRVzxff8kEiVZ3TCL7OnIg8OYq9Rndil
L6ah80igDZBUmFHV486NLriLW8NxmmZCd1HdComEPAMKxAfujcuygD4XmNsSyrVR
CXG4reYokSB1nynmzhSdAaMHhRVMM4JC3O7ypyBqtn9FetfBHEnu7DPjhB9ivU94
On5h6mNW6kggCpjGAInkFXFHRWslqx/rcK/NKtF2dimgUKbGNpfDmKaKKbkoZ8Yj
SN+H0utj+MU4LYBLbfzEJJM+dYe6AY8bTa2f9oPA+iqdjCRVCyNZkuwuA15vpU0j
fULXloOPvcaQwwFxJ0oGA+fiulCF4WqdIZUTi5GnyG1boNcEbv+xTD1h/GTkVpf4
wmC/0OOJZ+MNRB5rHlvKavOGGhxcRmDFX7htosRFPnqXfrUeSdBgZTPTrtFclq8b
Mjk9/RUEGJVpHEf7TqVGLt0jUys0dI23Omv4/jVj0gRyuxDfWAIJOXNgYm9zobsm
sWLjdMAszv0kzAK993f90kBXFeo316i+3lLHOurP7vJuqoDODqgIk2656utKd4ah
/adbt9s0o09pAu+nGVxCQio3YaahSVsDsOZAcfEpogl9dLoF3mKWNCexEJeAtdB2
HDLdLrJx03ZRY0+Z/OQSEkTB5P69Vuc4ocZylkHmQM+e6KBRV2L/K4njGARBBghv
PdlYk6Zd4npYxPpj5BJ6YH4cwipUAQPNOPBpr6jYzEL9z6Yc7kRgyeNmkyjhpHv5
MAD5NNG+ob3edptLGHvN3uDH7l7qoZfYqFxfjOBBz80GpnTlezIhMmTb71xmcFL3
z0r9mrJgl0moB8WVTC5GffQejBZxBio+fRsfZXZXSaNnZWUDWgZ+LFEhxl7gDieH
mb6PU4+7NeA7GJ+xuneWKbYmVUUP14H0IwCgxaOEMroQw6cWRYKhSIgJ9lnD3p78
i58nJURHM8648ZPe/2VJ596kAWoc3S/1eHr/l5HuauDawRCUxgEOwhZuWji6PaAT
2BKP/LJxj1jGFdh0HN4GktoNfTXj/vPMGJL8HHMLHhFY20Q174sqIUpS7L1W+KUQ
hnqffhuH5wNdVayx7BWjMr4jyw+WhJjGC/nIzgL8o+eTDnk4CGrAqa37ShlxuDSg
2pvs7XEDpkoKtyPywtLTqmjgkg/ADuJpDgXSWr2irrT2qpAPuiJXlCYdWgsCgRnK
CbHYHo0saAHhS2ilBGKuGMk0WOuzjqC2eoXHJyJeMvL3c8zEAelktu1Mux2F3bN0
WgmxjOqjV789Wbri/jFRcrmYs7KRzWbQ7eI4xBuLh9C9UIF1PpWjJir9CCwbWgQC
5+kn+dAVF/lEPOerDYlHQUkzSHAalKqTJvE4HPYq0KrmyhnXurzhHn7NQvCkzlo0
rZMdXBc9QGtXCTXhcKSBHIMOhNf8Xb4SOro2Hx53BBhTyy2Yeoa+UWO2FgW0rTbV
9BdWSRiI1yoLbLTpSV0X0X0RrENDWWE13EpesakEo0NejrQZpcrPNnunvky4Q7zn
uC0SdJfO2yI+ipFP8JpnmOOsxP3U4u3ZxJDz7Wq/qok4H4tdBilKQDTmq2O3vnWj
+8OorHI8fDLAM5jA6scyEeTVjBcoV94ojIBAcjrb/cyNCp2CYykx8NmVlq6Pm5Gc
BGs3FFvsuofFidcftWB1XXbHOKq/WC7FfawZi1nR/GjFFk+hwxJ+tXN3DTWImqLh
QrF7ve03aXkJoHlogABj24KjeYG6Kn1Nlxzk5Q/Gy7MhuV9a66jsTZqhnlw4ps0C
C8fJFhwKQ68L/4dvCsoHJnu+rp9liBUUWsN2I2JqqvIr672NDt/Ha3OFyXn6wFLy
HOoUoiPbZoLA9WSpY+nx+qnXXN0pjeDVFM2HgoE7RQuFEPCAOmbCfStsorJDqLmh
tR7Rc3StWcH1VGPrIGaFgYyEx0xImx9/5ECWaxC/frIKHq4YArB2dXioAWOrbBi7
ntkuRBiZGBUezYOEG4Xib5Z2XP2sBGKnqEd+f+e/JS1DO+TTG5f7FmoJ1mLyyWll
GzPR6Cem+f4FUTfwTnKr2+/sT3yq8wld4XfpeGv1WKzo2f/DEJTrQ9P/bGZxDqnp
uD0MLXMVmUi3yf6zarcCMt2zaf/MuJOENS6gaJso4E7VGkZM7kL/7bE2ol4C//ay
+IKqheNAxrjfIQDq+Tk4hwy7gGtSJqceT27HmsOK7nQi2ZC8kWpgdE2UXnTluxIE
uBfjnXn2fy9iLduThLR4vcCtxpwsUPiIsSjUIv9ls7P/essTLWgZbnm+ksv/gTt+
oXo2Ir8VZ2KdtGQFfx1qOTjFagaxTFdBWTeA03n0ZVAa9aWO6bE+G8pLQeU7J3Di
xn34wRRyWlJcGVxsbTBCYpD9otUW3BNpZiyxL9pRcAnbD2iV5gc4ndAQwnyroyeM
kly+8t49REhhpVK6UwCOZmr95TzR0F04h1z7WChm/Q5EhBgImz70XcBABnWW0jLY
JzFPCxLvbJEPahssCFYsAzlBkJgTqIZfax6IUXIhhoO2v8VX14dl+LecA6BJsYzj
8Fs8wmMLHrpQ/7suQASzulCTjuB+1X0r8aXoF3DN8tKQ5H2uy7OP44xTdBCUIXSD
TOKeW49KStWtycou/xMDYt4XhojPQ1slIMZFU8gOls3p+Iavz+Zg4eccYEO4yRIN
V/tZtJ0+lnoZxUSBxSXYM32Yl3vCe+YHkYiRCKIWnDkctojDLmisvdKjoBeLlJla
1nLyabpMRxjUKXgK7kseplIPBD/5PsvpNGmjZk8kh5RBaNGpNrt5ODhNA7o0uRSp
knI8i0ED53uI+GVWlvsxFjsX5QUrUwL2VFB6vU6Xk/fkY+uGqLcyF6cWFgmGc7hN
7mqlunOfu7A/LQUr6ZUpRr4HorgHwlU84RtDrn/CEg4Mr4de+LvAusRD8Ky3Am00
7afWR39E06THqQSUqLzASuByl0FOKuY5YVmVNKQXbK6S1DHb3LycntB+uKeK48OW
4pUaIpIx/z0RObFSgHG94q2KApTXTc0MUWLA6ga6ErgTvftI+kuVDf+f4zUWubZp
Qk4Tq/aLGuJfuxcZFQ74Y8gpjwPQLLUiioSiJruPZARlxtshn3PfOC3tSn0vRmHj
zYZNC7iRNkNAb++mxUCgqQaD3K25E9U9e58hl9Xwc4SEE2nxtBTUTDcmPfgdIuub
5uEG887GCyuGvWlB+7EwpfYPDxuoL3hwQYLIG5IfgjGnMrrkdzCMxXmQ2cTNc2bW
2zsOmZ5cMzl58eoQMZIhBA3POMbPSsNySe/FCuFaM8eMqylLjXEOnLUPYNk7bRCu
165R9XaZgvvJmf3aLARgExM5FOVTOLlEQt4CZiFC55MpefalJGlAzAKJrwfGWus2
9HHDH7YJyMKM5BCo/sM7RYSAvAcItMiK1KU0FaGL8qeUE1g/89dYM2nwWDIE6ir+
1YIvB02cRJjHCWpABjdKEmQYrxV1867igh8nOkdfQfaGTFHlnjOqwHx6znm8j39U
JYHlZNO2UXxTPqzxBC7Vmp6bDPTikGjam5SU1k/vFuquogmgHOwWCDQXoj+WZWH3
6i5hspOMxkwnYQ/bCUVVSxbMnPeMCAVHSQdUhBPjaK5r0Nj8O7TcGZnJT0ZzKBTb
YLe0E21QFaUBnWKBlUrMhdIHA74qlc2dge5aYWyr9zzo49V/89v1ds093YYtH06+
OMj0lmlMAwZ+1Tvc/CRsLgW1n8E2koQQzT55Y11lxnp7xRo1lyxUqGzfoiSYtU9P
2eJcvQA5MHRz0f5V3UfPHyhL+o1nVFMNazjCD5cuIdWBH0hap7WHXGOr7cdFXGJ2
A8bSm7ifQmkeFgXnbfNX4YUk5YQ/a2Bjhwj03sDAiUvkQBSZ4g7Vz5PRnLJPjfgM
iTFTVtz+mAoUl1IP4sTcovrrn79i6qIQwKa+yTExE64+459ZzONDBMqdKQURPeeo
8cBD5iKxckAUBQVjrvCKJNXcZXWw2Bcmd/yHJPJfePa+jaA2ogiIjVblLepd0PDI
at/FKf7T3MGNb5ELtxBPdB159pMHi4qCbQHG6SpakuHumXWk+Op20todSiSl9grU
cZKdNYJ1LxNIgGlUpIqnrFVvogSTme4ikGwu17HCEY25bR24466CeQtvavhzJbxS
c2ylhkZqENtygR4fvoGWqBF0iiq4R/qziRYUpqeBgDAWNVgrLFJHWGwmhORKV5CQ
R/h4Rj6UmboZCDhH9VgIYsCS7CCIQPd54zG834oX+lALQ0dcvNbs+2ducqKW6TGw
ggiMCDxvYorEDkRVFa/dWDKWMg+8QZR4RfuItecEVBz9VVek6wNPVFaVS/ue+aiw
TGDF2CtAPDXl9jQGQqMml81d5cwHNDvsYkn3y4GorlVRrFSUb2uAMJnlp0uy+tQQ
FIGKqRqvY1JT7oubCswojomdoJDdR5vzOO+xlLKSRTkB/36Z9SGd51qmgv+vLLST
5pX6pI/WBy41Y1Fr9aR4MV55mQFAVsD1Zzql5CdQQOSZZ+eSmasCzsMhknmHX4Be
URVDb7QxDZKh5G36CfjdBjpMej3kPtEn6GSAo8dvazKc6xV7LmW1ZxTcO72ceJTB
O2sXVIhl4HB0FhM2FeGo3os/YpXymw7DPN7dR6Ur8saj39pMDyrIWI7NJ2MHboG0
TdutFYTSdWcMMx32bR/fKtftYqM9zfamlJU06ipIBVokrvrkd+EuVwoUF8893KNT
pycBRsLE7HXespzwUiB8rlTCPSK/vtCb6oW3MAiwtaQCqV4FmIvaaUzG544TyuFP
Uw4u2E3WASKnRjXt/ylSh5ecj6xbEUsCUCxCfI73xSAhYNkz16KPB8lQFH1c0ivA
oP7VfCzu1d/n5qBVpOAGk3U6Cgoqvb1dij+WlyQaEQgZRw6igTYDisSRNvcnKTkY
0qvPhBAePhmbwGzkG2vfwUThHezqhAKyIuJosDRXe0/ucIex1HcBzRyLD+phsRxR
/Wl8VTsn7vCwevn27l7Ha+ux+eQix/CTrKu+SKw6JnN+lrVMEidgm8F2hNoeZAgZ
0sZXV6vE+f5rKppxw1vMzDS1tAU9SgZHxGeqSOg6cbK9izEpo9/f8t7om2hrIaR8
O/xHZL+9/OmiMNftjwXspif3t9o8k6yhDxkdV7T8fOLSS3UN4NdqIZTx3176MG/J
ThqvWUZJC/pFu/xJmZ+pEJCSj9LAgUcCQqVNv/01CkYTGgA11zR3/s12bgmHaSY3
tL86YLASb8grHfOwqae2nGtlBFIDH7IsyTyVVXAjnqG8xFIwTj6JHw8+9gMQ2jtp
hbXpIuHbOWgthSR+dMOFmQquo8FauHB2eK42v7HxmGJ2JC+n8WhOMQcJFUoyvbQ2
7VSOw50uEPGMdTyBQXWi9fFjh370zAXLOz9bjyRP3PHUu/BLuex7FiK9Ponj/cOm
B7cnE5Z5PtDuHHR5SCvL1T4WGef2uF7k/hhWS3mZ5I+U3mDBdqQEiXwn8w5y/DNa
y1eXJ0B0S9T02WjGSIVS+YmYuciDf/Axj8UYcPTyo5CfY9qvu/CKAPz7Y1isW9cg
KdC8Lpi7VpkME8c8eBgmmLclSO6b/XKmmfgoQl6aR8J13zP9DRU7BUdE3TAFrYsR
L6j36dhw10ouflpU20CbgP5X0tSISfaqs6eDLQ6845TS75vzYuLc41boTKVG+pqy
Av/Qhps9riwe49DKGXU6NqGzguanbHDe+HQdtkaCXc9XBTVi3tVEG0ALeWyl2kCF
gNj1vHiiIipyapaSHxS6nYcxM8o4VHqt/Sxwjtmgv41mUKpsR0m9o+zL/jNUSmXz
E5rncUDI3vQXB2Zj5mNUpN5NsV9UHXfBZqj7z/DwiCtKMqwl97hRsYggzcsadJWO
/lAiDXNCIbiwRX85uy9uDyKQ60bUhhTWzaPHOmxbbLuhHdC7v6/MjHd3HbJUt3s7
BR/vaitrYY6VyUxzuaQXSkKpJ5Fqzb5vKK0z0DJc91zLHeuAfVnPBq57zcw1UG90
3n5JABQu+eMeb1oaKSw+Q2MPLthzkRHooVCPHULMvoIU00MnVcwI9x6v8z8UUqJS
3hCAJjbI8oYNOxpwQSP/Mdsfg7SyCZyKf25U0dT3fOWsjQ+mAc56mln1e0v8VSoY
+jk/klD7pFm6Jq9DQcL96cRbvlrzmwAFNOKQh8z71LaQw3vbOBnJoqq75yd5xAsK
Lxnz/Kyy5ZzQCNjRukhGEEu8M2BKlNIimsXB1/Iibq2OAcq7QAn62B6QaGjAJzaf
M8qobKyu9rHG2PoPXISJmFss/q7kofH1pXqy1gQ3Hq8GbnixjJTP9fXthtnXzV1y
27ZJSm/3bQ6sI75uyKmr1f5d5IKgi45Yb0eg0wp9vYuQ45oeI6rCmTU28LaNtxoT
Al3Ra66+FdXki3+CRTNCH/qzegoe2UvOhzJ/5ml9GxfKcnDjs9MOZKUVI5AIPkF9
HMHkKjUglL/99OaAB40mqxgCbGgWFPA59ssIfn63xTlYWbJ0vDiCO8Q8dhIvyY+6
nDGNuNHXJffLysiBkPNfCGWg7O50NiFQMYfi/LBPlzikbUUyXn4GDPMTrkg6tVsL
pqeLJFPkhM9vWdqDM5uxXsZxF8Rpc7Li6Lx93E5/Mkk3CMKdPit2m9tCK7PIUPsm
TG5pwEjxEhnyLEptWe6nntDZ4gA9iJIf3alsUIYpblTzZPW8RRtj4bQ1GjbOTjq3
gkljijFFJHqRIrXUIDVs9wq1U5uKbVcDH+SfvfysPZ1YAPpJfFJZYHZ3oi8gkcmX
5mRjbQrVQbQ67V8itBTLLYgnEaI7j/HPczajfyihsgTUa8D//8a6mEveYNDcQr6Z
dnKy7Wb0al+MdrVxIbSn7O4YBdiIqbZATlN+2zKC+iyJR9/MmQVt/2Qx7WpL3dvD
w6r+nI2p+6LXwtnybTPZyD/kPF64J9PSCnYxSonhkq+P0k8evxwTsHVukdLfEUcw
VpzSR8V7jPXk6GXifovnXIcfFlcLYWW8egAuKya+miR/mI3fkBa92vWBfVQrdKIZ
XzFmptKT1xNoNRyoDvhssPu4iPSSKHkoyzKTAFOOX0t4G+CGentjWse9VruyDCGf
UZjeQNyKVgIP9fU+wxFnjcNbxkCUvZrYiVYU6EkEA8BaZfXgIurbh1iGJBM154si
NOG+t9Y86iC64tdgPCGuVASfOhXEdXs1K/tFk88H6zDwYi3KlxsxB7knzvAIQxDI
eJaEJcZpSAFBNrGYMpTUERKmDVbyi5ggHcHo0AdDU4QTy8CYNfzLGqaxV0JxrtAg
+YMWwJ2amkh5B2i41xZyqHFLQPOmPAOby/whPkFFi+zomK8XuzJqRVQNhTVKYQ7k
AtwOSWa3yI1J21m6iMAij8sHqj2IhTXopkLpB441P0zPow3x3CU96J2lvNUQOzCh
aYgsc8BxlhNOyAgBiHgxpSz/FvMy+h4z9JTCEJyF3DJ8J/rB4ZNSulI4+I5ZXF27
bXMd7yjCHCxvE8m2YbXdyR+/4rNW66T2V90pm6bKl4SmVJlxBr1mzwHiae6llO9N
9TNId5xTAb7uPG2QVBHKU09TjSroGGkJKq0NF94oiKnRzJVpfPdY7iEJhambo/3t
UG6TuhcxPRtM3e2R4MUpgdy+nnsXjgJFIWfBdoUy1x6KhdZX8eFZ2WnNtdyIMUji
Y9RhzV5tprfbIkTrJdnR5+v6R5RBKsP+E/h0vJ7zB/VFlEbbn2otN+jMmrT3IIcp
b70k67PuXl9OQvyA1QioArk3YJuPrdsNtj4aLgJZgtg1lEV6imsMhaL9pPi2vxln
DOXHF/QmKvWQSABC5hk9sy+JoP8d7CGIjaW9bAWQpkNCjK2eJ+W36KWPAakofsQM
+ppi4bI5gB+12w6QJ3/2kROQHiL1Nh/EaTq/IkK8DGXSDtIrsT+QKGXWjnLzDkZQ
5mMtptLtWuAeITxXksHqRcSmCCUgei0k/LYIqg8jg0oA8VEUUkn34y/PtRmeP3ZN
TMH9scvXLhq9G1MgBInKLu+5rFDBc+5srvH+unEBjhssD7Jb1IyJAlvxPqrJ5MIA
FQaaCcU237caj5FnnWy5ptl0R3I7WL0eXVAoJayPgc1Ezj3A9Eh1n1uPvBkqo9hr
LzELBJase/kwiRmClWvsdtFSLsY+g6MO1TQyuY3HLiP60msMlKqtkXLvRSvawzE6
fQzk7LlXACo/Mum3yaB95o5K1Plm52fNncQAEjvlb7DNJyVNN7UZ4SByvW8CTOYw
wrhZ8V4/NGpH6u5LyTY/j72joF2fuWkwNAZCI/9gbXAwSUWU9SMF+WQ4aWi8sc81
Wn53anxLkS1h1EhixLJcUXV8BWwBpQ+8oougnpqp7Kp/4d2RP20G8RGKfJ3ZsXpr
B415h7bFDdMx93zYGgMzFfWI8wAJYlarMsGA4Z/njhy7/A6nPfsEDzzq5dkyWGDq
Db7x5xOZuJt+YvYG0X4KiP0SPiAdH8yH0N8B4GmNdXGXQqk0HZ9HmXvX+D/br6br
RNz5Leed07nxIxu671nO9C05fULQuFyU9W3w0wLBnKpiysLNVeVEcO4kufog9koZ
1IP5rOUK+Ig9qQRjqti/TqYKTp2Hz4Q7wm//31+iIJVqCbr6w8yCk+rBr4o5LeVe
xYuqj5wireyqvRWvvtEI4Pv/K8LDHJDrJtrguq2/zgZ6yFMM+Hvt3TT+03/rXDWv
ut2aDM/Nyqy4lbYLuAE2WelZaSY/BTRTumCAIYVTBevSKH1r+EgELeexW9uiut6/
+uCHXbv6Hoa+PItwWGapQqvrM3gIGkrPG1oVa8EcgEmTPHzwLvj2Jpo8pft9jckn
GNCILy2fPG7/oQL5PlBPjH04A2HzTrsXX2kY3isGrNOJv1QBMaeQ80skJb4T6uaa
fZ237D4m3/WFrgzy6B3ExgqUZwMupgh263qQhlMr0noaQaX3zl8zKulFmoeUZuco
0gP2XOphZxGMZc/XEIyhlMwgKImUCLZcdHAJsQtvWwH5zz2I3vmixlhr9wS7DjIW
0C1pv79XlxOsRrfJk1gyCorJuEMeQEBC1LJxizNxRF5SS/qYu/wJjgWz/cP6+Z5B
0P3myywv509K893LFYJ+PfsyYgedQw21lwHr88oqZPsz5cececqYsxwzlbRbSJQp
08A1fZ+RwJKOeeYVra+MBhpJW9Ijb/Cvk7rv5afYDP9z4+EFX2XIDldCadT4NloF
mt/ZB+tKImf/BTNknzLWOYmR5aRrk4xRXt2SVpUv8vf9lFUphK87yN5SXRdDXfIk
Q7fC59ANi36XVqAYLHDGRRVfIBPffbHmj9LtNVyVfoCyPntSObr6IFxzojgGxUdX
MTtxb3MHaBNohpUOyIvXiFj1o0Pzn2jGErFdvjDFpI+Rp8Ij3cEiLYgWJmTydjHU
vEJeCuJCQuMBMoWz3uJL96CMdyQavOrwWPvsXSQZ4SefNxCQ1EvPoRHZLR1XY2TU
FxfOTWy8dhHmsU+0NyLXEO6YtT3mzRYFIyhh7dqUyTox8wvp4chnqBQbKVACdE4Q
g71Pz5KYncM+JfmNdqm4XA3EIu+SctjbD5uywJgsHI03Fr7DE+x6AWCuRGel9hrx
LA2SYp7HJ6lZmeGh4+o+pVcLrZ38az3uiyJ0uoVptjnW6D4lAfiCjvyHdMe10l5k
OGcPZUpyFccqFegZkdrzJg4q4CMG2wVP7DuQLOFnBzlkiVwLnpnHVSPk+xePHcPE
Qd5f96vMVWh7LK8Fwld3ImSHOp5kXk5CjAlAQF2Tygcww3Xa17tJ/VtccSq3dClE
5YjEpybLfgYSbbI7iZCyY0qDrn50FxiZN7ogw74QsqewzsW20LQ/WlZhUKASTbC4
VLDpwrJNkFFP79z7whY1e2p5AD2J9djlytfSJe2NctGmZmNn0nxnqgoGB1cuM4V0
cu2ztHBfKsy7se7vVloC1AyPp/01M8aNAL2CbFBGutGUadCCF3Ey751I9HkOV1vY
ygAGCC8LFe+Q9KBjOA9NDkS74W3b7O6z2uvYsYXFRIijVon8fvJDqotYlCR5ajRJ
KbKhI0iDB7gvn0lvOmFkAQX6DCCGkSQn5iBBgJSyKXaxLwUk0Ru/M1OOR0cEFNZ6
CoqCK4WmKoxcEb7z1FFjOx6ip0BBSLLVLCjwPi9XtxOe2ZxddEtXRiWy+BoE3sp3
U53qtZNSG76M0wdW3iANAtQ4EtiG4fXbUX9fgA2hn5iU1tiv/w2m0thiGw9YDQkb
CbmhRkbLtYrJF712Y0EjaTcLueUYZ4SxN6D2bWx5lvkbuFoDVJGgeh/SqWEvlDYg
qMux2JuLhMupHrZe1GRJD+7OeXWhw4vuKO4NDsEjwhdB/0nn+uGqxrPGnJkaxa05
LQ6rBsvXbnj+IC8pl/AF/K+SjfJUoJrJxJF3zsi74dPCizjSHna2/JhLWgNoWreQ
B1p1Zj252+Fo7j3BUHoQJkwoKy+At9bB+YjSpVe0l20keoI3sQ8UlneZCEqkioPm
G/BjC7C3dJTkd9OjTxoerVW5ya5VkkWix09PTc1NSeAlFaAOv/hzyuwPeEelNoic
/uqa2MaMV/gYxJRAzt7L3l3YAWGk212hz0UMmlt+gYEwZsWTzb/Ch+Z/nr6zPh0J
UNW6Ou+laSxIODTX1e0PlJvqKPx4KtNW/1j/kHlTY9zln8UOeA/9gjw7kiJ0amvZ
N5iluhpDK1TAJ6yzEfzpksRgpugR6mGelo7fSYAgllinOUV9xev3ubdwjv5p9frM
29tDbMiHfcVJT5VD90302QMllaGnxGQc2DjEJudIlkiNA7hcDEQeDn/byeDp+tQG
PYI3mM0fH/0Y3GYbmDQq4Vco4IfJ4P4457mx7E1uiv6p4E4xuHGmkshnbqIXrUnb
OH55+pFrCevzwz9ZUN+6o8TWuC/9K6+/ZZVe4fDDSnJWI0rr3fVQ4MPHthkPTfat
r77wi65PkgFNuf7qPLVGhVXsjv1hJ2Yh1+q2URp//YQFTfmsyCV5TFNl2YDXaS8w
zzbXoAu8KQkZ4VfuUOtp+gvNuUDbhy0Avw073Lsvs41krd5sRkaLojXRdBf3ZZlk
fucwjcHtfnqaxmXL5tc8nWgqKzUYub8mx9D30RxxUFveCcpD0lH+WxuHHE0EUdPY
ICtI5Xj2KB0vk0v0i6TiO1fyn0014+YKD/W5jV4tNaKvge4JfkTYvDBKG4FewkZi
uTS3lt8+aJl7K/Ev1CIIiUIND+9Rf2oMCo0yyQsx5QcvMAQMfesbFAsgVBbLXS8K
Sv4PH9XnB3Pqba9mTR+mTgSEq9SqS4WIf37FGC1qG1hfBaU1qjpIgWF+GFBRp3Zu
CM3PTjOHSP35C+KamQG5ed2Eggf4dRc5lqU/tImn2FdYRVZGG1FVskDLKzGpHjl7
18rSw7Caok3+N+6Dogu3/fOY8KvhHG9GE1tcmfgxzeCweXu8dJ5TqyTXrer7SDiD
dZUWD+lpEPouuszLiLUqUesXZXwoHAfld+KjIkCJ8X0aopoOuo0NLLAGjcI5hqPH
nEmWtclt0+8OuIA2bfRWWO3ZhCG3DmoSZnn7X+ivNo7TQ7uFGmCMUY7PVe1wegr7
c2Kgd+KQkbuNhia/SoA3eUzFfXjhS4JOLiC1iLgLF2SV58iszhxbvzCgLtQoJ9PY
ZJQK04ishACybJFOrhMey627InFfn4FSrXGPJQOg0q46AYjlMvOl9oZ9NAAw0YfE
gH+FzftZ1qSOTmXzEGoj01MEFi6WKQRbVdXkD14yzonSgOuggZJZNJHvQdkdd5bC
rUQ4NMyTl2IjhkTGRlbPUkSAMYlLzvNNc1Dn8KIZC7i/d4/k6j/Jc27Is2AflG46
Fa3AH0QwxBOFF/QaCZjCUEw9gp/b0hlOjnqWk5UrMvW4bV3EkJF0gL2R5YrCgnjc
qwVU1VsfklyuuD+W1LeB0Y6awnFEOf2EpthgZTlOm1Buo8BLgRryp8iV9XR9SXCs
A2jo5CNXdWxQtbI/ERywPbdy5nzYaH5QKbLijL4fZwHnSqUXX1mwUF21nT3oiAak
GZt6HisKjEVmv61Gs/ckEqnFcZjWJG7zJUQhi8OItc+bOaJPHItvQRzprWROR76q
o7JE9jOm75PINwAGND7xtoN/a100rZOSuyWujxMQ41EpuBPuNL3w3P4dRVCQQnok
3MzHKHxZqaDyNieJE73mwqM6bu4gdXXgMxfPCmVayJuF2EBUbdivXI+ggfeC4to7
+OOpJblhL62CUuTE6rUxc7JT4UH8TWNWCkLHCpcof4fThqkA2CENCYr4vs5PmmeE
5zoPoynHJyelNnO/jr+7x3U0MSgqGZFX55IzgsdKz3UAmZvNyjGfsaaqt6fzovMd
S/N1cONHAkf31XTQkU1Mm+s66JP9MduKjf4uujinGNH55H+qlof+JZkT57SGgufb
HT+1Bc6TXn8BEoWc9DUP1TcI2TfO+Y+Py8Q6RrHXgxiWFQW8wjYwUocHuq63KVtk
9LZ8tQVxphQb8/npMEZlienw9ZUXwuPzpgXAEvwmiw0RtRUgBvLmcMCP1q0YOJBL
K2mw0hqLm2KwewxVr5wWAK7XH1SHDueULWEn0qJaKofWMT3RfUVTQ8cqK6TTFWnW
Ou6hcn+G5xogZr3dD2kV03uSSTNxahF4cDQArf24xaZYkvSNLzVuSar7ySRpWDIH
lz7vAJgw99p4ZE+5NCP7U0ijLiR69lFnMUa/SuYkEsVnEb1wcovA+TgkmA+lTmz2
u97BTwOfhM1vS9IkGkj33eByubDHRW4uF0XKYSjcnEtd9dK1ch/FByZXx0+BITum
urDT56s/A4MWQfoaTv0GfYgvQ2qZS14ImGIKtVRbWMANbbxLBzxCMzjUvWquSt5p
G+0ZXQbIHIXEtAgYYbNJEC+k96kpRzTzXxj0b3gmpxCNxY5/0D2wzFpmAYHWaAWI
8LF/hUVWUxIS52meHYZ/Aa1D2xCIPyGgWPWiFvC+Mx+SSO529YTK1B5BCsXv4Aze
A0H33rQw+KB7OoPW/FwCwQW8R2/KG6bPTVj0o/TIVeMJIDmhQk7DzaBBB1oR/r8u
tOuJTIORvWq0oxH2QONjYSfwWR5C44T/gVik+hHacagxSWkf5l6C3SrI5tsdCdCN
Uec2JBXetsY+T+F4JZqlQmK6L8g/eMtXxsJ6fZaP78gnJQQ+/v5k8ldQyNYdY2zj
IsdVVghqEebn/2fHfhbRgmh/nWB+TCKY6edILkCijwN68dTPi86p2j6F6qjUF2k7
17vZ7BUSZqy3yrqCDd3G+R2XdvfP/lQgIHt+zSx79jN0AnzdLisekivG9gfa+qJn
/LB8H9FPdesDAXMFsqxwCPK0ys+bNEUy9W+A6OTLZwfkPqzUhsyPxjJYZVZeavn5
5RVBe9K3Nk3o7nISKPN48MFVAAQqUWrnAjIvUSpEqxr7lyUcCn0yGo3ToamZnTP6
NQQcG/EovFKrSO1ImqJE/NiD/sUZhyLpx2ngYS5TiB6Mm1KRNCcG3CWDr1kg5Won
9Cy3Y6sChoIDMTVqzEqpU+s+TC7ds685vaI5nwRm1CWVasK+P/DpYRLlDMZEH5ZO
3ubxyMShhEHVNEK9T5aHZEJEY4ndZ+7PCrfCJwgaGWdEf9xnhb+b80/iJCpOlB5F
3MEFHZBIQohTg25gRAddajV07q+qc+pPyp8val6HYHrXlArlVNRm1RQjY8VtUAzi
g8B6In0YI2e2Q55p7oHQqN+A1lDyDrLPOWOrl9/Z2Jk+DkM1JFibEh6CEUMCVuGZ
/C1jLrHJv2trlhD47R4kYLFnuyOy6MPUaSXvXhrk4A8PQpq/p6+CDQ13ZJaFjZh/
FINwckIfT0bHdXV79gSMOVf/ytkuwwBAJ3LMTLCiQQZ0cdXY8gXzkDBT+h+FEq8p
ihgv2A/uFQ/jDPgdlAXeQ8ieDZakCXaAtE4pB2KV4Muq0TSx66a25hdF6e51/drP
gMeII3NytlvtKi3gRPuW8NgCX5JDzJrrnyJHQrQL5lXLr0/6PiW+9bswlmJcCvhF
Qr7fLIOrscNLozP81Y9gqusggAfVW74/kNEka4Fa26W/6zqoY4Zd0A3FeIuL6Zht
iQI6O6isEBoOdPou49MLhWlNIAm5bTJ+/DDz2g+MxflPrXc6+EJ3l65KZNPq/G8z
b4xlIeGzLBzbbE/3NJvpNPA2Tcb6zfrw8wJ4Z2+yYuDt2RuS84pgQfluncsBsEje
pIldYWaMLI4Sv4f9ln93/kHpGO0YdCKTDNrSCTAXWvWCg4jw2RHcsx4RrhNVj4Nk
s7Dc8/cpHNbmcM84yvHAC7iKBuShU6Iv0WCHqHoJF5vgnCXxY06AZ5UjXQckI1jY
AEMsc82DpZaLTXVtkL97knzCYUS0LtucB+0oX+x6BpuUgATX9K5frk0vozeVboLe
/3n1ZnAnPWwKmNzf+ypoFRwWnTulaZGj0p/P0N2rIggTk4WcRDFYbHwMrA1QoxeO
YL3HEIMyGHyaEYa7bPwwJ0XBcNjZF2HzeRtUtHAEQ/pNwu4HLURh5sUaUhx7e2nN
AL9nkFhtUJafhtAKbuZ5hwAu8YJ2zzN0lwbx+eHFq0C823sPKnNI2x24zidsOsaE
gE0A6zYmmrmEa+/Jwmu3cx60izl040Cao0UkD+H4MTGCHSk4Qagfeza+NM1HKYlW
wofXWr/nsk9O5oXVgi3tY+V6JEhejVgUHAGPR1XNzM41jJUI163LMAfeIteUJhDv
WOPgNlXneBzlJzqUhLC8aodurY3JdCo4JpHs6mp21OvVsoCTDh7Oi+T8ZBgELSvV
bmXF/IIsrgTq8aEvfTxKASR+1+n66y7/lZ6hZqt1kG1weTwGVa07ikRCM+jgVs7A
lwEg5/oNqk7HiaK+gS76rVVqhsV6MKHi+Mtkoiva85Mppj4vCzon+CfCBPzrb6VC
+TBp646PhYaxBym1l8EeVRC1RVYTcXCr6UIJsBucv0KeKZ+QjEoCDq7cmtzvnI+g
baoNZUsEujotk91w7iDPJjuw5MFcfwFuUvDRXzNBMezJwmNeXxonl6I4nwZQVv33
oR31/FEaZe8M8/TxBqIVJjm8+apol+0eHKYAFAMqYhwcz+aS+v7eXVXFQtmxca9G
pRcdyur4ELo/uN/SG5CIu0E2rX/ZXGYF7p2omUxQnnVNPcKM0b/gylJM1C6j8bCj
D7TKO44PNJ+a7WTymH7RwASUJZ4fpytf2D+B4RYY3UsewEQh78aZnXN13sBuSRIJ
k4Yt7B4vBLhJ0kh+PHsQumjD3JUMbHOg3vbtaPev4UcE/TvNzDeHKdL4JEIjFkku
5b7EaCDIlMvNZrR9oOW3PDN4vvPYOr1rq6QdNbMf5CLt2WlrQPS7hazE/0SfF3b7
o29n4ZGA6riKy28qS+vE+28Z+u7NRCakOBdPDTCdSh8nSgoUPxRrdnI2A994X6Qr
vdhwUTZX89caHpn/j+2y4dVfMIUWRx06I6fFN3VSzcpvKQrDIoYoDB52+iIbCyxB
ZMtvVTNYpwgqfq00qzseMJhhS0eiBtYm+3gfr6LeLiRGeJiSLrvkm+JVUUJnb9kF
98KpQP3qL8/0NokstuZHo305o+yuouR4DBh/1Zkct83Jcw6D6hQC1lBHo06SoLC7
r2n+YZOx/NLNebk+Xd04LnteaQwixqZX6hBeqaHk/SgPvquJ5sxtdmEbqVGURQJt
36CBYQ3Ruc3A72MNAtiSQQyeEs+fEVMHxExM48WxDA4STudeEj0FUho4ir4+ongr
t34E9suA62SQ+cwXAnk5gZSXYBvCuSCS2POllksCJTUyHyZlye1gTfJvHk6tDLfm
qyqDA60PygHvYJ651CgngvXZ4lwTbfjyOVQYrdZejNbZyExqQxetozfgjNWxnQA6
A7V4LQ69i3+MyTCTCyrBL8Sjd9IErfATdWvhacvpmOFSGWduT+sxccEOINWrOuI0
Svz6iJVNDdMJ+LVOL1MpcUZCn9vmy3yxiWtMqJIX5OXW8ykAz4QnSaYyY+JgMUlu
kUj9Rx0y/Rua2TPL6EEJ48Nk/I4ocI2DUelyrCYsmOpMO3YKgs3ng8yStI6xpl5Q
BaZkhpb0V1i5An/sVv+Bt8WlHepB6A+qxqCc8vaIqG7i97esLShY0yjcFNmo2w8y
zZ1x1kgsWzLp5dG4bk9IV3nfIp0L2vCgx2Y86gjiEKwLeiKU3jnUV01qhIH45Cdv
QWhqtmxmLXUrEgooalWbTPCgERxlWgpyWDizolj0kaLErL2J8vzs+VAygpOAGLO9
neYevXgWERQVMnHUsDAqxAE3S9aCUex0rK87z7sWcSKb+rYr+hRK8014iMmEO8LD
EP68gUiZUCVyESGYouQBeun/0lASezEzeswLSHiMXY6/toDnkoXGWJa0E6Gt7BPF
tnR7QSIRA3OAKNw1YhRJV6f4ypJ87JZRXkyxOXZJyDBBeTADR5JloQ1wC7PIT4Je
I7YwTC9xOB+EjVvbdVwdcyjuyOigjntnb9mDVO5lsVIhNLidb4TrpdCLn3v8xgXt
4ncDaJHKQGVyTQZz21ANXvyPD9+fTLKI85qEZAvxHcf0ffJ/OUhFo1qcNeUMDxAU
IO7FVjDkkU8iOtnzB1GcwSBaJbt7s234Z+W/zPRGHRPHw5LJWqdSPQdcF5yr5Y9B
70sJZj3+4NddgAVs0HqhWQ8HFSc/DlKauaKEyU+/LKhF8b1FT7tQ9M7h4K+V8GHJ
CgtPjvM9OIBDCQJ+aQsU9VKq7h+A1AFNt6Luwbk+F2CvCUaQLvlDhhRR2n4pJeoF
e+JUabA0u9cAQ8TdjMP9j1j3EwNFVhmz/eRKoqUXj8uXAuFP4kCoSNoKn2etoX5r
GT9L78jyqJ6PZyNonTCMHi4ul8dSbFPhi5btqVXotktzGaDBXs5rq3/+ouBL/WA/
HD93VrL+C/natgykVI2NQsD3BlkFaCQ6aR+s5Fn+jAx4LnMH+km2z7tD9eEI5ARX
iGPtGRNphaDLiYV6VXiXoAJRRlIiY9AewQ9DbN6U48iC1G8tYxRK75bPBPYNN7xD
B7UJ8vv/DLDFidBg8aExnrH60w+SIFRZW78bca1hX3k+KoE4sQJb4hrVYEdUvybq
NYtHZj6XTHvnmqL5WmxuYAFl2ZrvtRoFXuU5oSMQ09ar6cfH7mWio7i+R7Yx1WoL
2bE3HftW4MKW7pFXov4vZfG+YpIibsyOVyYynLVHt9OMNrp0GxfQk6VnYpki9MS9
BTNd2ogGCiBiB3zvgWD8+w0z8cBP7kgntxVczCZVzECJJWZds2HWTrPkUvLtlF6A
YDcmh+140HIN0vuj7dGP4twPp3E8z0KmOZQ6hwYh/8f2YjYV4lj9ApOKyMrtxKTN
egXMMDpXhJN8JTSx1dejA5GZnKchXlAZSb6k2EMuFFJuB3tZSX2gB7Y1g6gufCfZ
zXzuwLhSugPay2imsrcLsx09ktN4SSBVVYla3mgKohuXp1e3c8I5M3b6NZdolblx
oi5m4DkxxM5UmsQvFw8XFPabTCObY7tc1I9Xq0c3VGFEY/+ekDFNNuXRVNWpi4JK
cPkdhEmpMT6b9fB3EjTgalVCaztqo+2qBDbdkBd4llmamYQQWysyzACQfGlpQ1LG
VVPXF/V5lPAbEW4itPD3QsltMuM3xnbOCDi7nzYBaSdTusO4kku+1SCI6WdL5mfL
xJuNEYH07Nka1wQa+ud5vDN/Dk1qrblfuO9PK7U90TtUGQTi4maYC9aJCHH2+TJU
JfxOHJ4Ue6WVUxbm1IxWxiyokahaN0gyNlzoh+EIBY4h1aTebo+G9X7PS/PvHvBh
Jn7EBLZccUGSu/cBhtKncZoxcNCbWQHBvBSFOzJae7L4QqRLhZCh85TVwrrCzneX
n39ip2YqG4h5HRQ85lag6QoVM1t9mJXsNJzN0gjPcGAMjmMiAEPxcHu8x/sQUDkJ
ioC3PF69206o0bpso1WMtpi8Gcn0FMGIupyxP+ToM3bwfri9Iq9/AndtstgbNOsW
3t3bOArNlOJG9l6rjRurqHoErRm38ziqyFqXA3045E5d9rqS9gDOcOrs2Bc4wwjC
txN7smHewIppjJ92r+fPSTGfcz7WRIYVal5JC7IHpeA43LtDMHg/aW9LCm4C+uTc
2osmy71eL3bBo83lNxE5gof+p2QiT6BgxuNx5vajY67z27XUy1AD48PxL75Xnvmp
t5honGXE+Hl49gcXovDG4W/KSJqSuYkE8Cx3fZ8NeB8Ji1n/2cyCCu1lmgVeBw6b
Yhfw/0syKwp6nUIr3+R3+3eTPZw3smTNCDf/2Su2wqMWFkha0upfkgpZtwZx5Jkr
bKq6cv2w9VP3EH9N0O4SAfHRkqCA+xzKP84yFXPLsWtbF1oQ+IfBFGaZQMLq9q9P
5e0hzxmlBkWSMBMweKIzj0rzBAfhUdSX6V3LDUvA0v8vtHPUkWTCJECG2npSVIfS
a3pxL9vlYOmfxMjZEXvp0egoBwvGfFFZb3/dXa3qQBY8XOSjjSv3p5OwVvLv+Wjk
gm8lT9bppaoDU5Vqnp+IXka5YMrzsSo96S8uF/YWNVwpggDm41py5s4zZj04qWR2
8kiqvSFTWT5NGbAo26Uh0PCWalU4NBtgxfC1VrX7VuEmwCOJLzOv1wOtuatVjYY+
vPieABivLIsRoNKgrVEkl2vQ4ofbDLYdwRDmmClHXnq9PyrA+ebUMA2WgxWjt38B
4gVPWWgh05hVV2NC5itsRxY5+rFQd695cnzPZINXdk7DDLCuyheSiFBFNa94j+aS
5/SomH+BX9b1ccJDmdk2P4RTRRdrrTLFs0cNO3/SeN6n7sxuNEpF+PmoDclxzLit
P3zwEH5NzEOcK6ICpTe6alUwTvw4lI281H+kV6YHwa+/w/hy/mqm582PbRp2WtWq
GMkEacSqSlfxUg6ZZ2rEw+tN0joHdvSm+L6YbPMaojNgMx0RKyr15VS7FWQsIQqP
qGyy5NxkCs5Dk4wR/JUaqBKP622mWWnSRXmpGPo8FDqduxttCGy2vT3a6J22cJip
mZxbebr3pzZg0PtnR7u/YvWGlUwncWA4dGRZc+okwF7uz/XYqJDgoEBOKPE3BRBD
gnk4HTPT6f7Oj3WU8tV1JAL2RQiM7a5ijrWNMfdUulCu13s59tttfmgvZ1jfI8qr
ebIF1/Z9zgAUYnBDjYs5cX7ZGQ2lJWFkbOugrFn9E9Sz8W0DevY4fQNwz9Wu5yPj
N/t6x3c4ORm8LIq8XmrXhaRk68viG2ySf4IiDaaYFfbRkIGZZO5H9ZEk/QmrDMLk
RWd+YHEraV6OIEnni6pn5spTXhxp3yOguQK1tcorVaI6VrEfEPq9VEo55dPbkYf8
drRdxYIuaq5wZZyw7AAoAzsoTnSU02urIAjkLFbpn5hAlyHR+/Cd8jZE6bjFES+X
8JFoQ0wLsK6pqYtYEiCWXwzj30SDE6RkPICcOdksKS3KRFrTFoELHj9RFO0husB6
rZdXatN6KGMDUHTorv21vt4CVo/YPT1hfx5UOOCvZhsV3Y3hUCFupCB9f9GSCcOZ
ZdonvLIXTBbSid41vaSzgKTtRpP538wKLsFA7CyhSi4Y37iANvz7jtPxSmj/8xJx
f4yDcp4KGekrg2zbse/jcCXpYKy1VuUDsOpuDAFzWQEYlc8/+Nuajy4IOa2i/QMD
rFiltJaTlzf74z0xnxv1mgH8OnUXN6ImIdhFZN5OsblWcntbZRsQBUQ8JvMufrw6
Av6qYdDzURz2T7lSaFoUz9ZbDGTg29Hbwvyd9dwiKGuVt6JyzkF6kepyBGohjGQi
0tjqMJ21VtWEXk5ltenu8QU0uq6NKJiPr5YkC/oR9NIeOSH+F7mC7poi1WjoEMvg
dyKHnolBsdr0Qthzc8bCowDynmKBTfkmScsecUgGbtkuuDiWiJ2Lt0WCjMEoOhWH
6BxewSK/HCCsuOckPdIT2xpWuQ9k0DH1qWoRuLgG9Vl6eKpUaAJdNd1Rjz4id9Oz
mdU0kmHBpAwY7P6imoRhVorrNIcGGWGugw2jI30ZYpHDKGF0j5/xX9ac4gtI+J+/
w/Ils+Be5zFhfKCHdoMXcRMpTCSnOUhy1YUXG2maG1+JBrJwAqN2AF0ETq/NupaU
0li3NYMoowqjFQh5ZZMqtqo+3+iOMkoxXIaLqCFPyoEpDV9wFq0OLwgpa4ASwuJY
JoENZvPSV4BDTe9jSY29xlSL2UJseq+axtGc87Tt9n/7QJn0J+/nW/hrMtYr1pun
06mEARb8XYMCkPmq1uT2FJhNDtlV1y1y+09Q6UrFiSYiTMNVTAsmZWU+3Wq4PB+K
SQiDZG1rnI4STFZ4xljHQyZjAvm8L3OCapk9OdHKbQPe+i8pHiKDbXvWApVOZDKh
74wj3BX8jVIbXI/sqYpqPYthrrU3a7E3N4QHOQqfuyfHcH/6jUcXq4tgj1BVAXMs
LVWyxJ7QUBltxIlYpYMsVVhUw5TF7GE1EvgB0fwrtcfPseDsihz1rUJGUPu8aWUP
SqaV2DjdJW3pNIdRzgSBlEWIZmolkHSZOmTcYZuprePmQ5rwyDKBORPJKIv67am6
F1O5nMmoUtPygN8xoyvPtMtOSQvhOug64E2fZV6tIp5LGveD2bnF00dENGs0c8F6
w+UfuuDZrFckpsWa+S9W9dVq9jUAdCsj6CoXw8PtNSk9Yi4K8bJ7KjsSkGGIJV6S
aCO5T7MlnayjhQPbXszsPCpWpLVRwK48G7NXf6I7mSzzFdM4ZW+L+0uK8EEcwBZV
NSFZyhVWX1Su6AlXjZyGVtCEg5WePsqvOlBNwnaEttLz6+cPJ5tCmGNznw2YS7mK
l6PiPeqg7MgW6jcSMfK4e8WIrmTDbRymWSFPLc8P+NVauN/ykIUB3ULGd9Fu88XI
bFFdIX66pObQkRQTXw8ncgV+PCUlIk+iW9ri+MtZ6FUaMMf5IeMd4BZg1wc6fbRK
N89cHEXQWdQN48tD4pjkozZXmykKksRrZLTe0xMjGlCNjATaVc/k/9JAkD4soDZn
i86wwY+0szvgiD22iu2fxlfErlZ/6doa0XmBzRQ5hAL0P+tP2j/57lWXp/l5hgzY
/UZ+dD/bMJHlqhoqUmYVOfx3LvL4bXPift/G16J34Ch5OCwRiXFpFTlLqUURSKC5
Rm9HghCXbgXYkCuM6oyqpiR2V3QhXix55S+fAkQY30AiQ2JhQ9T/fXLk/rKtOBDX
XCOgIrGD/xjfxffRqGSVqoOBWsiKSuDP4DiStqrflHwVlSRZdmSO94IrQXBirOXh
UO1PZHso8NnigAqdy61begN/QmyDqhyKJ8Kzamqubfh6wiBw3rS9d8Dx3WMaGuQO
jVblRl+vpfCgwLz8WMITOJEHNNHdbG0cX0gLBYDYz2dj9E0bZAJPIoTDMxOJhQ4T
fbuzBPx0ZLG+GZHJOg2E6GAf7tTAY8WV1b7NCKCqSgMGQDjs34ALiikAnKufbf/e
hLK+zK8gXyZ/6K6bQB48+BCfWc9AXPVfi1FOzbquFrkmhTuhTVlEw2bXdF2kTWY5
PU9lcH6dMRs9bSw7Kjg1d6MtMNzu5SFFB3iQ0q/RVtAPNiX5/B6Yk0x85Q/qbYfU
qGAhBpg2L4fYvTeplSEHDB+4P4wXUWsjXndldHMuwbbDhqHjTVGDbxsDLt9t4xTL
yjR5MmF/zA56fnKQRTRvhKBSM8c7fdst/R7gt/H8mJ3/DIFcdzf28wIcbT0nmB81
tBNSeSTIivQVGhADjk8YLgoGCzTlU2B7zHCez27ryoYigoAKSpYO1QuUyboUp+wm
y6+0SYe2Pj5QefNEbVMPNLgS1jCPGBfD79e77jAsY1ARCTyVzB9zE3W4ihXArZME
UiipUKBwKvMGcuNZLJZ6MPiPVe5jO8DjaZ7SVx6feVxvj7vCzCIgaQWrvULcGUTo
7b3aGPHtzRgVSeJGVmL40BC6xuXFRfvDOkdsO/GW3cpLZDC8EdwGXFA/s9D8PHTs
i4eOGuCoOU/iyepwjblgGK1dvdov3HIldiOsFXZWfY4scA1oGDDWLRhY6aBe075h
yEQ0VZGsWxRn0B4Ddt/V2bLKqJiUYd5d8IG+/fXFeATlgjfLVtlvzrHNbqEtaD7R
18AA6RvQlpNvID7uoJe9grR5S9YEi6PqsEOkGndj51cTOMYToM7PVzIWu06yvJs4
toPF65+PubRSFe5NiIlzc6OJbMz8VtSXwgZlcx+4mzDP2SN9+LM33iVQsewjXFuJ
LTU/RMyvSFWRj/E9a8djTTbVU+9f63XdQntU5KJ0EtWym9J3qS4n5/uD/Kx333vJ
3Wf49KfPICXiLFLlJ6Y3TyO2yHWBVxeLwLsP9SBgPnk5q+rWsrCkb9cR1P595zaN
pOKelLw8nRXqG5EIOM9poAEs65YwbOXxv8QSq9TNEmarHvUfYnkyYMd/1C1/ire+
KWah0Q+3BLcmBKBwL0XqDUENFNmwc31zBJX6uAa1PtfJ0OAOLOqfi1eDVWTe0N8R
jFUdaWrGXeCbNhbnLVkGokpCpQudh2Cdi0KnEJh0JdFlcfEqOvPt/ZQ79s0vsfPF
AL2FxrjaB5htgEm+tWHJ2zWNrTUXpQkFKFPdQ/rPW8IX49liMETzoZtNgVvg5h3u
szr0y8w68flSbSe6/kJZLKSjzrbnqMeGvMDWxRtKqrtC3c+BNvZxItxkF0SqrIYL
9F+gnPmF1Lb1ulXhWiddzHCTOMhLj9hPfIIDPILLWWV0wWAB3lt3dPiHMhTTah+1
Gc9HtrKgqFMfNRjvDLDFEEhPHq1oV6Dky1itehzSePDn0toB/LRKYsP6aiakY9PJ
mmVzE2ts7C02p5BRMwDJ5acta3ninNIMRI2XPBpDbjE+6kpEyQGDQSQgEKDsTLzQ
/RaxCyK0/nVLZYeXsjm2QABy/uQx8OUdYVZzZR7dGkm6mPUlXznB7+XY/yQwJbJJ
avIDRZPQFVsR5CaTuKy5Hh66MYqG2fz0ieKeEFXz1UexaD2z7D/x5X5aQEtllZmF
55QLhad0Pkg3Txtj/joGdclQre5IxdYd7cHQxBzSDSxGMeOiP6T87ewQat1yf/X3
67JDilzb7kheOU3tu+3I7IwEq84ydlrOQiL3+pkgEDYVFvTXXIXo+rglyMMDiThQ
hsosIZzlnkGH6UuFMblZkbEbtoS2/yqL4+GXKx1ebjLqAUHCc9MbjPuLPTsw0Ck1
04dCFcEBb6J/Enh6pLFZLGOMEvh1dqSxTPM40kJZIu0YDUbsuZsFc6qanGb28SSS
5U/ROuq9F/iwZb1d00D8ZzFVUKi9XFrz/SK6sbtV6HORGU+RcUT6DMBg3fgOR58g
l9hQUCBOyMUVNdr7h4BlKgqjnNXoMv9yDi5m19AQO94CQm+38kc7Se2OC1XrLqgx
uavH3DgmAheUDFA/fIkVcCXErqON5FwB58Mfqx457rxOCxig8RLRQDY8O7wmsk85
T2N6fDGv2I24wIKKtiH7H8/5PEAG5mx8YcWtdkwp7yL6OwHsv5b9xdoVeannYyUr
KOAzLGyyXExgRChPBX0X7svtMQ6gxXdTbKk2EcB9TNx9j74Kh5nMhJvHYfYwPbwF
Y38gFvXdk2/5zurVq8Aq/N0VIGdX9mPFHZ6t64sRWD5P+s/nObhsNiRODtVC8CXi
RinBXN5vHpE1rT6B33cGQBxqqcGJEUH+hVZm139B/n8kCEH2eGCjSNueQNB4PziB
YTVF+6ys0Od8Z/wP/rnEMKAC7a3mbBT8iE0VZC417h0UxhxV3DaaSsyrUDAoueNW
oIM2GC+w4MLDMNYhtlOYnMMPG98K2H31rk2b64xNsbVCjXqOA0stUfDH5rfBlSw9
90647kLZskhsHJLlJdXxlxFo23rlVJ7FiFflG5MBjNMBIEZEeY5C/tp5DDyqbFeM
b4iVeLXskP6gsVtyw4OEnIr1LxU6Zb3oFC1rMbXyRKgTa5HvArbFnZ7l0+RjAcNV
4KVwibcYZiqPVzaAvPDmmiq4s6hYZVjigB/6M8m0HC+IMz3dy6EbzVPmFd7ABZFD
Fql84CY3vyuYkfUulAOh2qqk//mt++hfdA/V7Q61rDtrzqjFaBwNnNJQi7zEQiHz
/o/qYW2VvVpn+86QpfJXqgqLZMZQy3F4nUkL5tAcUsWS8rAFxr53r6SXfHZbtGYN
tUlP/innyFwA8ayKU0xVrekgjhgp6SRlP5ccn84LoYxPEb8mGhiexKrJ1Zg9UGcK
ru6qWasxL/7shqpjLhbVjS1wI4mwOXUcYwuLYwoVXofQY9cVRyYnK02bjNBwjGNG
8+2DwgI+ojkzNCILWdWrhrTCrHz2at5xcJT/5OSreQPw6iZZ9Z0wyfUTerFBXaED
/oN5KIebGO9LsgGRh9BdEEDM8yJGlP0Bg5iBYk9jWbzG/cEgqH9jNjxu/Ot42MDm
ghY7Tl2JyRxjhuLQ4VvSysBsPk0l0qoEUKoMoF19XOXIPYsA1SU3mSFqJMiJFCSa
ewHLQchZ5bTa/ONLcI0msTKfJd8rGtYEuBSUAHM+dmPLGDM69k2PXtefYIHH8c1i
wjWIDVjRQtqQogg11WZ5wI6Q1nNDKpo0cd/PM7rBfzIfEBphdBId8V9089c1gYlJ
V+sJS8/0rqdS7ZsiLlfBrbNCnYPZgxf5yRlqJZIW2tb2Sq75Fj4IAHK3C43rWDxy
DgLT6X0or7mpnlmmqLAFiBMhg+t+uhjq0eXd0pCBjBaknuaJrWMk4uIVSp4M2h31
Edsbap+r6hrQhC+wfjoyZ60esX6hefslRLETJybUXBQsJpFyQ3aves9E3AtHvRbd
ktaRbcyG7NYjxHIHJS28+JBxR8R0DHuxD8w34QJWwVNIbzcDVSnxbWzBuOHc9wvc
YlV/4nUeeLHXWT4iRnyIAYqo7Sb5gUo3RNcRqVbrYAA4cWv9CjHYgoP/CPlUTRsx
jmF9mhTBgbjmHtApCmNvt30MRndGOXjzZjwsrEJ1hnfmHIi0g1ZThK0NSthZam/g
29WiWV/HsxlUMroAb6dAOrrU1bBr+kaFnegmOFLSESwm/SSyEHspWZpECwVchEGh
DRStp6pO+//uGWI8w9GSuj0bLDZft5g4yg9JtMbVjOEzCGmdV85cZf+Ns0IDyW/2
KTHz1hpAxjIDIOJ9pJgU5UfIu1TWaZnJFyqJnbvR+tmNHY+VkGU50+gRjIUb9Ad/
qNyCZUsRaWFCUiU7cAdNBtPyY7tpBdWy+5s0t5TmprTMnSsS9PwM7GVwbIkXmVIa
NECnyk/i+i6SCENWCWDIoDuFzFoC0y9VSKOy+H96+9yeIs/pLkkIkoURPggvciPC
H5z3a/2efytvKlxCU8/tTF+mTlc8oxg5ry+lEBHMhKeCATUUtoKien5TWsyY/rmx
NYhYiL2gocI1GL1qKYGe3//AEHn7m1zMUhY4dRdJc1lFsJMYPGLmuKoTaity+2Yg
ErU5Lql8kSip1T+bHtjxAoU47ynN/InxwH2gPxoqwcWTD6TSAJ2SLWTM7b0jLQe3
LVa7Q7b2vJq6VO115UY09PTTH/E+Wvox9KUcq2s3L54WAyD+enm/kbViy9dteWpy
P+qikbjhbFJtD3hK9/4+ypEa+bXSBJApPfFUdoa/YAOxTThDmTjg0TrT9cDbPVW+
GFMOT6NmnKj9wpY7j7g9K609C8lQemcaOYXJQ+FdcXyaW5Kc7UHLXPnyAHrE2rW2
+UwQZwLJ8eLJUo/JA0fpW8SaOMhrcDf6rflBKHHKOYj/LgqAYOCs5WkBgF0xzjmV
ZK2Ft33uLYz9XDr6+TbrcCe7r88Xics7s0DyzG7/hw5XU4/4VwupaZy9QIOWNtsU
1CulpXCaWBkGH2YZJuHdWu+xS7YDPSMtBVzpF9WX8J8bpXJcCJYzcZkKduErsbc5
+hdZ4t2UEW/feDV1Cv7ep3sEZfncnIyeH3v8/EagN7tI2UiLr+Qm4ILrvKaRSFeQ
Oqi05NqSIiWEZIaUcYOsYGCPD/gEKyrf9t4SCWujKzG+Y2mhjwOv7Xb756Tkrs4j
cN2YrSe4FaNlEuTpAEi1Pi1zJx0gr8WmCZcrMCyXqqs7ogX1zF8zssYYEMQrFlXH
rGY0G0/SQyNYVUhttWH1ilLBcvdRRmTDpOgRGByXd1M9ljE5QCdpSEooH2NsgdUD
C+y0JI+eCgo3qtcVswszWkvNmt9gyBso9jAlYHFfKHEmBwKt85Hu7RldVTGrl9xd
hfUXfztpugbFtVTLTLyAyEWCJqt5Efpm8Im3lWzWH69wW6q89kIxzwYmlAd8VfUn
eo+nxRHI/5JyfemoVzD06jH9FQniLTvrChyfINTsaMximmUwhEg8XmKVodEhtRJU
AcpOVtu2DgwQ0whNtHMrktWkHoEt22VtkjZ0TPYpzDgscU9Tm94gvV+04Ff0d048
TCI0QjPjalU/zcp0RmljqVKUgBgCqhBBslXkWQ/0LuyCf8VuENc49Qm4ZPvUUX39
KbKpLYrq1jFiji8P7n7upZ7elrhd//Nb/HmRKcxVaEMYVImgcCRcpaRtK6ptigXs
VvCO1w6VhLkQgJqS/b6uJZ2zRZaK3tlkaYdAN/14gIIJl82dL3yYBmfudRrWYFp+
cCfgX4qqhIF9SetLpmiFiPRh59PTAhZW2DL5YPw2pHTSokLV325ewVDyIssCl8XZ
Jz4XDwyWItpd4q5T4Hul0zbFrbN8U/v6TqmwAXS5RuUWBJ2vbVMuEfYI7RDXlaah
ego3ut9LaB1kxcuolW4LsYpNS0L0bzdrB5h7ilwN52PplhmdfW+RxggenADFnYrV
qrFnnwELhYnJbmD8XUKNibPwBaSE0WSborVFECfnbrFcfWyfJaOwD3jGuMdwaNB5
YWwMFGwTE+fX5MsVZRnO7mv51E5TWjJLBIzqwDW5Iut7coD1rvbdrhN7SlmP1BnY
ESocvl/fGXD+vFT0hmFH0P0SsjpMEjl20WZKHFiPfjtqHhgrs6lUTIacNv2VpjXH
e0k7p7YKl4fciad8sbxxHEFsRmZZ1qUB9LMmmyXJTiOpRt2ZFobVnT8dgTQGl5Nb
wJI0Fe93ie6/c9qa0BnYUaI/ng1x1efd1KwvqW1jenSIp4tKyp7eet61htg2YGBV
hc50KBR82Un3It4dYW6sc/NUUmQLolx93/RYqIY5ku75nnNuCc93QVSlFqcUaPuh
98AxgTNzOJHvl9TSPov/KErVvrM1XgF5Y2sdxDLVJvLnxzk3UqUXc3JDuPfnpemn
5wzuzkkdo1p7cZlobwFjAAnDF6suVYJxq0eRuPpHgRet5gCCiHfoiVBXCLyLcwVu
AnHEyB+IEOdfoag4Qhw9WdwAqqdi6v7u8KDwlj/S8SPcFRyWxg0eNBeWolBw8xsC
kl2vY7oqboUK29HO06qZVm9oG8KfulPnsL56awLB5t3sJn3wMxicjk67DVbIY/EX
1Ivd4dpU7FlTcB+celVnWP106I/CIc2ypoSQPA5zHDqUfVrP3UTV+E534Df0GKpR
zGcwhTyhAgJXBl/HSjXzz3+B1lN+evKl+N8zfsydk/SqJyCqJ4fS9zkEzP6ZPlaI
2qH/OvfRaP5+gYdywvagjE8bCbLuycZSl3LTbjGIZqiE0dHEk50wv89DyebC9h6a
VgPTfQ9MmYbao1WB6qd3GRcrSnN9Cm/Llm3+1BiIhtNnibpj92Kx+4K0zr4LOkFd
Pr7M4B2R7wffMcacCWDm77zcsAgwmDhyNWVUItC86rLgqK9G0tKrVpK2VBpHweON
hi7nmMIDMR4hIduoQGXKete9OCVJmmpmpiAc4fexmnBVkCvIGO3zYJ3F4VbXJTpu
tqDefgM+wGUtDdy2RvUnguvC8AHSF2Xhm0SlyqF6IRUlK/gz4Uu1yWvBFtAe/S6o
CNoq4LxaUPGHGNWeXin+F3poDl2jFoyuwgqcCAzxiddwVutVJV/+zB7EloUeQ0rK
bh8ruk+goZRGRq9Ox32ZPg0GO/mhqZts+Vi0mLxn57lsDT1WVLH9aGf3KILIIYW8
z0KTeyPUroE6M8hZ1sC5XKR3xPCRCrvvmw7S3eG8u9Ib2a5XArbecMc0EtfIMV2L
fprd6/MqT+JSYQSEg6yLNSwzJ+1FAE4Y8pEqy7z8ppuxPRv0wbYwGQJwjSUQajAM
Ej5eRoDDRrIHMLq2VrOAW/KaTECnQ1Ep94cVybu+xWcDe5TKxinicSsHw3guIjfO
w8Ez7r932jGwcro2NmJWwW15O8UUMZiR80smXNJ3ylOyd48Um5YFSlhrPu4gxhPK
i6Sce/fNvtX5Cla4dBuZDN7KGamRltedDnEq5l3am4+TwS3SWPWiD34Tj8CbQ5R4
pi1rHKYso5aN0aUW/QtyrzpQU6MXipx6Ug7cAZuowCoU3XjUL9i6+GccgTOqGAX+
muGVCsprz9/tg17rAmjb9jbuRC26uvFVlHGaEqmjDGbP8/MXtvYK0YiJfCzoVEgQ
mDMMCdsJ0YdW9KQveo3p3jt0jXn7U82cGjVPrPUrDKCiVkmFKeeSFaTE7tdVdlu/
sL5joACT78CkLRwn1eO/ijRy9XeSJ0p1N6h5HHu8b19fa2nC9r3rpG0I9KWqBxF7
TL5Js/mR35ljijEhwcge+gNL+mpxzzeIPO2IlOq2UQkkX3FrchHsTWUR0NT0jhja
16Qu7awwPQjcOxBRJrGEqmz4mHM1HmRw9vTfvM5THk02reAUJ8R7x6Sj0Tevp4u/
jz49P2syjRFAkqzCYua2qima57LFFQEB1Jf/DalFJTiIhrH6jlUkLbc/sKzD+WhL
DiPc5g7NBnaT9l1Schdqh3B0SUbeIYwRkyFZ6xfpgOLNF1luI/J+ef+2N/WraRc1
kjQFT3Pt2PYfQhnYVwk1nsJDSbTXSH620fV3v59wVV/9whmnjUjVXkWGsB9glC3T
1e+e+557mGOG0Vj7PFoCjN/g9bfDAS0ZLb5gJYKFY1Hy00m7Vfl5Y3P7P28TF84g
iadbhByD+plrjiJoQ6ginCuJOAaKdAB8jiVe5bKAvK94reKGr+OguuSR4sy0EAXx
JHrJ5sNahwDUHQ95mOCSflB9WJ0xUearVUMkI2NMs+gkqUyXUUtUU/zcVFngDOSY
LQ7dAFgQpefFhOrhBDL78ZGmW8JWx98N53wLhZz0VApq2GaI/cz85qK2NZMw1g9x
FYT7byr8Z8H+wUlEe7IABqjfWCYU725P2pUUybiAii5gswO/7usUJM82bjTenPAf
B2FYzqj3i6FZKxshCzs8YUs4oa1nbtGeYHNkbkoqcQbPodP5wMNqi+6PKjNj8q1e
hjsGJclJ1tBqGDCIvLE1NXgG6tv+9hS8dpvfkVXhct0MyP9Cxww6e1Pr4y8NNnRN
BSDq2oQXIglZIXSuvUZD0oATGhWUptE4z5toinEnaEA0nZEUM7WMbFjnNzhenkU2
sKVyu1QgJVcpl/6UtHEx+H9lF58MzVu0prUXrF981SK7QMs62j9hnn2clhjxXZ1g
f5kKcOal8VyS5PGcASOPsefM/x3bl2ECvdVpZx2+BptwnL80wyk0z8zw1H0mFx43
/1fSQ0v9nYZEO/llZ++yBAwOWmMrcZfqG8FpszctQuJTbMCmze0iE0pbbiQeGMBP
MYcXySw3bojJvqI/6nVpobfyRf20LtR55Gbxc+/YRgQYVvgpMNkg89A2+2x/OxTC
yB2U7s+rpuO8LxbXf6qiv8vJRryroeyeREx0H0fY9eWKgjwh0YgXvkPxscpYf0wM
HroXpInkfEEsMFapHHxCD3pMHvI7spsFrJFt5O/LOxklZE6dvGYxV/zi7UnUexqr
j/KrwUajSwvw71DiMGGNBJWoTKdEJ9qXTGwMEAsIt/0iJZvbpwOoWAx8n2WltrK5
JtrbzBQIAySMVCUz9/+e/GIXJ5UDzlyMZlgbJIYq2KrIrI0QARchMl3QVlhJstQ2
OdgToVJvQHR6S8Tepf3bUTbZ8gtOt5CCIVp/1wXordyT32G+aeDeAGoIoZkoCTfi
ma8NtqvQTVZmztLYqF4hqdPSlGbgWqL2ep8+cHCvZvATv3I7yr1Ao9vzdkZpO5Wh
b1P39OIKT/RRF8uBXyKkwmbKRENU1TOxZmazToPSNR6d7VnbtqYHWGZe8AuIoUc5
9biipyVVJRSID68Ej5FL1ANH4PwvXqtzgytzjO9DfgmLcApw5Lh0urrQGQqw5Mzu
97Z4RALMskFyDLdGWO1B5IPL5FccFvVWl+piVHL3eFtN1k2XXDIz4JK50BwResDE
OQ3BROAvZikUkTYGwVBIdwCU6Fa+cPn2fgME+2SRiAj/o+M48GErKLLv+wGXz4zG
FXLpdsgGn7FEzU9hHoojnee5QpMrJrafyvqpnWUA8jqYAaCthuPaUmrnDkFkJZDi
dHeFMzWyQjO7S4YMZ7LfT5xh9SrZU7sQ77g0SDBSQBMhLsz5rr2TAPTjZ0OfIzla
mzHA0VXdcY1m/cI0fKiSdMGsHOf7XTD51o4zQqp9UbYaXTjZ8AcQLYRTKfV7Owr2
CKFIUSxjGOBiPLVsBf5wR04Q0VRxSz6X6/vzB71dgv9xmGeZhJNwcnu6VZWdaxrt
6Zh9z/wMV7akLTKTRuxOYkpW8r3AFPABBux3FCZ17CxBREwQdUBl6pM43iA4voBk
jNNvPSX8K8oaOOYYLOyYi1cQ7dcub1tHoNoeooBiXcWgQiqTQsTiigVPv4j9xrGf
PopbcbbEXfFeoO5Lprrav08M3YBZYP0wk459lKumLtRw/KjTol/1j460eBQkd2AZ
w6tJznTfxQIztwK1JKD3CErN3NH6q8+EGbEi8FhiEMfhkQsGVYzL59mLoMFiHqMB
mIoWpyuU+x1PukoiT1uoEVJT0RzHnDdulNch+/lUaU5sodVUvHCUmpNaRlXWlKwf
05rEmJvuNFgpSoyG99NJbWjLQBJB2vxb1DXmznMIkcRa2tTXubFTQoWdMRHsncJK
ZG3LCEBYZbgSY6S5us6xEcfNN4eXUXUHOiLcMUTihoM5/NX4bSltf5Bc3B3d0IZN
neSr1OmVRDijWih9IlmTJlIzXVcTUM3syxAFf5e93gQ+2UQnmmqmQR0C+MN8WN+2
AkqexdO64Rv6ZmmDBC+a6cqv/3hltNT71SGl97SgDZRZvq/EqGMhLBF838nKwKU9
nkLz5ZR/kOCTMDxhBQSVeuyIYHqeJFO+1t733NFdVyjrjbAhINaXjuEZCZ01l6Hp
DtXzavJKIgpvpTz4rEhmnVzaKU5i669w+5BYsRk/OawK+wG6ntEUKGU23PWtURni
zi7RR6bh98VPdNe/nd3a5sPvGHgWM8pHpGCPFXIhs/YoHB5iBgoi7nLkMHVO7vrw
6r7CJRfWsEFqy7f/weDjOsP4UPBCamt+VIvIHNd5UP36Gaa7SfHTiinA5dpxp1h2
HbYx1ltFLBVfHCRCffZksvEwp9ICVym4dHG6Fhq42ervPppL7NIeLIqTx1WzB4dD
sXW7hyTzTuaimNZ5OxpDwG3Sb7M4kQtTy/ErYpN6XVT2dsvgCaBF2TWCfmdvOE/w
71pwpk99A3sHfee/+daq9ARolITnsnx+musscdZ/jOOUKEzJbZ+aF8MRO6QXooJZ
MncUenteX9K3mJWJz7kAkYyr0E5nBWGUANMyfWOBxv4VzVIYCCi6CKzg61lCQ/T4
n48OVatR2oXmkQJONxsxS5es1pPHtD758M3WMwdSOXL250b9EjLzeOugNkK9Savo
P7jo6Wk9lpEOcAKyaXWzkFBOKJ+vKo8wN2464kZhjiOYUruOsZ40BaV9jH5Mwqw0
kq5UAIRbM0PnFjisn6MCFF3svdV07U676AQNEvELXTzuJI8zx+8N5Hg2R5rNZC/U
oJjQo7t17B42JlqDwpsMjwVjxSNuE/Pl3zgiXg8WgAr8svMv9mxkIo2EGZJUr0yN
1pUEiCG9YCjUv5M2AxgW0WCmHpj+uDcMh/PGsyfZOZKwePrINTQOYBSoeu3eYpra
oM3xWGSWHdea4WBOR50okOB3yB+0FPNupG089YiT6LGrBBwwoEgj6WBNQyD37mN4
Ya3F8gNwpmszhtTcrMg1K1lx1gOUQs9Eme7MQC2N+nXUVcy11/yP5ZvQZj/Ao0rO
wmfKnufOHs05JeMJDks7FzMhNJ1gr6NEoQLrweU+FZhvZCyMmB298jL9zUnfmhf5
/F/kAXJ9AsPbA6HVzk+bffmRYts2ZZ9cVc/N5xT9EI2ut0hXRJ6g8nmqCSkQRDi2
Y1HMAk2lzxeYTCfZYMqj+NST64Ejy3myAlli6lA+wFpMKYfed9NRiCbxQr/g8GGW
qfnCTIoYHrTp+ljvXd9moQB3kzWDs8h/kn9VjiPWm/D8BE1fhPbGAhD2tlMs1G9u
wGkiIM+1Y0/OTuojOJg/7s+/AxGDT3gWokNLBhNfJAxCW6NtRvTiIPY8w46auQiX
M6CyzOcslOMPwBvboPlKwXrKJmHRcO8G6EmUBTEBH5WI54PH9UkBReJsoQDm9PXu
o2RzPUUji4+TCtRJ8ZxMBp3eDRPsUXF5cGkVYuzZPDQEVebKsnLNS/zZU94nVW9l
lQTCDNrtcLSA2m5bDD6ZojWTMwzBvUrHsl9hVCNDm516GkqE67ub+uYk8tDUNIUo
Xd8gcMd4mmIfzvHAkd56+EXVWswwsMpmIp3yiU1GcQEpbGIa6qm7v/l9gnkMWKCY
93EecNbsTYvyRHsrOxBuvoxh2c4+W3Gx93kG2ws6sneONhSY0trqGaak7X7dYNN3
D3rPYzrfbEytLmDjPwVgpdeo4YWNK+bAeeTCWmMPYolnHiafkFtLEqSvkYUo8nLu
QIi1MZVhLuXPjfwa8drA0H7aP1ZKcS+AlmYnr3L4V95D6gXzBgJ830vT/r30SbTS
yaDM9XUdQyvjxJ5EHABgsGVwS93Fi+kN8OaOLRmzeLBlgYv44ij6B6IJ7Sp0x3Ze
3vcuLmUE7KnmcpYvqPQrOGraoggBVHAVT/gtepr9kJSbDjG9ezKWfFgBSaC3A5Vp
7Bm/8Nc6khw8El3cue2fHyKGNSoGYpVZTe7lx7JDUgAhasJxEiPJS1W6BZSpW+29
YJKpx/GiRIv/gdx8jX6kysK3ILAz9blxGCY7BFUdvo6q3Gf7JqfIifXOMx0qgzBI
AxfLZrfub3l25wAOGZTOMgwPvodg2/2JzTf4eVyAWQcvPod/ks9MFLiREr8YZKU3
8Z6o603CORJr6u2u+HMSdkGZkBvBPdyAdupw+OvZyzgyC5kI4wxkCDWxf4EPrcE+
aIYZZ5+xHG9bv4TtxVH9CFstMrlJMPWNmb0jlyRdGsdyoYfFoMfQhgXMMh1afXHQ
EGLZBH4pwVc1luAMdOIuZ+EVR3gEsT8buEKJOsEvbAh33+oaGdB2/j0bIP3AzU7n
YDVAYx8QAeliBGgglmV0fvMtyYtV81LsKe/wHVWjEE7As0qulbew8SPKLybo96I1
ULiMwUkFnk4mtLAbSZ7iH34k6wU4wjZsi/xEwPmuOk2aDONCEM1Qtc3S57+gglw0
dQNN50Yw4L9pOGCnHQISKZ7Qbm40Tz8IMXoHyJJ4q9EO8rmy6B/vSw404TgB8aQf
vXELTZMRITjLfFzs6v9428AFuF6OCGsHq5hViXhHajmBU4MHauFLyPW0SFD7kxCx
HhTMvBc9XhPbtu+Q7W4k9hNderJTDmaJCIPBoS8rOxWYhjt20wkptr1rJyG0ogoi
dYF+yK/OVg+xuk7CgjCqrEFePAa98AZ4J8c0cGcG9Zt4WV4tnA/XIzliuu1Pj+ki
SCg8M8LPuFjC3lyymwuLnjWnEO2WnZvyx3CqZEHa03RW//VmfOSee2NuEQkDv4Tl
wJnae+zDUGUMftq9PqXxhr1vPkITWzSZIjgVKhcUrXywjuIRhMJLBDad2O8i+kql
FzHkJGA5g4BmFpvGE3W7PeldVikCUFkWo24jwZ8zmBb/4LwrTSD9DaN3dxIWI+Zg
5tCEldyMh2pYgJAQ08cGA66qsMZ55bp1UEVi+6Nkab0PWEZD5kbraTktIUU3hOqM
ZN2IUe5zfHVHgn6mg/HIoKBpdy5vihi4rZjahUiqdTfeaAfrcIQrw8pbuO7hCt+W
ZWuLppiqS48hkfHgRVJIT7LhRV2LuQuYAZLLFXhrxPyFo5SRE4LxHB2h9by3LD6r
CO0FBfA9sjwI05valnp/VIMnLM2E0hFFXNfly94jXMTlf2eUGMyPwhdRN5POBmls
G3rYVNzgPeJQOjvffzeDKJw8jlSklQztJxE6LPgGNshnPG0BZc7STtALnhGllIvE
vZkgS1LiX/pNNqb1jBZE48Mq40AspnSHLcdPNG65BpHfZRKqJQf3sbeN7aXZu4X2
vgQ8J23LuA59np00OXl75a0cPKLFElWyhsvmJCCR7S7MedwH+92OBx284iW8CINl
pIHYHSusW6rsBZDfVxePA1A15+RDnNWC5Qg+FpubNuFED5rPqwcdKyUTd03SmNNK
uEueHO5wwne7Nv+LEzcWvO5WDaNlH729IRBimjHx9h+5jUb8m9ilSqGA5u9qwr4q
JVVgvCLsIM7ouLUhGna0F3RaWQMrRqbSaMlo3+s7qJh3hXypKaXAz6Wc4eVuUbGi
2bFiCAMToOjumvy7quGvUYfszUmyAAl/C6qy/hfCPQJbORxwxVPQPfxM4xL5axNK
oJFx1jayLLqeE57ZhUuqZVXc6iCb19BOVN857fJMWfJ3XwzImlFr8c/yGP8EEv+s
S9SJEthMxEty1J6fd7qef/tbWIDCH1j6O5i2+2JyA4efi8ZGtjQOele/uUk1hY8d
I3zeM7VOLlV7CJi0ZtqoFs9NaollbHSgqrVwhs+2GdimRAo56PC+D6swzo6P1QM4
NzfuCFHT9u2Ew93bq+8+vnTGWuD1Nw+IPpj+QRucU83t4tWcEsEMg2b+H+08LBmo
T2rz3MgBwMVmbiD2Jh+uderty13Ue5YMYhR9dli2Xqi0MWB9j2Zsu3MdjCxRYuf6
oLase07AF7gE7QCZ/4q1uuns6/lQ/J3PDJPiiKGfWL4va7RsKbM6+OsFoKM4rMpC
4BFL0etLySU2ehvRWzdKLXs1fGO31GRC0TiA6mNBav/tBbKagvhV5W9RSHNuc47d
nUsS7W7rpong69I0mx1Ks/YzCc6zklwO/uhWLDOBIHvpeSA8c34DLajR91eUpkyO
F39AwDZAygiDRckc6pKvrnP3XBUME6XpDdJNZYy/0FQ5mqQPYvBwzfDFTSu11hya
Eb9oK+7KDh2U/SHNqGn/I+VfL0FdyakgfLL7JL7XbC9TN1Yq5eNvrYOzsvpJiFd0
0U7WzT4/stCtv1niLbtfaChj6OTQmaK/5CFKJjCYEWjfpNTs8PxV5ww3p9qGOiE8
BAkNJVm4ql425Zpp6v/ANk9OpUpTgEmpOWLG1JKkzPlaM23oEABiJRadwjlxbCbh
MuPPJepzNU8JhXpyk1Z0I+wJsesSXmQJ3N3xc5EssKkBi8uR28py9zE81gvVagKM
iWR21U6gOjQS5xKX3x2Rgj8lHByd4zl7RumD0jHTn014zN9vtbFLQj0sSxxxh6aB
qcIfm8GjB6JSw0FpRt8HktU9fxPWxDlPWx51k3v9ZiayBZfaWD9B+KTJL5iLEEfP
EG8gh4q2CLv2DjOoh18inzsgAw21SML/8jqrHWIFGlYd9bUQu3dTNjmkGFUlCc3Y
bnBiLSPIgbq6LY1gi4MYlSgwGtER9i/WCpROFMEp/USJNFQMbQRUHknR5Vt6q77Z
Mm6AeUITvctVP+0duqbdZJfong27obyTpHQcrO+aRX8z9T6pqic/1+sFFMMFQ4hS
GgAJMEdweOCOWt61eBjlUBUFfwfEAah/7BDFW7MoD6VRxFOrxaldEjloatiN2p3X
pMvcOhvQI7EU5/t7rU96gRAQI1U/epnPpXW+6uiB+APwWB3wS9KjlBIj0WexTczC
QLXP8lpUTTkVmVox5nae85y9Rg+bj/yruhMso/FH00W3UXNMSBuoPgn414VcbGEu
8ATsBpmmJ9Y1EEiURLLqJgqAjVx4KHQSavmCk/Q2TFp+Eym1rlwrg0oVmh5OTjiD
sjVGHNs+6HwccgPT7JWoXPgUuAWpgG+49Wn0gxtDw3k4lwFZ7upPkFmaNU4afwC2
zmkE3yutqGO8eSRn4ScJjhO5iC0EFGm75U+B6kw6C8/Y+URacGC/vxsHsS4LQnwl
TxPcoVLtGzzdbx+QCnJiNAonbWxOfi+wgY+7lsfU0hCKeFnx2UR8TGaro+ZQkgUw
e/KRhS1nJJAM7qcBbM2lOTlJWH7cwDbhUOnJoAOtJVDHMY1UXvtL+tM/PZOTf/nQ
lD9n0R97UVAT0Dv2aApUNSFrPRjCZbLzTuWZ7lhQI0pv0ecyDGt3mi08vl2YWzgY
Fh3NgqAV9YeYq6J7ygN7kleud/DOpQdld/PEkSpAfpWilX2bLjKm8+mRQ7vP0Puk
PAYbBvYJqDjbPSHgeC87HO6GLu0O04sB7ptwRc/xretQZO1c+YzGAn6i1eAvG0o+
2QWakd4T1tYtjkeWIIsHmIMIMvhZWM+Y82Z14APDXj11yfsvJtKn3+ipNTK5y2/P
Zrp1VlZSEZj4y5LUXRk+eIreNQ5ZWSC9H6Yh3yiuSd0LWdXLhg8TBziMry/kJlsL
BaJMdADQnHxX3kY9Sklvuv/c+HJvpUsVnaaB3adR8bm+G4bZfQNWfBdgnMLUwr5u
gF2JMHFBjXmMu3Zix6vSZ30WF8/hEO13aQKbP+V2MI9T32Jsy0J0DFOqqO/LzgG7
OtTk31heDwYD1qvyy3NRTNjZ1ZHKJnUOxop4oVyHv/cggK5mlGuBIiZ7nl1rCMzQ
oBk92Y/0TVpSQnJsNUlJgr13svjnIxUPOAApj1kTD2tiblHt7uiWYXuy48oTwVqH
lOGrEDjYc1SyR3I396UPqBIQpGAH39p1jWn50kf/krKSYczQd++mT8iCUgxMQ4Op
0fXHXfTwjYEUnM0z6E3d+YVSVDaNUyn5xLl2qItdl4MS4/5jnTrckDSpkcgGIYFy
TzzqjfiSrZjUY+t8BY6p9WamLDdPNFtnULCSF4Vcof0YbqXfzRrEd8puht9ndNJt
9JXivndfnn0antmF9ODyDwodDf8OIVehIYIDfdLc1DKQF2MrWAXnZwudQf2EUUNb
r6q+peTbetrGisL/qdZ5OviwnhrD0RCKBjJPiK1ZZ2nBwUgf9lLOQJLxJBLaM5t4
AI+AemV7AvLC96w/W+Dx/CVO5SmKXs7tfN3jWnfihbDf1098fSGJHvANFLF2lL8f
IjgWNSBtWOf2HOOXn/NzTybCeBxAIsSwe4Zj/NM/R+JE57UD48wVxDG46kiZWBJ+
dYepmGypLXQQrCKy/3PaHTp5ro6jhstK0diW2cqlgIfbgAc+PJQmrnfD3duny4zF
I6gAmrojLDodu7SujYVdqqQcvnitPJudGs+YewfzKWh60usN9nh0TSLSzD0ls5Us
HbnTxzOvunfI7Ybpjvd+3d+W+g+233FmwJmStIWWpfVApA2U1FXSeZcP9V/Xxot/
JsMz7DMQBA6j6Ost/fhoJMO9VmmpCS8dflMdhSLndlMc08KMpBaYwFabWeWM2ZkA
vjfSwoyTRhPkOR4Szof2BRDV7iq+oyCCTgpF4jHmcHTCXRqKIX7hsowMTqfjIP7U
JD1ORUN/0yZGsceWNp7RlS1QZO6Dsmj2C8wDOf9CPoNjQ1X0+H0Kh3095ZzoYEIU
0B8I00aaiopOBehM6aKxNFAYtCct1n+HleHbomITJalGEj2Rr0Svi95MAf5iLG1f
ZOLTm6EFyu2pKotSlVE8Sia2TcUZISL3jxbcwkLyWt2fy/XnuGSZII0WuyP94DQK
P3pBuhiYTL4RcB55bQY1M5zygSJYlcQkApCWbx9mF8Nwz5CSih0/Iy+eAAbzcgLk
UvltgVlSfNCuRBfDg8yc8U6OmYZmZ2R3SD2BspwtuArLiJeO+dyRdYFwsMhtAmPF
61Cu5YGIyG7nEBKgefqtpRbjvJsk5tXaBG+T7PDxsdKBUFDaxTDN0D2H3yKDFxv3
ZUOZi7ts+LuE5pnXfh5RO6q0O8BiwsSyK11iPTT4Mm/HBXcgNo0m1LBpQvUb4xIN
fOFOJXoCYpV/XloBJAUWK4W1S7sGDnFtB7k+MTo29fEIgp182uyHhhxtnNTsH2+2
iAHER+++d/y/oFKrK7we523HyIhA1as2Zg9eT/cSNkQkKDD7H8IKWjgFdNjinSHC
ORo9TcozK/jfP2WAEPzYPUiDBhaKGdFpx8YnWO4satmgP1nbQQoNRWf1CG/OFfED
/mXXN9ca2WOiSzibQzXgYzmCtTGyFRZeGQcdbAhQ6spcdrLMVj4yxNxw1u2I4DDq
i8t7WBdO/5T0xy5gqjhB5+6l55F5SvHQdyePZs4f+8gABLjT2Vo/CY1bvlfHCHZ+
gzNwsDG8Ukz3rHqj0oeBPyVu7OVL7XE1uQ/CsvzSbhyrjN+jWp+CwHqzH5uJOH+x
NZlON5qAoVsygQ5hNegIT5Pz0hIwPDae8kutm8wCNISU8L1Datl55i5HGmYCsFUq
e+JgZYR7WRtsZX0uYMh+lJkdjbCY1QFeijPnpxwlcMU=
`protect END_PROTECTED
