`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IoPP/p3VeApZM8Zjv2d/Lvr8sGOPpVI9+S6088cB1+z8ITFaZUcE3fVxx0apyS+j
mc6n8RpXaPQqqKCxG8xxummg5qXL/y13tViRcDA2eJGeIDb+5t6gSXKZ+3Sv+WGV
R0qWSVSTrNtwEk6N8lGPRaQkW/9B96L0r90ua6VUnIc/r8L2p+sQIkbeQgNXHs32
oll74AGEVUOR+jghEJlmgSO+1BnekKiKjm3wRDMpdNrq7rnqbdA6+kGIWogNvIgy
jdmuSpWRk+Xxl9z1XA16zHGCA5fJa/E6QG2q0Prio7gmK5vRVExkmcgpDRdUDnU+
Xhu1d0tCoSQeJ0IwBEWM2QRBkMggxQFNbo3ho2cMJwksuW68CsGDGhHhif8J6dAU
6DNQkHqSVmLVRiBboFpjo4GLN4zjLFOZtMhu+ItZ/EBmiVS8ElJzqLceba0svDp/
jN7/SxZ1KETVRcfcSGPngjhV9d1wwWWByd0Bb+vCEbQO3lAk/s/M+2yDjzhqU3zG
MsRGATBpmyvl+W5nVu/KtbE0cQTC2Xl0mtftS39FBrOyQ4IB9JsYJztSdUhgFuUR
GQ9cC43A5o7YvChIFBhK31z7aHlhTXyx5jxaQHnjNwtkXIkfRnwBX34mlxhvgl7H
ycUXWKRnF8YfQvzNec5qo+VdEOr//7tkxEZB7cRmXdiRMOXQJuhgbdFWsBm1XgLl
DFm55ycf/7js4MrhXw6sDynrnigXwIPdmIbGY5tzrB9rMgzMozkinJ/I/bnZlU1I
JBlq5t91FeRKPIFNY0rJq4YS3PIUVWDvDt9FdAoB8DgxconxljjsN7EyDoM777sS
pQh72Q99qj7rI3sugMTsXHYhN45S/fS0c3Wa5/yJ/twXiZdVftm0IQW0CTcp1aWA
IMoFbPaDI68re114ugJIbzFA21AgTeIsVN4PJzo0WU1KGy7mkjQBowd6hkyi/UVc
gAG4Cr5sRNem3IgyCJIlPfv9DeHrbP7VtjOhkEv/SibpblUtKiWqTkxVmkoEhsqT
uWc70Yn/F9bMEM/8qC2xRZtLtGR48zmNqyUKbuwqMKd0m88OXF/R7UYl9J9V5dWQ
4hm64GdCovaBpK3Zz5NBqKybBhI87dVLjiA3VcgBP1DOQrDXRLItEloYZZ6RJulD
ji7CG/dAl/lqaxpJrVJPSt6rE9guEEbd0Rz/tipJKa6JVk/gsvoHCPiIrofme2Zb
3b/c4HTNUPUsk9CV20TO5qYzzpHPg53IVPLq8zcVa+Bt/oiHnv6uVoSDdzkslRcj
TnQzeCbfqH7dIMZYJNO8C3x25/zXs0VGA/1XFs1ambFIJgq8vz06/uMkguD/iHA7
xlpoXdgtfRPQR64yFIfm21ajMXtf6vFBpWBgNKwwtmfDxkRWtxiVVroA18jngSHl
xTMBUOIFexNpdu/I5jpMWl46nWdZomsM78Ks2Cy/YTPvdZny2SeVr4Qi2NukbWoT
b2kplft5QrkatlrIp0gkcG89zR9h7G2YwkRMBmH4aAH/YSByYB8yj3vSarlALQl/
LGJ0i421CM7eJ3XAn78TFO6dCTgDErcu4CzZ51pKKVoZbzwRZG8AF5lKswezGeSx
Qvt+opWpoPGaIoPnrtXw2080NvBTLmFkWD7o21ecqq80l4phpPsTB5npUND7kVtY
QFcHnZSXO2ISTjbSwUIPdRzpV4qMwae5VHThlNom9t1DNoQSEZiddXW1IHWrqYS6
1YXBWHIVW2Efn4doAa5sBXi9MZtihCFEa4U55RdnOO4tuZ4VociYSso3TYp3nzR5
iGMrV3aY2eVkwXzdeotPk+VlIEnzaPNFCGMpckPo2iLeMHA7DTazETH4nZJYD/xZ
X5bSBDHxuEHYpv9ufcmXS3yE6zt9VMk59Y03C5DLUB7gSnN1nbEfweZZicUoS+xL
7lyX0vZc5Df568tIfn0N9XAr30W09lJAqN5j7vmltWVkPXD218hF6Pu8gYJMjbZ5
qlR9Eb29+VsknqMj67R0LOxFODjecfVfRo9WDAZuvbii01D6IQQ6wDpU98Cwq4z0
ka1a1KQXTThvoc4/S607KMA3onQFaXAbQ/UVUcJz6pLJnSNCJ3EDQ3MiOPZk6Stv
Mhy5W/1qGQYqaWFWzGJv8oHaZiK/92y/FjehwnhtSfawLbdSOZ/7S/qVEcDJjTLY
piHQy8d2tUlCs8PRl7Puw4fXQdgqMzI9d7tfFHsoVa7HaaqP578LUY7eCOwPLhW9
fXU5Ew5O7xe8CNZhgvizuuofo7K+79OcTteeQjbD8qcqnKl4TRW5X9MC2j0wVlZG
ZXLcuYQ4KLW8PrA33Vpbe8HxiF20LJqQtbye5+pArgTFR9ubhqdwho+M6aYdpqQm
DBmppY6i4bX/yPntxMZiU3peLS6McfJbWa29VV/sGOfO8A9EMnA/hDOsvMnXlV/V
sJx0kIDJ7moXAje0fev7/Q8IolBv17DrGb+XaAU76wFw/RziTJCylobuGNi5CXkI
EUpmmXr/XQU/W+uMDKvdpgYa9bXf42fnOxCeRfXgOiCw8zcNIxEvm9rmdnXgEz/I
hTPOyqeH43cgJ/pvFkUSHMGU58K/5jtF7rbYIAXQXkS7rZ3oVMktMlshvhfIQGb0
Xi04Z/gKaVh9wjMF5b5PPcroFN2hBUb5wc/pLc+NIfU=
`protect END_PROTECTED
