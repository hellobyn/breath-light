`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79su2nbmIbcmwOSsxyeqELvHZz2vm4JBCLbQjHOVLc4gMuPX2GMthwaA3IWxBbOD
e8LSH3YMo+M3K9IzodkCX9yTz1iP0r+qBPht97935TjBaJDtJjxhqsfvmTJYJcHU
E1vmU09rhxWGx8H2RZ2Y4R5tRSjZxiHapmyVJV0jZorU9qiVvkLxTpIt9AaoiKv4
bgCgaP9GRzAsR3OsjFYZs1vzkGJ0LR2DHrEHzApLqUPLeGPie7gOfqP4P1Dsqqo0
cfY6asvB+hLADYrvddcuy+xRyseONGd0ama32HS/TvKn59qRZu44Y4kju+mA9nzi
VV6MwjwRCpgJwfuzAvHNFTSgBTvu9e1hqIszMh8+SfdVdIKdAFwcKx8ARSP8bV6x
WFzO+F1FYFoDUu3Ji4pepEulgXpSjbrlQIwFfSJdsdAw6/nmOhu+RvtFaj2NNOBI
9RnUVQER9GYzlNHrlXh5+3fppyINg0VJj8JIyHj6VHADQR2Nfn5YSUwz9yZB63S6
VWf4oWDUllyYUwYeOLfJdvAUNHqzT0f9B2zMHfY2i8JpdIZcnr41xThcW8sN8KDl
QVb1bm8LKN2A9gjeOYAyGvutFUCXeZobkciY0B20nbQUuuZ+g0RsN+WvHehdFStr
6At+WE/CKRSfTEMXAVtg7o3KGzsY5pf5U3VZ2Dbk/J6LXFpI/lQ2ei8nhTydIH/A
t4kxqo2ypF2loH9HRCrSHOd9fxYU7HFPv4J8GzavdIOb/byY79IhcQPBCjfQkeYr
MuNpq4q04+JYolFsUtQkkF7UtszfQbr67p5b20QRcTEhWG07aAdgFdBr2XU1hqQw
7RHIDauUjEXmJR+sOla84HBTB7u6d8aJM19W6atf8ZGDE4tT2zijTW15/fe1HefK
CZaKvu49RhvAyI/Fsp5onIiUoR2kIA8wLYaZQyyjlM4E2g7fZp8vvMzjMS3802RN
5CEwjRcqRlfPFvPSi3XY8FdmFSYLksX8o01DeXMPGvHsPaI0/4ERuhqg6F4IgtHo
rG6ZKu2lynW5iT+aE6CaBTbjEoQ1mKz1NmEu4Bjbi8yeMZyn17+rKdZpV03qOhoL
vBvXqSZW1lIakyDCBeAPNHYI8NCfmy+iik07QfBE/5teUzJDAwFPM7HzCnWQ/G+4
PzsvW9Ktl4aU00ICtR3sUBAZVrFY/n4cRM0xbNd9xsUaR1ElmtpbF9PIjiB2j8/s
KvBLkEX4Igs2nNWRtZwor1OjfafJs4TQno33fAgsZHCPFNBDs+EGDCCJ2pVY0IPF
jYzw5whp8UcDPT5/YetEH4F1a1ydfUTGw4NhzUFFAnenVStrWM7xo76R57GejSeR
OF+oQlXmaHzyBKafqVbjnienI6ZdiXv61Tyq3EzAgdE1a05oM/3PmyIlQgQNdUGi
Pc0p1Tmeg7Bz04rKTURPBBEJPRBVQjQj2b6tZFADcgpIJCdsa6APQdj7RMaMwUDA
j0g+VyTT0WyUEF6Fxuezn+Ebz5ZKW8rxk0RBvbN/uEZkSRMpKOQLqH6io3knxaI3
StgY1JeljQ0AsaMa+nso1NNDkL5I/vtwIWuMwGMMM86Edp6vWkeYTCqbrCX1gcl3
pTmfXLIgPC9IH2CSXGpnrJI9rD2ws7aZVgVfJKScpDh/rdJ9n/K6avgDVShSAGxX
`protect END_PROTECTED
