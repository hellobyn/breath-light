`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Tq3kvdt45zqTvu1hcswd156yiZLHznq6CvCdi6N8aZf87Hs+DZAAHJkMo0dRm1O
3/XoBlgrNRmp2W9mUUQNuJxfw7Lo49CAFZVTOzq4NXcMbIYn+Pt0t3+ZGyC4NBdP
NTHjDjQ3tDmTQy2Qyu2RPaBl23sESQ2ZI7w6tvZHj1u9zPKfyXdCXg6EcmcsKeV1
o525Y1SdlMQ175IdTIyLSlJlIsARPVafSb001Lfei/m9NrcIlkxsQdfdCUFabCyD
dDE+m4+BHDFxKZN4wz6+I4aVXiwmj4MwDH7/fKo1Sc9xd6KWlx+vHw2u6rkqDZBB
GfEPS1qEJPtWjnehEyHahny0MdcIV09vuS1Lmfj7RLOVBpWa0LkF5FxVBJ9M3JbN
wzj751J7Xls2WCfiU+d2fA==
`protect END_PROTECTED
