`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBmuT6lUkyUXSxCB5hsONnE+EVwHrr0lukZ1JWbBdavRaNLPTWEaNYvED93zGW6B
SOVWgE5oGFafd2m1H+11NmwH8z+WtXjNu7O1CGiKsKR+oIkbLmhnIQ9nOyKnNys3
FgQUKK7PFhGHqI7iB0yOlQAKj5dtIvG6YyhkHsAlgtKDGq05i1052vYaJ8AC0gT1
ZCPvUvZSO9m9J4OtEGrwMdcWy5cHTUOWMFDa/YLA1WxCdOC5G8azt14KO2y4j/zO
rd6fIT0lBjkqQX2X4Ko/6EaGhSllMkSBYOQDpA4agOUPdLy+d/STOnral11tBVuj
L6MW+lUdyWwdrFdx0UNJDGApy0nszjUealKNnT4g9r+PRq20IJxtwnK41ZQgVr0r
gM8rfd9nK/hAZlAH2AtX74ecLafokninlrs3YOB4APiG6B3RAHv1yO3KuBSM9FHC
MPH6dV6PDVW9Bfa68+cA56Fs3nkTApxzETVGa310LkpWV7MZbzuXhjO8kHvboWo1
VaYhOoPaTC26cNPt0FCaXHw+bJnGVicl3CKhG+R+ttSI/KktbpLOsC4phAblnMBd
JFL3wMU+OmcZPS0OsEEegZtmxQH9H6QydF6tAiEhjLlrbSCvnsFVil7dKmRTpwjD
b/uDurD4bLVlcsN2q2V7jNjh1ayEini4LNReMJuGzBamOh5kKCc4+R65ZTDo2qUt
rI4RhaB3cBw9dKoCGCP19Cl5XdMuw9UyDt4t5r8cdZ/Md6n56PNL2pOoRHC/3ppm
ltBI9xXxu/ORFcG0X6s159IMn3O5t9L4nptSV3yG1sI5KzA6L3SQbwfZhSOxd6XK
157GzRs0Be3XBUuTnDZ3XgBwGlQbZko+YdAN/PKYrIsJWL7E63Q2e9Xpd1zCswxd
AN3hv5zCBqcS2eIfKcfJwsHJyYg22plE36O+JsqM9ok=
`protect END_PROTECTED
