`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ClzHohP458dFerOQwa7evo4qXDGtu/a6zSByLvi3uMAKTCzdR2PnwnPcNjeGiWd
g8fwqTjz8yWHybagSgTdMZHNA3LWs6/0W0OXc12K1km2eofU0kX9eeUkeZCiHDRG
m0JG8/Yq0Fz45OrcycPvyIQ+VtBs+G8VFc22QvjeTy8r9r5ZoQiFy7PoygglMI78
HBJaEWezNm+S5dUNToqfnxnvIpAH1L4hRPUv//vG5HtlJSB8EDJuytqr2Ug1z0I2
ZH3JRHqgBUoYbtyUo7dJutZxhvFA6RB0SfafVVOnT+rTtLXgh7BOx+5rMBc6N3h9
CMgV80Fv4YoDDgL04LYjALomf+oauBJZPlCe5DT4HUIISyLXd7Rr5pvrxQ+MSzdt
6P7e/6p2EnHKEKs5eOrhQB+v93DAdqErrz78YQj+sGwe5EgTBxzGonrkpX8Sg3HF
IIHdVnY74N6Vf8y5EL/3kDMFCo2d5/9Hda0Q+Gq2uGxrBe3PiduOPilAoglSkmjb
gW1Jlfkp2kkElDlfJHdM15L7064ZKoDkqi5Jvov6LKfnCkP5rD4707/KRL3yMmpS
HRcpmI7w/h8xnJeC7X/EFr7T7GDSSWK/+MP2FBmoMMTNQE6kleVXsA+jpk5txXfJ
2vHQIH3/2wRT/w4CsZFOm0r3AUBDQO+OYc0E+RFcJ1RL6o8Tc6MZtDvO8YzR+UqT
nnOcrfbum0jc9r/F+rpUcPzgchYVUHWJgHeWMdTYRuxA5sXASfX4YQHUU8tJ6KaF
f/TP2j3MEcUyDmidRL6/RQGS9zteEZ51CMYsO/h5RlDY0sbFSO7yJC9xOgGh3wco
qrdveu+7Fm51c6k9zE7Glos4VIclL0DDOxUbc8IdWv7UwflbYkuF2CnMEOVB4COy
HBO8OnqQJorDt69iY096vvqWCJ4RD0qgWtZJqdZtdQyb05JDnm9z1eOVb2bu9Fpz
67sDZgvvkEFaJPBDRK5TUERSJ9xA5TO2KcLqt/cyca9b74C/EC9mAHjUClboAFP9
Rz239tYkT4BtrB0fq3ta65bc8eHoeA7ek5kXlHC09V4xHl+WM09AuAcMjYKpAHaX
Xc+UQAXCuIQfA8oejKM70HTYtb4Yr6Cljzxj3oZsyjC0zcCJH7VwNpv5rBwWveWn
0mJj9MaP07gfrkL8Lcc9YHQyYMpF2O0o4RoIvN7DQc0TYVF1LXcfp5BCogS8q/v0
7717I7csp6O4MKGscW2uoZhT7KZ2ZRjBIZAkhGUr+nEMdjrSZAp8AGy7pm5CPE5u
9fh6Mn7OOY6wlJ1Bol04rhsQJwGPAk8ikH/zYL29+CEUtQmpKVgTUcfk3obKvZC/
aKuJ+xmXSN/Uc5B+6vNJNhrButsYI6VsvjBzrAN3/kxJgtCTvLDt16MSTtv4cVus
ZhWcy5B8JrDuIQhMcyk9uSKpV4Fpz6wwoUqrc1OUazHdD1oXeB0WWMsrDGMnAhmC
m43Yt+xw6quppeTbJw1OOmIt3qTfQpQ99pKLTZ+bTS6Se6ZJvCsjmmp+PO8LysZF
sZ1PbEUCREjWBdnqHu1speZ3dvon8Wx8VvBKl+S+F/mxKiMmYFM1tgt62lWnp59k
oGO4X0MBc6uYMqitUB0k6iOEyMypAYcA6rGOoe+IwvL6tdcJy3DjJ7l2xcM01cxW
RYkEQF7oEMHfWJ6L0hPWNXW4tQ+ALargY3H6zIEsdnwpcowR9VAUK1WewKfrrWcx
6il0ZPYWGY/NQhrq6Ej4r0VgpCyt8QKkRhs/gSQGN8fnkN2kCOF7D/p5NevAgjoz
fXwWqJ4UY+fLUIlmj6edNnZreZt0IKyc5xiXZahVmzllg0hG9NJInWfud1H1dkdT
O/GzpxNY16Bs0vImYxflv8m+wjgcO+Cajq0V8pLgov8HBTYran4coH6JG/L+3EGo
YXqXidR1Os7IE9icFYIGOsYgeOlWg44X3QVTM5y3NtmyGU79gAaM2b9TkGjllf9X
iZsYsq8JOoRbSa+rgupCkwdMkZkKeJbygz3as9GDbv1m8glw4Pniyhu98mUUZbHu
NxufSAl9NOgmG7Nz6qBu0y7D29WrSkZPueMP2M8qwQf0A0FnCBhprbfdcCqqxqDR
/tKFuL9N/LERERrPDFB2DDgzDaDr8Xet0xEYV1+O4MNorwdgKulb+uqQkCp0j1ww
IsKIFllUcm+XTPJFMd2+VDNFuSkSFYqt3VMOBjt8XIVns31++qi+2rxF/Xi6bqt4
a647u3uiZSPYJi39R6omd0dKQvQLY41fu/+CAy/RVV8k/c1QpFLy7wWBU3AEyXAC
cLVKyRWqe1afzjVnhby+lJTatKHnwd6CcoGZZuLWw4KU7QePl/dFTyl9mHtgKgKF
ReUOkHHk1qvQy+R1RLmcslsZ47+fKszuhHs32MkUOJuzdWhSbk0pbaAPkZSqdO/E
qpbY8W2VRJvNJIygnHZ6iBVNgWzXG8ZGkLQFjpRTnMVrfXrb0wheszDZPC51KAl2
fAX1/QEsVtdo5izs8QrDwi6BTNWT8K/oqpuCq4DAWFfMiBwXs4cHXHmxpoNhOGoz
Qew1JBxPv89bp4DBIX4gfrJz6WJWKchiDJUNK6VrPKsiyc9C4glxTSvFtHDzw5dz
bYXbmnQhnFV0FI1YMTx4vRtSehhvB7WcvXJUtRAo8D6k5FjhfiYMDK7RiO+Hb7bk
64dL+Xg8eXdmWo2L0CBWMnbW/wH4cwXnNtVbGllUTf7GhSqeVT43iqgzrAxchj6m
HCQe+pmgC1CLNDusRRqGuDA0An5rjMY9+yM3kxmAZTE0fYjDywco2Qbz+ydBhILu
zOHoQQyvmT1G6PkOEVrw5EL1+4CQHoGzu62eJ3w26S4qVG7YGzKD8Mu7dvHv6UUa
m7rWq+yW8hYaQ1hCGftfXuXfHOJyLudHG516f48rx0SJUpn+JC8wMb5wmlY6Z0D7
5WWcvJdzpsd8XZmL/vZpDDwdCdv94iR/w4e4WPOpZlQzqKQTjTKUMD0BoLk8L4bP
/jbcS0gSlX9elbZLtw506qHnyHlnbD+0SpgtD+jRaEsLUYgFju+DIo6zSdu5czb/
CRRWDiqzd/YPWc370E2R+7+1fCFuw6/1w+HPYib1KfSwEf4BYWIrqSciob8VUsCj
XB7emWOAYFl1dX+v19ppXM1YPrqaTlkkkZ7NRh6Zwa0YL98NhX9e8nihpvJrvGs1
E4VuHAninsqqwAcJR5WITkLNHtDWYV3aUVRmhsWlTD8y+SaSp4vVl0VXujaRHKud
wGF0GPvTMn54S25rvLIOi9riXrSkRSklfIQG3HgZZ2RdVLBfgBCkU/4iBXn/Ojs5
j6zJ7eiNHS9wuV4HvKzSvJcdM63FkioLqUfFE05IUcTEidkxsSX2v6k3cwY/X7xO
L+njREuQJNCFmn002q3LLkzKJYXZhh6gM0OLv7q62y8dXk9HhUQAQvlGAI0yrcLM
XhYW0/UY84ws9Ro6WaWCVkFTkZ/aUC0MbnP7o3scD8a4DEIbEYKTzgtKiiYQWK9z
S4SQ8V0rv+mYbipXcWtxPMt6Ed9jg+LOTRx5fTYp6BDZWVdSO7OVUNGFLBC8MlcI
I32kK8YiioEInF4oebm0wNFKDtU94HhOaDCc+ht9C5qeoMPmIFMSav96A4JPO4fI
OyaluK7iN/7w3g2YEhVYelbmjETH+2suwLr23IILcPK0yik0zQ7bJgPcLFr6Prcm
I7Lbm3Mwv4BG3KFl4LX/kUqEvIZEnbu+F6Z0eLv6pcqMMAv0KFP+b/B0i7wc2yQA
i0sCJAFM9vHRehQjO0dvkNZ85GFX0IGqTRGb7SS2iYx4O/zUApmCSR2mIlFwQtQJ
xXEkeLOlBHiTxe1eeMuc2pn4RLW+bwjsRh+IB/CRf/xKUXNB49c6AAV623g3YDqe
OfYECYy27OWdqfdACtG8HPzFOJFjoX14+oETt3CLTMgP08MTOHAbDbz2ByxH6dqY
AjuOldDIuay3tN7+TzKUCCBU/QwZ8Jv/lJnf28ohmUoosmohDydKkhZXxhs63O8Y
/Fv+QNcRMGcgne0qJZQPGRvYQLzDFfiXz9ZNAmYI+AUS7LDilvuYD3gveRzTWxNZ
VcmGm698emal3/26SNf5wGVIoMztF616MwowBYH4DJWyRbdVrf/HZbUjNm7XqTMn
c11l4lORTXawz2nmMX0FuKOQDjCAeMDeNADPmfs6co5A4xH7fu/PTHNSPGaeCJuS
LFrBgBzDhhm2SLgx9n253UnTNT84O2u3ZWEcuNgYPOf2T5e7ox4YW/GDbSxJMgSj
pyTMkYV06vBhaKSyEfgid4Zw1pv2eGlL3pHwBjAYi729WLZWbxJ62nIt6NdKnYJx
3zGxKAV5ffAT/1ZsgwH9GjjF0gK9kNQ61cUJD2dLA9OEHJlywsr17VPZM3JrwUi6
tFVygiyvVrcfYo7BHh0WIyZb1rF3n/6eyMUDZNbFXug1I8TVch1ZysY+Q2G+UcPZ
o+ZLdoGIWWTQdhCKsxj2xPOvwTor1z6ocA8M5qmlBRNxS999JMHSRIiDijxT32EH
0HpiwbuedR6SnbURvLrKTIMNP+8nFZzudMETy6zM70hKA7HoKGzLU2w5+CTX8KbR
Orxm18SCs+l8vOEP4glO2lUyM2uZoRrDFLkFjwhRn/eri3UssV413gLEIgGBUFGe
3QxlClNw6Sbdth2bCLLDGeRkDbHOJiBnHCf1bpkt6LX/TxnPfzrD83z0bWIsYzN9
OV19h5q/4M6Skvbt2DBwkwgm7Fltn2K8jyS3RJf1wvPhWX1I5w3JYL7pVi02GxkU
bd/99DYBLB2dEnQ08fSr4GFwuiEqKKvLcyS8kk/TXgjw+sYjp302xOai76HkZX4B
jQWHoc+7HLq3JmaayrHdAi5N0xPADZE2LZhwQZFnN7Wfz1L6mOIsLaAx4/db/7Uu
Hp4hJ+9QdX61GGI0Wla0z5VPxm8tZzeUeAa6EnZpmTKECzx30hdkhKEzG6W18Dk0
loaqJByYmn4wbC9zYVHc1e6hZa/r5uG84ZC+Cu69SBv/feCN7rdscYiHguI90eGr
1gFxZyuwfhS0pgGPaA0QJ7PWerYSFUnRQtRRuos9NtI4jpIukdKIr4vK5k67+dew
KT3UDUl92mubPME1sTJ4YKoZuwzheEeSHWZins4gchKcWSjl3Y4Yh0YjYsxfclVV
e/xI9ccQOeZlWpW20/2PsG8VCrG+Ew05DqMt938eo+rUdv1uTgxDxj2xpwU6hAWb
0zVBLpj2AOEof8l3ja1ysDKqvBIgqHpkGe/NG/eMhi6gh9xr/vy9H1fK5kyOB9DM
cL91VWd55svu9xVv7qi6BkSkbeKadpW+6GOFsMBPs0xIHAZ0rujo6tFH1FUnVnIb
BzdzVy6GBrILzQP95BJdRhlEAdBe9jtjwcp5cf6nDqdj9yS3gIm3tNxBVnIzUr/j
bU/YID697IxKzI0s6/UAKnH3BVZAam2tIpk+6TLF3n80yjw6h4o1ZGkReXH1XoE6
GwZjAfoHMP/IE6q73mqZTHG8lkoqkgxy16Sr4RV7RszMqMIUjhVRnfKt3uCh95+7
41sj6J6Hqbzf5K04c6I3UTLz4zibo7w6erbIUH9stlBfQtLVv9i9Oo5EsH9EZIMX
3jMoUvcNGGpdYVH/pxXqGMe2J0T9LJxuAAB5u61WvgdgoRiK/vE5ZMOqALr4OgRO
FZ7/XJOFguZAZ1GWKIR/jNBchEvY3zQiogJfHN+iI7mxAoB5HktB7IYX0jh6KEji
LizsTrWeWPfCE0wh+E55MJsguEqK9rlO6oQOUwKRP/tnDORJuCHyvrA8NQXdrJ1p
eayJ8VWUEOelkF+rNN0MOKlbmk0LhfUTYJVce1sb3n1v5Vp2mduysWxgQ3DUgzsX
TgvBI/M6CRTnq9yammDeMjM8Cz6C7WrEsTQwWFMykBbrIl/goURN9gdTeQ5f3bDU
rrnvjwnBRzc+IVSMd6Jp9Zj3q97XiRh0D7TCsHAC9twd5hubEZ05FPlYTjIpkHX2
iniq/3tpCKjOTUR6B8sozi7DbVgWjMqMcsXhXF84gb0wK8mSvlmU5L7gMV9FBc9a
jD9xKam09nNqKIbFmV4SVjdfUQeLe9c3sRFNkbJwUaFQzFVgwWIbBfsR/HFJ2JLE
P2xJQMmw6C1i4EQZYs2lvAsfjoIYMle3iWjuP+gp6zhJxCPWJZhjar/gNMuAQL8l
jV/W73/8GwyaLTN8V1Jw+aHlavwdomUu9VIEHggdAleebn5pfuW/vshnHIgAvBaP
U2NSLivGCQNqROTeb7hqpIpyFO/gaxrBu2nR5Ehcub7KZ6PnyMw5vRNq2lKbxmrE
8CTiCFdSvPrvq4qUQ8FoC86MSjKlGuKg+sBysjJuVeNyH7dnqCZd9VJnVR9On5SD
pVPD/3IWIfraAyK8Otos0iAuXdlkUhU6kqxsn8hEgGOLvVhTPMlVXdSlEOuoWDIn
Z9Cs/SgOUTTK2L+IclPs+1cLaMjwNDq2dZ5Ov5ZHXZPttHkDHJvZ7DB1merWdySM
EvBuqgthZ8YaBUbyAzvno1OkgrenC/LCFyo03imzgEbz1XtUXnI1at/5RoXKW1oH
X26U/hy/IvBhvWSt28TKxvdv7fURZqVVhQpr1BrkJYBqZhLJyrFexcsR5WPym6KI
2WjFgYmviik4n0zGXyPfCe4UwMgEuJ+AWnpByRZSd7CIlrBzZ+X19hVtq8H1zE5w
k3ESnSMribKiCGbz82heusPwQW+7vsCY6mc62X9NSZtHN90yfmrlEnz5fLCZxHqC
wan/0vAyX6zUKY/PqQFH17xJhidAmEsyIHMps6dFI6yykeFaO8hL6QbplgyOpxpC
TH75kdTpcygaIzBArsTez0oOws4i0TaKfFhHYpXtmizVjGPCaaFIDGja9F2y4iv5
+zrCFIa5FQw2D8aaxP31A59YEYvgo514tfIBmSYRJmq7siJ0DghD0uiraOa0EuAt
2DBnysBMcLS2cZZsttXuGjjtFdkM+DYy3u+6DddgMV6WrnIsXQP7jIkwZyScHmYi
ZQ635vQZgCdVBrloopVDOs5muAUss9w9KTyAJn6XMlsfRg82LD1Z2VjF36ldvQf4
3BNS/QfL2qJfno2LDTYn0ddOHjtsrcqVi1xD0I2Ul8Do1favRbKNv291X8LmQ2Yz
9X1lXdUcnEsDWBBSc7BcpGQ2qLOnTWmTa+aPTPiw8gKOn5TMJ9y9UM/v8FCz+d9G
Is06PpBOjopEmnL7NU1yM3azTCrg/9r/veQA+s9G6SEFcS2p3MzeI1PzczyjvER9
l8e5U/o2KS84caQU6BWB4y4hhXdoqJvuXQDI0motNxlbtnZ9RUx+bgWssQ7bbe6i
fgTFvC/g3Qe5iiONOiISdj9Xat1cgwOgn+p+xKtW6zbzACyhbEiCCXFUVod3/+2c
/7wyrtnhvOtNOkyKVHUtZhlqCE/gmzo1dFLy11/Q5iouco6QbFTdsipAIGX6Lngz
wWvM1OL8pwj6+qOV4d3QWGTLVwR1k0ucbX8JCR8CO/KtW7EWgRuxuQaEOBunv7Bd
JtdOa72UhN+35ISWB+A6kuDf/Yb2EsPUKL3wRQkE95XkcPR5LRXm+o/IasSrXE5Z
mIz8Tw2n9TqGGescIbD63jLTvsi9oIEAnAIC4pQp7uXpa7UHnWjUIIwMxrS9ckAV
hR38E1m5jcvprf5w/hUwU+NgLusVlf8fQEcx81Q7aFaBr0mvASEfIHCVBqQlYBa2
0o1yQVT0iGrj3s+tb34Ab+u1OywPhOll9mMV69vkh/2sL3GsQXchfAKS6znSP0y/
oLnCQ3Li5GUt1KjQEYoKnCWoVebFqLP6DELkCpaDGP8m0sKad90UNFpfKMp7W0pA
+kn3e6JqMgLWWtniKKMrDq0TxpkG4hGbxQPWawPEyok85+sYxyVFhNPvMqSSSMwf
q62s5eIWCueRBMZm86f0lmhbNjkNLBz4bvZXaWyBq7KuFHGKp2X/Q5VFRtKreFHN
66p32IfMv3ZJfe8mS+p2WW9gMAakX0oeVsAqj52xEOENcAB5pK0m4Q65plolyfUn
mhEc/DL5UXcgGYfJwH75USnFeOcED3d5N11piZJP0xVw2Biq7UAPegb0K+80DoyY
kdCfZWhj92OSYtOrbJMzwBoVFNOEvTenoZlv7xu7rtBvqEAdB4A4uOBTZ5hUkB0J
Y9js5wRcPKLzpPlTe7V30aPu2mf4rPGKe0Ds2OP3Lfsz5pXLtufEEZMqQC6vinqO
pmy+MgXxQYClS4yj4mIWHC8Is80imlTbNpd6Gt3u2dAAw/p7RO5rqa0nVaFf7+8V
L4UkXRAvvSFctGLuBpSYic7AImFdu2Rz5+/WBM4/d6vVhjQIlt7kbASSEbfwyWTq
eKVw8TaFc7Jg8DBOdwSXu2Cd7I6Z39YgPWzhaeCIA+5lRmgMHdzIkyFnlWnMcr9w
hjWuvHVWrxmyV6LHAVMqDlHRa53iDX+r659WpmNsBNXmQGo0uPC4VY2aSGE6s0AT
3hDyHRbNHGEHJw+meDa5zkwi7PMJRMRI+wfFKsB7Y5PJe4RwZiJPNcOHvma7RH4B
BcnR5sj6lozJksfVnNXbTRWNzeF/dLdWg6CKncPkT4zgsths/0XY6qbB2D3zWoug
bUMI0duZUdflWj4yGxwV/sLpBnyxQcOSlApWPa8sbHksqakoQ+l3mnYNokh1F+oy
P3yVPoyN3ZZrqtH7wMZhOCUANYW99QMqbfEvC7w9mBA1/7Gt6exA+N3kBrEMkcP3
3cJllPXNpiFO8aDD0MTLSmeaXMuqILXvevmGYdYbj/uCOMvHFyacYurUO0yyAu4G
p3fy8RHj92n9HHLqmfYvPWDNoG1p7D3TonJQ7JoCui9/mAPQ+6VRRUmXPAod3OHc
H5EGi34ysQGQGrA+GLMZgFDUIzXoz048+ifOEx4UbKVGUalDyjdaJv9YaG64qKyG
dRnZaj1EtO+9Z1mi5yc7LU9D1q8WM37zewm2EAJdmqaek3E96X1kIpfZbNUDRcVK
mEo9qycK2B1sJ9XoG3DL8l6qraA/g3TYuz+z7WhshvuorbrVkUcRfDL93hk1UNWb
xnaIAFRcYOHtTvTvZJ572z088sI/MCU0D/ZM+59llHFnCtetGBSEPOEM7l2DrHIz
T2o5gbaE9LDskKcFRQqya5eZBDi6Tlk+mXBCygL3UNjjQ2iocoTqTVo+Fu2U4FHb
EzjH2yr61UpAEyIaLZOPKqeUBsGy0t3CLRZDk8S9DsqB3eD2VX6eMB4/ScWbubqx
6CivcJgmgq/lnEP2PL/7knoCTl7Ci6L84pMRFtUgdegIichLYOdymX6ty8b6I2Hc
AZz5gy94FM7Pfr5hvncI9abhhkPNJa0rEEnOvfHgiyjEI+Xt3rnMDtsYe6+EdeI6
5LhA16NsO9ZKQwiBPy+FAoETS1PqucNJVs1/cbTx30vYRbScg71EHxiIyF8AmlCD
LkE09/+PUlJwgk12zQoq+iyVswitmsmPMQAKYVwRjwSA/cyPUGKa5qCrLpJrqo9D
4HbI6xjCIFOKwbngu8g0MGUbs/PNjWfLpqmbwJkp63cKgyVuyKNryRzZ+wzPemSe
AhxMrRqwKpVK1oVKE/R8nKK9YJZzIJf9Ehdd426lgGgnraUXK4EIVSTiceatFlsL
FGVt727KHCJMrpJq5/SHVzRLXsWMs/J03dMr3HO4P0Chytp5jvfDe0glVR0BbpHx
PIE+zCAhA2bgj7ZYXXLGCtjn7Gv2vLEsuUtvlJfzpBZ0iGq05cqME12SdO9g+Xbo
YDh+NF/KsRkXMHquZc5YbpsJmPIgwb7/HUGNXt4HXSwUbqZYLTXyQHhETRlyfKJt
dIuIiTRmhqLYUzi4Zk4lkaQG61wys3ZsM4cRvTE8GSx2EpBfojTdPJAKTqFGjxj8
DAIHqSueWHZR42hUyZhOBn1Cumy21H1482sAlE7hpd2iHFoTv2RjcjBqciblmG0C
19VN28Hxi3WrzQuPHzjLLlW9bsEs3RGOvcM1ry7i6kSrquoEEu3FZrBDqnWwHQn3
qD6BzqrHhc2vrrZfINseCjE/07qdE98vKoLvxr4dHZHxQ4L41IfjG2c99plfCMZb
2mMrofXsXIYOR+TdWL3j7zT7p4oBaLHo5hsniNn3FebLxyPvTypCRJS1j6l32IFA
fUmbgyGOVvytu/egYG4SvQ6lpTQa1CYH6X0Jmv/NMWbqEqFDiro6OO2LcmoShw9t
9US1A+nmu4PM5EviOF8DCohGKqRZKZfCJx32bdPKk+9nUFuN+S2v2mEBKFcsdSkL
qCEZASXp1m4VrTsqvQRuM6n/9bo2JDyubB3WxzqyWas1yX0LfpKI/wOIoMF4VwVz
tzWJTfsg9fa6LDq/eLfjaIPzi7rX2vnwZ4bA93/I2FzyzqsNVYgrpQHv0oiagH9S
megxtM5eikDIkEKFC0BpT08PzVAsLu6aHioulXNkDisrZ2FRlcwXwhTMuGGPCYfq
Z3Z44ASHItIK8cS2aNyha5iTCu5+mf4M83PfEioTa5nAae7QfAWY2psQg7K1rYEP
kr4N0IpApeOcjYVGh/t36riBdRmVFkOirZ5Oz39pOEahGLvG8hHrDl1nII1nFNR8
l5rVGNUY5ABBqHAygOeeW/uvxopro6acjeNB+4uqBcfE8zyd/pIPLyIvfrukBJEK
Ex/6fAnfTlaOvMZO8bGbOR3HNj597H1g5uj+bxtkuNvn87mDGSIlWT+BrBsABOoP
TgRzUyNPGKRq6QfvVMTFzbiDdsYBDvAO1ZfFDhTBBOZxYXH5q2ozbprCMeprrXOF
YKqcQWm5V969BjXF9mF0+vVyBdch3AvBOPtVvaHAmheWnpZTen0vbguQd5oS6ni0
WNiVnpwpV48XEFyaq+5ZwGRvYKfCmw2IqMidmk6WXEhNFa+YCxEt0nqxhiB6fWl0
z9DfmkyGcYUYatSTHnEZu25n1sCr43SlXnNSEGOwTVc+k9wK4RYVrPc0oXZuMaQX
UgPaKu/X/knKVRMaRv+RGumAzl/iOeyMX0lMvAPQj/g3KJsT5urZXC0ztmrNMF9Z
3SzU0mr47hmmz3UwOsDDpND5RoS99hHiCxhisugwhLVbUT4/Ewi6F6JaPNmjck/a
JMxf+X7jh4SIMF2fP8o5f3iuQ+P2OKulvGaTpO2KmZQFzEa5Ntz3edouwYu00rBg
sBlRjBBmtrmwC3XJ59c47X83gOMp8GiuLklx2aoMR7gASbNleKc5D0YVv9SdV4mt
j6lGxuJm6dkjgqVyayt7FcJ7A+7TDSX5TbtFGuzeDy9Y64eRaYtgyq3cIWW1ampR
BVUvncZxkhAk6eBsFc61WiuwkUS4tT/vKZ9gVOE4X0iWSDAZZm2ETP1fEVNRskle
bFCoOMHNvpoxFNyKNDs2++WqELAQMIL45uqTOIWuLmKMTq4S9Z4M4Tfeyz9YZJCv
Cy6F2lYc/XAfaNCXhG0p1USt7qZeND3jGujHqkg9OrbmS0ZW9IzpuF/GWbP/adsz
3JSjHbB/gYlnqtLcgcm+94wnc92Me3dfd+fx8cOvC8Brnc1g5UonN5xLbRzO6MaE
Fes0/n2cPYjSj86JlTs6B6cGUdo+5QSFZf/pzrPiUSHNRLwac7CNNpRkKhQg5YlP
MNvrYnpbvUqrZduI9UW1mXzNcoyuPxLrYPtZI2c4qhP/aGLLP4kFloOiifepg+m8
Yx3jJfhV9cht51O45QLzEaOgdkk2loVem1Rit2Vi0cqS3MZarX7baVtCavW+BTrT
6szUGKdS93trTCJUJyqUd9/tz/mmkOYGTvFvmDgKooNRTdr5iR2GRXAYZFFN3iFh
nOL726E7jfUnLwNsz48qwV1b3dlTwEYlmXhp+V3g5dr7uTZxsxmUiJtVPlF+9gYU
6OW86G5x1/x6riVqA4BFOeEiDmQxisyFGnVEOaB2ZTHAk/RFZxXoxwPuTlsujHwE
afoR2hty3pM4M9wRCHlfbGqNUl6+kjfukFczMYExk9fdspt3HbcHUPYCGiABRAqO
D//JHUIu0EX5TJTy6Xm3LvE04BF9wpPo3lyDlP8qSZECCaE65KlRFc17RyF0U0/7
lfWy03JWM3ozewtIWQSR1X1HncOduyPHiXbA4ixsWuZ40LQbUBzSmKE8UzhsBulo
TYsIV4pFjHcl7KrF40FhWlSvwlHHjz6ZOjIX6TbbDG/GMAeZN5uzvbkmfHuKwv5d
vg/yXjfX0furOlGTZtMTQLYEI79cycykQcExqXyjUnSrkOjMXlMrh73fp6ugh2D1
c4WIdsk5c6mLCnNffSeFa4Od+UCKBMn3WjwsgA8GdRhc3DAOocBBJGVg6IiP/7ZN
xZv4yqdvrTJehs7/GR5hExP8yp/ivJ/s2DXtAlg0TEExrG1QmoyWMYNqlVoD3EEK
EUwQpwCtfs9naa2pFjgA/qVdlGe7m8C7jp5T5GVwydnYa6w4cCHjs/bSDfEb4Gou
`protect END_PROTECTED
