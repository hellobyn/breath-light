`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HS26dvEHcP34wodsN2m6vIPCeCRygw02q6Zd524Hq/0Rt8Vh72nVWkoChirhJ4j5
c2YSIM/szQOoexSZ/9nGTrFAVyf6cXrIQ5xnWzV1elqNmhvrPn+TWW+zU3k7BFTa
3kIoo1vf2UugAQVxdwc46EI+hQghH8hxSRoiwSjdEcLGZVcXBgli4JDCXjgiPE8S
bGEqu7AjLyKXKHqCLY9rDaECjDKt5X5eH9Y0KdA+npGnt3gEd4mJcxW6z7rf+D/K
VnygxqkbUdMxlpc9yMLL1yovwVuqjHTUeZsg9zkE493VP39Fo0J0SF8AT8xqpT1G
yrgpVRuwgjX477UESnteFfIMzo4bKw1OSbkGYtorliub44tFuegGWdAVnq+Y54jI
P7FO6ZBAhu04Y/DyQ4FJ/J695eAQqygpjvk/AJno68jJEzDU5k2NKTO6uPTEwW/G
Pr6sW/flDCCLJSSTCdfvzYnleH11+w6o+HkLHLYTs042bvxiH9bD1FP7ORPm0X4s
lOXm9+zhRCxpMZhF82LT8uyVcKihe2ewXVBH3ayUkTsWxGSLb2zY8sUSFgWu9fYL
IcfAsMbJevetzBgtl7NzrmIRpQ9EEtZZ92qWbBxl4MmAEKoMaCtbTYmkQbsdcBK8
oc6sGkjdF8RPwFOUnSTl84G5yLXyzJSzPVboz+1H2hc+dEBYTWWAcNYBMI2DiCyL
zu0ZoTzzFp+0uLejQhyXbLZ20ErrH3eC6w+DH6DJr856L7FJaiWVuq4WE3/SS9na
j/76F3AtecKH7GAdtfSn0wXGCDJspNHm91kC7CIsan4j470e+E62rmdUgx2urDGb
ik8CdQLeyqV2+Vm4NB4zoV+aJPhaTJAZOqc+WMueCJV3WLDfyontLAlX1AXZuP6K
F/CIj4nmFLHfQXw17XeLTBm0ZogObLNKV9I+mbJ4Xjc4i3UKZa9eW9vTN9EQG6MH
IoPGccGM3qgb7SquvmgS3J/dSeWLPz7E/lqXS40Hcg8AS+ScrexSu/xd3y8ODdp6
CEJaCznt6rrkPKmnuHmZZjpS7VCcjfaEzjh1yfES4UfNglpKi+t3dG/3juDv9yJi
z+yD8z6E1PEvZHCStbeC0LEyPLb7hMDgi0q1nMa/3karf9x3/TWRTj9Jw4JhVX1U
nBSjMEdWKa7MGIma3jCHxe3MF0LQOXaX4UZESvJa5mJhsNCjSDuSK/DmkJphpDwm
RDJKLUy9/NuqctLvnMyMOtSEdV8D8FaTWE/a3/hrBcuDgP6ypb5nyqoP+3nc6Hn6
tSrKS1NeD30xS1hQI5nRLQPicckaVzKn6LYSpMYGtrew0iQy+kZOEHReXmgmw49r
tpM+Js3Hkyq08Bn3wn68eQiV1dolMl74maMKlFZsyM6WAYhbQ8HzD2hutmhEXoAL
XTnmpPGrFJQjPBkUO7gNkOs8gXlC+yeddPaWOtVkX9Z77rLQdZ719JLilfKpf3TW
Ym17xBJ6OVP/fdKamxV5qam+QdnAQznBCNDuj63QB+/XqHdYTkzUPvB9fjMUpmnj
qISNc2NuUHhEkzZzuJBNLR61o5NJNj/l0CWlqvAimn26SrKDztXSLe9KhtwBG0tC
fSN05nygFRqXV7tcQXz/uoNShAdIWLzSFl/K/xMgaX2AH/56kru6+l00D4deIJBP
00WFCXCj+yiX/lgkAApcUdtBVS/uo528Y5s15KmUwZisf8bSgRweOXGgzg/HtA+P
hpmJaOgtVn80666FoEd2RnUM+ZEOEzUE8eL/rIm3JI6JBWwG5OhHEQ14M2Gj4j82
5vjgoCGLmYddtAP31O1xryIMDGlKAA8o6IoysGwQgy915Z9WO9hXY7c6pfZtCcAn
Xs+IWHgaGKeL6JB00RT1I6TTLKvUfwRGm15rKYwUNz2O5RBNpD2ZIiVNSSo/34BD
xn3nCofev3+PmR1H/0DaDYKoAci2VW3lLvgGKIh0J9jXGCmBf0WRRBtU5w9V366b
t+PpDmlu/hlrMe0Kd3oNeM3BGi8r953UPSwA1huIYXO67PD+BQeKGnGD6MtrsAn2
BIuPRQIG+hj08j/Xe1k07Z75mO+7EEFZOcej0z5GqcLCM5kMFWLDaKV2y77yqcEn
7AMV8xBgoqmR3HQiLGf6qHQARDyXGfodKFDbvNp48oVD0IKJ0WM0CamtRsZgOgZ7
OJDbOB4xyphbvsbrzx6QyG3FgXWddubB5OJnOgD8vadJ0cK6zJq5wV17FxtdHxax
LfG/q8NYZ3EtqiJiRHcH9Rj2hjg82Y57uO5TYh6TvrKgA/jdSTAyqYWirF6IT7a/
3WF2w7NTOsqVrSegjKukuGhh/1M0rnHw/L8exGyAEbOfaZ4SNvYNwEKyCF5NHwBD
zQF09nrO1ApNQGcg0zO+A/co75/9Zy1zpTXO5spKZVS7PY0L4hQ43f0dGgsAEHS4
U8H9Re4IIv9KChNFUdNBlzBrYog9L26EwTBqTiC5yUkQRxJqLq5uhN9H1BnQj/lE
bdVxcIm3QruFfRUscW/Mw+jYgluoIxqtN5k7pd5Df8iw+Wcyn9PwUQ4YbI/z80tv
jtf2mlxgJWcKu8PNfoXt69VmXlmF9oTlKXnMS0OUXgW0RkGZGqb50ye2t91H+9So
vjmcpx04nLpw+VzR06oQr1iOpwL2unIhzmAd5QW4t0qyhCqsG7eAofrn71zvr0oS
3CIJ3eM2dyNNJ6WT6jW5InIu2+Hra/RFInQufYCNHZrRFJE7weEtv8MYw7FU+UCs
YfKPJ7Kg8DjR/88sOvXJutO7J3sYMAvRZa3VVASdlQ0ycK14q8tO+r8b32pYWiHa
juWpC7iF0j96/vjOJGEMsDXLrvC3Hem9SzOrmsbj6aIe6Bmvo7vhtkhCwSWCj5BM
st6VXaeNSzidGNiGDcZGVyy94AA5+b4ivcvSDqiFLd2Xrmq1kUGpjYlWbM8i/611
fJ95xom+08q19YcwaTkIOA==
`protect END_PROTECTED
