`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gNtHmxIvsmSQaSqZVYp9bnGrsjtFAH9rZE9E2O0QrpQP9zlWVZCTcXum8qAS1mZ
3hSB7xnBmahbOiVJENR+c/LswwquGfcenlyzrmHA4uUo1NieVSD4JfVMPR1ffF0H
iFkEQ2gUbKaTIQYCqox6UbofIoZTSxsTAmLG49Q5z0eNZjr2FXsnJ+RXg3U5TOEO
qy2CkxM2IynovGDvK4e3OB2eEZlXsCzWPRa5JDqFDM/qV+Rrw/oPN4gAvjuxbdm5
HxwBD76dDfB/VbkGhz9ZdxAAmK5a+HxqXaVuG9wrbTKBlZgqFQKnNjZPOMY3hFKn
DWYm2ph6Zofk1i1QIA8OgDCgiWaIzryZTT9Rr1IhYGBy+AfP02N1lXzdQJynbyRH
y09XBdCap2dEubInaMZFjOtlzZRktOQAuB4qYtFbneDPe/DMEp1kYTB/CEDFUD0b
zY0mfKoyBIfgSBt5zM6nXbRqQ7a7nJjEqzKdoTtJNjKbIXk6O6oSu8BFmpEDNI6t
zOr7zpH8WtdJIymxg+w0a9vyS0+TdPNxSmGMrKorh7NEwi7f/cIWIHP0M4EV9Wh2
iQUIKSABMBjf5S4OLLMzDkvfa+U/l7lIycMSywqY4KXR3k0kZLX380ElTa+CQPGv
Y7kCjrO2m7GXkJM2VNohtB3MH3Xo4z0d2Hb+W5au1QmpJIYqqPL712R1LgsmWT1q
y+h7liJQevQEMTQA79LqGpdOd6j+s4EiPmPeQTMfOWtuZ79kU43aJ9uSfu0RMYdr
O+/Y4lYYHlymjiRf6awnVE3+XQjWTR/DUaeclEX/g/vOCNeJoSU8wqxA1reSF+Eb
DqmOXezFusNoo/fsjfcPCE/PLNxAeFu7MPhbrI2LzzMTq88DjWhj65OxfrwM1E3v
xjRS75LKn57YzfrnRYOPjXWDd5cqV2erIpsSn2zNdl3s48ATsKZ3Hvoi+xofgIKS
ytWNqWqj3R3n+nHobWBHCNnfCGRoQDlpWKbf4WIBBFH6ZiZoQzG5SrKpYksdJ8OB
zzYsvgL9u2+ATw7Bb5TIP+4Cqtlc2yeTm54IqjPPy6Qqz4uC2XicVkei9Knt4pzM
4G0biqQNgwXlLHvmcUhJxS/fddV0LEtLdaUG7B7BzoaiFytTI8ksCxO+yEYSkQch
wEfVgJTyfBYxeAjtn7jaMMbyS3x5SdxCVuPHaCxfMBj+jGe2LMoupMs0obodBUNf
84e/mQMfcAYMTeCW1z+rlBqCYxoI1LHbDh7k/wA5rp1laZzsvbQVmuMHPD6gwz4j
jVxyukNo8TSoJAVeRdzqeqiYC8dWSO89uAw0lSNHYRvpfvwT9IoLItQapskWwPKh
+NyJheBqSIsSNq60wgpVaJ6DzCli6N00rZQcoV5mQyypjNjKHe+r3CvKr7CRXeuF
yAA0PJSzoftvdSdX+LNusxS8xqdgdmEG7GwrttfXByyz35uqdZ0QqG/x8CnrP1nR
pXbkc4quR/nt2JLUJ2nIBAY7sOXbsAdpILRUNxpTAHxfoSUYCKmtAUjGP0O+BjOw
r/blTojudd+Euyp4LPSeZisLFY+oDKU1aHchPKuZepXcOCCpNzJRdHig/yfjHSsZ
+CuZG45m54nBnwjkfoOHq+Zrw2YOE7TYiVxuQchmAPvvtgPrrKk3cGwfRC3wLLvl
2vSNwxGl4W45rKTkVoLfCtbdyqTOlozfbdNu3/8suHiBCilCFoAG3OS4OffWekJX
WaFcVMjZnjR3lOCBocCHURhKFo9iBz3StyVYysbbAsxiuDoPNTohMVGkcb1nCoQ2
ZryeBmrxIZ7HFYkC3NP1iAN8bA73xi7eSiftPnBqXQ38dCwxxXKHdbhv/AeQmvBu
hnLKhtiI0Q7Jimwu1XrLB6c6WIzThMVw91L5MKaXl04s3jz3DXIw6vlrb5BxSqW9
KV+fdArCKRs8hOpcH+lbT47io6gRcFKWMZ6fMUIXPq8WkJdJM57V6ObjKWLLP1jC
ca9tB12Gi5bPPu9BxA/w+s5djaNJT59cUSa8BiPWxawlZXZJDV3KooHhE0IxtGeW
UbnZAH9E8SUJM5zXdLGI7wCCdYrVIbphk3xsqRXgghMPIPUtyqJGQ8a5zBNPb4rJ
+e6G71JXObOP2x9x+T5bgZuyCsQnWMEhsuzetKdCT5a+tUQk/fdwnwg0T1LYMYm3
sF3O6LcYeyvivZ33BuZm0vydvhIyhrqkqVZPKw9J8ovnsLv+smh8BV0Z54RgBvKJ
cCsNExZGNkkzBBAE5XgQo8Tcm9tZQxFQ1f0tArdE/3yzysVRYP4yitmrGgEX/jW0
JnvgSLRKKcWW6jI+cNVeKjl5iNon4iQtRaau9mlu/iFVnoR6DMkkremd/2Gu6FQd
LlkBoCjIg9AVZ/wTj1MYlxArZXZjp3oQStV+qK8xT8Ejq5/JVY8RbtH3puxwOG4c
3wWUujLA3Reqq2gyrX6KaC8bw5oa2oxl5vW9bmbG0HxaxXGJ28MxKzIJBwKWyrlH
Yqh65t0USx5Ys/5jsx/Wf0v2YNsW1+4kseIuj1R94xDisOcpXqMroQa8+ycWOHG+
lvAAH2e7jZfVA+qXADpm0Y8Cg86nwkicPstT5nIRz8ZHHEp8snYCvMCBOzoCmGi2
Exa2nfhhRlUm9hR73HtAygPi0ageF4Y5NbRLx0jsGCkiZFbKC2OOrgqDUG/njfPI
HkozgCTuisHXJMb2rN3Nk8J+2el6wAlJhhqsGqX7EUOyZ/v2R5oVI9Nga4rWH0wR
H+d+LH7V9zBjWqxDLPhS9qZzCZaSk7Lkvfmgz99pHxTT+niDMrlg2ol6536zqzrk
VOOvLxBno+8w9zEGVV9C/F1/JppNstg+YE9yvDat6OixDkNs/e60Ub1oHuMmc2Xn
+VUQZhgyyHDxvLH8EgJX2YHvNCyP8jm5KS4+7VCZ+K1ABRgm7JLJ6R7yu7fGKM2Y
qBco+cRWLYYXGPzHWSfa1rlG6MdHma4Oimovz9nObShgxevXp2OCt3XyhYbxCimo
AApXr13IKv5dMwxMbGWGIpN3TpL0eNTeBJqIaREk3JkVMTPUqiYBYAFLECala4yj
sdSj6EsfJbPQ0QSX7O03cc56wE/tsIwjwNvOKw5aRipOv7nWTImgcDxSCanDPbzE
XNH4Qi6E/iTZKuP6B+k0T7wmtD9nLVKN1vAbrERFqbpaGERBiPnFYW8lpl/vqGNI
jhP11dR6yMCuqKzGZcb8w1UR3wNIVGvXej6vQty/H9tJICWdiPMwA19VNnwPT7vI
rcL671Gd/idKJUI69om0CNNP46gNPX24I5/+G3qs/ieZCqPWKrozg6S4I0NBQSjX
mfDIV31LT5m55iNTkI2YQt1TwaWBvHuWin54uHd7cFT2JmOw34bMMi7ybrdGJ/uP
tSxJYPCo1r8digQOzFCKjJ0gauERORbs+IAFOKTR2Yv5NpXXbhq6jnL2RZIffYfW
Ij5e1QWn14bPb1gl6zXfqzkDc4yuxASIbZkgNGol5ROlclp+0LuMfFwzEBFLz2js
fA868QIeh+Lk7J7REZnaWqkAgd+qAqC0O87DaoUCa6/4MWWAjky4eF/NT6dmO05e
JDzFsPCJn1hj2dIuQeMhakZ6RsNlLgU2J8rXea3xQmJnH4nzeUpwibDEddfaDl2K
hYZHQCqUncKU0KJ9UcWMtZw+MtkIrLkxCQerv2qUhG9WvXCj86Fcb1FzTB4tXrRL
pKZdf/TYvGOir7myPS061DHL2uk854wjQT8p8PrtHwj+c1i0Zyt1QNhl+cbJFBu4
0RE0FLU01/fReQ5yPtbixWN+AMfYuoZYHPx3T9fSYXn+KuHVSzBj7ZE76vPJcpnv
v/g3JXcwiOZFBReqL/W8QaALbJZ0dTl8iiuV/E33Vb0117tVWAEuM+STzqzzShSe
+4Cv7yJPiNAEr4pIe84viRmcK5lX1uuQmeZ698P/F5UIdaD+4mmPdu3KPy6nqJEh
CbHMnbk9ioAX8+QU+ZIATZoulSBW8W2NHk0DpRgvE0xUuWpe2+Yy9rlMkw+etVst
yxxoo7BpupV44uFwYbGB5JBvUdPmQNURtUqnTYyPjz546QOKuqMQGKUVB+LF29Nm
s6W+zOGZasMq6DYmGMj/i4sVywlu0S3MadMmPBLv+096nFluT2YQ0nEafpSM+JHL
KYLL5GyNXTeu2ndqlCqnk2V7UjAL05ouza4GEpp8Z2xsrSxNBojcYkH4vXNtdLBw
IQ7SoYBsm3zL1gkqm+7lOXsyxfQauYvTlaQLf2coJBh/vuZK5MJCQxbT7YIPkhYd
jS+72Tyw6ZUvEpURQyfrIdyP9Rh/rlhv7sdyhdPi8wMgxsUHAwdBlJim7/qA43RR
ajmMXJvucMP+krcYbrqVSk/NJuAtCvj28M0wppu8Jl1IOGalFAweOrceBlybKupF
HDDjIXfswhZxfO5cHg7+iY2UmqkoNEmzgFi8uwJYRgtK35/B6ZiEgr3UgcSAAwz4
C4xlmcO6JN0gkPQlqGOEx3yy5HN7B6IGEEWos2m4m2Ley7epwfmquV63KsCngsCl
C2g/L6154BAOXqcLlkmRqfTz7ZTaOVYnWtZqXjY2Q0TcMkyEuWKC9zjfopX+LqrL
3uVHw+xcrGst4bAJYMMRByuNi6WOgFaS/JHjBK8adxqnb2kcYC/J+IPoUVYF7DBb
d3t/Tr5v2ldm1j8So/8eCg8ctk0EhEc2PDzAXlTRMiwqV5B2P2rOtixlomPJQf32
DCc8IIRKEXaqdY5F+Zp+PT7mQ7mxTaD6SK60WMdR2LcAf+/0EKbvkho2rmUHixy+
2CVB8c/vHuOfs5UiV6q62XOUPR8c8+hMHYRyBnEzLWEYPjX3czfc+g4wEdUKDoN7
TSBQjsCffbsdjGHBnvVug6/LOrUFmftO036sCERVBop+FD9kKuIraIC45060Lkww
G99RTfOlzLCGzMInYMGsfg7y0LcTw8ryjiUyOAy1RcPiyotDU0kEEJVYByV84Z8K
Wz2d0sFuhxT7n2Dc7V9u5kjLpDZ5lhF11I3i5CvljdBiEPsW8dnCuCbbQsh0BnY9
KWtPtAorYQlmR1fY3SgQY1bxdaLUPS0bz2lScwIWTxRIqRziB+sOkAN6wZyXHw22
qK4QqhSOS2Pa4kDmSRcm9EhSoub0v+614ezp7XIN3FS5s3biiu5ekqGHW6STyNAP
sEYkgTiY6xYILbXEsMeebQ1I+PzEzBs4O0uuSMAEhuv7QdMpSj9Q5IW300vr6+bP
b20aEJfUO+A+8YFnI3CWl4zCLUloGXtrVdOL5UkO+/wjLF8cbqRXSqoSEj+fHEWi
px5lvUrttfuiXGOsubY60Nqoi02teQAzAjznX6rdaXCa93wc+/o4Gyy0mPj5KEGs
VFA6QrzyI49UQCWFBztqNMcvLQIDuHwh5dG4+zjWmU0WqTVBXstoKJKmnJDzCTaj
umLnAxSW+XEppAXQ7ozGF7272W+OpAK4sndO+WvHC/6YgVDs+8UB/Hbg3vytd/w6
wiWq82R425oSRt2FOp368ElwC4NFt7AOMoWCgIPDQop8XC7hOGvQhtktmWy7Wlmy
eRtgCA7FHw/GbACbs9EDdO1vCTfZbT/OhlcWKB6j2YVbdHcFW+Lz0LAe1BdjLN3r
hVtI1o0h3BpFEMOvnLvSfIO8dR460a3J80XeRLbdKsnanHIpgfJ4AbFXg6oX5hEl
i7iUMe4JAyiZ8fSlFbMBkeDS/aqO7KmpAxP4ekHLHrEWf6RjohHYOZxaO701a1Gr
g3tiBdlUaysHxmfLLxZIiyeGWwyJ+xDV5Fmr30RXNs/l89reYElv9x4pbcX781Qr
idH04K7UfSYTrSwryhQ0ue7HwATrugxnzi3Jm2aznf/QmmK8OB9HtgtUxKxdAFGO
JMvra3WpttZLxl8qxo9slsvtTM58xgcmCMqNZTPwb3AKB0ekbwLKs4oC0GAgMJsd
MUfdBK5ZS0HPgSyBwhAP9MuC8zTGL872rN+wR41+5SOmjl/4brkl8pvSc/0uBauq
1WgDdfhm37VrT2Ev1mRJjvSbDMrxxAf3K/uBIe99a3XbOie/ebw43Rcr6hWjWohl
kTxRI5wy3b+wi+NtivLs+aunStR+fozxX+/OzSy4vZYs1OutebabAct8DCzggk2+
feo3fbxSiStpuFIrLtGv3gA5ZV1iQ4oYCyfOxZrCLCtJWfYvNNMO9R+sWTsG1dYi
k3c4uDNMW00StiUlj7RYAUPJ+PvM2o2ivJlnMdgINRWu1p/erYxUrwU4l2yMKG/v
s0Vv1UDrZBB8d+q2Fov2yu4qHgY3Z0WgURz8kJKTso5puulvasi5eG59e/wCD9jd
Yv8N1tJbh8PdU3IYzbAqlD32PziuSFly7JmKr9O1etlTmmuTHvHu9qftrBqwu7+I
S+q+YQJca0hsmN2bMQJ/bWUc67ePcuCUleUpRNeZQ/LlTGWsgUpcqX90aJ4bBYCN
yL3+vvkMDvdTcV/VIB68vc3quXNBzKJUChi/w9BuUBlWBO7GaZD3DOtmCybZGnTd
h3QcWIScktlpJpkPMJQnSW3LZF7VJVnfdoe/x78Uqv54h+UPaAfOPmTiu89IUEhr
n9P9P6k66WIqqBl6zEOCtKOOUxSX63+I7+8zIBjaqqKkUXe87JkYlbn+rfSarSEo
ud/vkbpUM1t8Fwqpk1RMx6LhpLiVpOWXsu32G2gE1HLNNROghaODfzEmLdh5S6oK
qpsw/djrQGzqVzyzAfqKUqcc/Aay6qV4mo+FkOZIK73uUf+HhhxQ35rlGUgLtcaR
rx/0E2HR8kqsB7SU3M9IXs3euyMILIQZ7Q0xICi++CXdZB4CfHL/OeKdutVXy4XJ
4JI+QrCOC9TuBH4VzZizy71e6n1/mWQv6Un9jAf6SxNuCH8lMCFDSaZ3ujHlQipT
4Lu+/6d1BYuI/Iz53IvD41/uOUHc2nW6hJX94b+8oGlA9hoNJzVCzQy5zbrmZMkb
eCZNcDlLY0RwPdx06CiE5af1GNKsEzkeOC/qh6eiuVU1GkUMYkhNC/R6mDaWSzUH
SI/YOlxtl7O+29CSch4SBAUc3hUYQ2qlfjDoCWICKGjBwcpB6E3qgxe+fZOBmVw7
NhY1BZG0FWgGD0q/RjmP2HVi8kiwur/0zyXAJt8wPrHBGnM7LE/nCzzCwmulujfL
akA19z5is5V7ihRzbtdhmlV6o92xe/RTq5Q3Gf0z2aguJwPX+t4cQFveARsd2XUO
wL7+3Jr6sgFGPGS7RtmeVzH031oVGzeymEJU+w83lg+CTD5s1mSBEnB5f/yt01N1
psqV3D/tq4NdZkHu7dsL9mfB93ZCtvFyBWlH8aZQu5W7iUiQ8oOrLW34j+IIB2bq
VGQfq1CpUyGg3C3snH5Ib+UhfSX7Ki+O184UJrBve3wCnaLMU2CJ7Dt3PCr90ZAD
kbwS0rfNlF+VhdNBfH9nRCeiEWEKu4XVAdB4E95qqA+Pd9V56OFsP2T09jqfbLkz
MfpM+VpVTgedVuYQBkknADTLhUYg/GEFhaM5gIA2tDG0ccfV54SUySgBZ5atMvcf
WauptFYXppspuXlZF1on0Xj/JJYZWdX+EbyZfVni6UpHlIRgNMZqfdsBvSWPj1uT
KZwsnsIfF7qn8QF4w9Lyd+taMWa/y9cJ8xOpD/+Ocb81T+zvPk3i9pq8hDnOUpiI
fGCZn7iCzX0W4QhocHQoB1kNhQtoANat4cIKYmjgczLiZxNS+42ff40TuoLw+3Vi
v5tHTiYf9iS/xo3B89lGZDSIrNCxtWFp/X1ja/mVpFHqIDKBFrs4N4vLa/qwVeTH
eX8azX3E+l6wqizgX93et3NeEGdde0Ua+njyIFdxU9jANzPI4pNNHxfQMgpzqMQe
IYgqiiDXh+LdLbJRp+mUmN/5XFrIU8g76AIooSlBYvEgV+gBsLyEE/1dtlWy1k8h
vYr85I/kSSBwLgMnSqu94yeg+E3H+BLrYvy81KwQSLbHBuaojjPlxnSk+gWjSLtK
Va96iHEvJb25GMFZLdycNqAakREql42YkfatrQDxXsYLQ4ck0hJHxUZEN/x0YB5u
Li7YMtDcqy45KNYtuEtuqszlT+nZW2WDS5o3I6FCyh/ohAfbNKt+p3QbDKh7pfdi
D/ZToftVsmVzSbLytfBXCjniKcF3UCkXtc5ECwRDvK5pbpnfc8t/uLaxQA8u6xkM
uE5C5VX5m5bWZh0cNKhw2bMrueVwupa4JP6DICO7xrrSdDnNl5k8YWjVf46wMl2j
VYjV6qEvJ3V0X3QkGEP9UpLMmY1QF43YiGnAP0E9VVmZ5fQo6Rd5BURl0BQrW6Sb
R0EuhNWu+yUgCoBxhTLuqfzzUxhzYPPax5yaoRzm7q0/cQ0Inz0L2yDzw4cc7PVA
gBoHltpumVGsjKY8Nruy5XLXGleEPreaMSVx7qTBK5XaApO1bnN1kEpfnlpwSvR7
v76kgHS4cp2nBntQpbbOm0ZxCYcYj2DMRLzrJ5Oz8uRR+z/YVe6QVObFuhxidsP8
5KnzEv4D3TmtcGN69id8b5sqxeZh57U+IVHEKtvGr+Yp24IpYYFvqEE6MDXrE6yx
+Zr5JkthkI+9prObqOdSQYb/PK59GZTaL6RWxyu6Y3PnXP0kRlixKGd54vzjxtH9
lh+bJvEhTbCDgW9GezAam6Oot7IRSDxjyRyRVF1HN+z2MlzffZXknqcmJ+w3iDeJ
dVLVOTpz1lrVFKRsd0GMbC4usDhIaN7JfF8XKN4H6VJxxbHv6Xa9X3YUqZyXqgLt
pPQZTzwby7IelN7++DS/NJnp5answUO5QSKDyG8m+ryBEVpomo/rfTbmun4Q455J
8vOQFsk5YVbliePtYhF/tVdY4aWu4811/t9EcPxowsAuFRpRxLb9uU16XsQFiH4r
I/dnQm2Bw2cW0UAJmvZ7Pp78w0Lv9TpqL/KwVoh/InH/VOOdV0yt3N4dlr2GaLjp
bt2IWtRN46kxI4vO5fVWXtgiHIICgF95Crr9+7NbbaRixF+UHbXkEnMewc2i8r9i
iSP2Fh2K6so8JxUzl8xtoWWtZ1Egd+qNRAloa/KsxdU4qZE+z/rLnm/8sUKbA+i2
GV0AT3TbWSxbgwtIViSpa0QpYKxZCHGznbS/B/Re4lSsS42jgJ4Y24OOtb0+KY4V
rPPLmn6G/n9Irlb8ycCFIpUUvogc0mxQX0wPhN9NS6gMkRoG5eL7tgRSUYtuF1iT
aPGd3Hc50d5TEiRMjMRzQME5y1BAR8fwVelwkXBpiHMyKfJ3lV9/Pkcy9C3D6HYW
+U7Cz3+DTY1HU4RcwFp3v9BzNqeBS8WeC2URAum8mDIx1hdtKETIFNwvO/rzYCqe
eQMHUdkmsUwzvtHpo3Crp4rZxq4rwtv3es79tMuGJ2xbrxTx4klV2noErksHcLj6
qRgTAQeeYK0fxyipeflv2j9EOFZqT3Sj28PjY2AHFA6dIkMuQs6vQ6yT7MHBgbWU
kRDj/PD5f9EafSkxEls3HFPmXNIXBI3knmmZRmTCHuQbSVILMA+FxZZvJnKbh5EN
haIMGxeJiTse5e+skv/CWAqiB7WPd1ixIv7EbI6cwCAb9+MjlP+z5yWek2HEcl7o
17rU8urU0QwAVzlZZM4RAdgPTAQIFEpKt39CXiZH89yUadanEcvi+1hkxhGlHqk4
HldpSi1OaGpIoQVukGf1UWIYw+RbhG2F3LQjbC4oJOPQA1BZ5PzBk6XSotKb9aDz
NjNYfH1UxWxl5aJ6BZpzY1XhFnV2wSoBdoHI9RQ70ezkzYJLZI1cgKS/uhYyR7FK
DaPsdFH6qDJ11DaXdyYA6J6LZiQLxCny6nGPm1RnhsR4KQYl7E9h7bsxIiuVPaW8
1DMf6Kt5ogYYEib9l5Vbkc/2cnjpBmyhTFPzrClDzZsFr0CBDmfaq4ex/CVd9Plg
FRiQhP+MjtnRMnTKrm6bwSsrhARUBdN5wD463WHWqG6vhrzk9KRKJ8jwTXp732WT
BjIRIQgqrssYLCznwGYqchaiirloUjc127sAyev5/VtSo6zovy8tFv6uUlwb+YHz
1Kxu/Vlr8tTq5bd7tssw0OlcrrxMANc5R4tf+b29+0pT+p2YGAqLPrTyKco6zghW
815Pv5FC7vEqVVkdLeyceBLSNNm79nMT0S7udOAHjWYpUEQ8o/ezti5tRYw3fwMZ
1CYYQUBVc0wUVMeeR+rdgFkYnvzOra1JxNpS8yW6Ct7RA/oVCQPqm3BsjqqCzTsr
ltssuEv8yqvra6P1SbppJ9O3oWsMGRD1qu6NsDh2zJMu3okz9eIlHwovpUPl1wl5
mHJpIS7KIsWGPwQ35mn475uni2C5VL28cDID7l0QB0WmsCGgHUmZeiNmsX6w0EdC
CF2wONj4yO9Hyx42xiwwVfvF3AHHMXorBUiyuiiG3O7mCPVZDK8BWAN9Z+jXNnYA
j592t59Gw6MnvbHCYNthldgD8Sd5msg0+C3liNastYfjiBNO+EyCpv/Ph3Vu4Ymb
Dl1Rj+tINxTFg5g4ITYzXl9hjnG7JWm2nYUL5T/dPZ76ghLWWU+/Y+q2CbaDNNyL
2aZW5aRPJhzVtvBOz4P+yV7nHj4g6uxLC2L7nksHZq1v7Wnzy+AsoMp6tmqbZDTU
MgkIZlE0DXwUCia+gG1zht2SOFjT50l4IGp0plysJPhKvGJAkNWtnMv4n/76H2aa
5r8+0GehZY+jx/jSWY/z/5SOVmrh3AmV/h3f/pJ9Oz+OE0Dhx4osI2FbdCDYl4wX
ABttCSaVN5ZyYrFH4cqEY+VDVmPCOAUzjqSaWwiBGbpmEEQ5U4PmgMOjMNhMlnSp
9r88YQc2X+xv9w7p+qEvYz3gno52U3xANRm3JdDyV8lKQhSVbwDWeXobYU+ASOYP
AINMaY+iuwKrMZVPjmL4M71+gt9OtwpuSCd+vj0tGd172/U5IMAeu06t/h9lkMwX
GMHskRe2iFCq+7B0EVicSk6wVElKf/qp4h7zGlLqfScXb6EVMiO6CUV1gVqEabyC
ADgdyKrz4aEFb3UT11JrSqCxdenZJ42HvNUwezQD026oXsVUdr5qSuoPAg/OfIey
3luqzEtWpuwtT3jYTQmhHd/6qBCLx84uDmnooKEHU7kb6RjRZQntz5OCEc+cObS4
Nw4plAs4F3ZKsEGiqOkwXT54b3zskhKXiFO7LqLxPmFC6t+9oaXKkT5mzVeWK42S
/bttEms3erzaZjE48tnnL6KrMResv6QUS6U4pDDpB6iEpyFBMDans/BRr5skUnW0
QFKeeEy5bh1Z5YRTUHkk389bgMpndIj2wcnK09LIWgILNNa4NcuAAStMPoWLRIkq
mXSU6K/WuaOcbRVFZrele6KiTe8W+xrLLGKXDx3Gktpxt2lA0JBa1vjNhW9KM/IM
vLNvk9PxNfbPmRuZOWCevJEEhnnlckfjCLaoCsiUU3TG0pqGCuyZNQeLJ6MXMA9q
np5vhcq9/mflNahriuJhz9jBVGlilqWc1z1WSqrouolk//q/2p6jbaaYWMKu3kTt
ytrH9OZxznI+73kBeJT6doQ3HX9SE48cUc/bOMblKsca59lpOQNh/EhGdFystDtF
QkqjHdud31a7rRDzZwwvr0j7CG9KtEeF0qfg9ilkTbgkFau5mF2q3y687dru5+/D
Q+dI58L4uqWHkMB2LhXHhiYlliQwEk1Y9VnGNF1s5XlWrGZcgthFtxQO+WQPli3P
ICHgJDVIeuHeOZBNgMwceDdgLckl++wisxzdH4XdioN43EkXFuXk1TD8H+NxHbwP
5XZvQ6EtItqT6sVOEY9FVrLRZj3Sy7XFre0aQlECcMaIxg23JRxavN8Zo03x7zID
+0IIwlBNZOoz3YFj9yKJ8FsZONtBjW0yww4EoM++4bnPg+F9xU5b8p1LkjcXIgb7
qFmt0HFloRWHUARyRnyjVI9D8ZOZInS5DL/b8UAaZmMHMdDQvNaMY2F3R4mq5IAr
jhMmkwWeMzmJV/rEOLNgLOQ+eZ8htYZ3NYynQR6nMV8lqZzdyeV9T1LsyGecHkC9
5zhCCeL+NJ21Zx4YkJhZAd25A/0dbP3egrPW+7Nx8HSfZa5iZ3kiDesGiJgCgO3C
L1/Od0x7f3rWCl9YBp613V9CuP/+urbJ9ka+wDt9l9VxCLg0ZY2LL7X3l9xxHUom
l+fmmcGDpDDRn3pvcpzVr7P9ZpSFOJTWHZAMgeTPP95z9h8uwa1cOWPTzi7U7+vn
eVR+8nQkkT3eDrd6uUmgTTan5ySctLl+sXfq36zhREU+ybcmOcvXCd79aDmblT5J
5/QfY5Lwc25OtuSy20UdAnfqQ5Dn8hhIhzDTqar9AiT8/nCa/EQnnYX9Cxe/8/H6
cKkodzHGewIEVizsZtGW7CXLK2dB77mmgisFXYEhJW+OgDr1rxLiBBKd9eWo4EVT
Lg8bVn+cZpVBrYiN/k2OOVjg0e/dM1RtMmO0XzK5fZ9FpsTZH8a4vfhqqf0s4Myu
8NSWSuC4ZwvAi9enPlJsKyDhzCTwV/oIOZJ2mhVOIS0QTNQFQIYbMxojmHLkYPUG
aZ4ZNYe1hWK7aNfqfJqds5vqSHerd1qos4sVgChAJL+jkMdITS6dpfOoUGjZtZAf
G8m+WH4XRheEn2tLTq/y42nAkFeaLrCPLydJeg0iZ7YMZWr6+0AMkb8LpL3rCaGJ
jhxhQdaaAsa6QlAI5KjtzbGqr8h0mH6Zd089Jz17u77MFNOOki8N1VZrsEVUUcxx
Xe3Ees3/wske9kW46B+RfmW77X+eH2eboGC3T3jQWmtc2/fqWvHXX2nIBxvfb3cP
tPiIWoo/9t0wrVZ6jAe3rGJvidqrKaicTBnsQ+W0n6lkEm784bbPpNmk1CTbGlgP
FnWomnJ8l6ramEKTN8mGS8jbl52lDfg9PEtTTj5A4Z5I6uH60boTtsmPLmWUKDwf
i/GH5ZWUBE0RnhZbLX37Xk0IpFb6+nQFV0ZH0Oy0R+KuEUvNPSOzNP88jSgDYR+T
ayz7JVdS8UGkYUjix9GIWyuYEPkh9T3qUMJjpCEWDW9q3+HUSWhzpZQCdWLuwaDL
YoddT/06+jVSHJT+O+MxAiw6IFYDt26L3sT2xAYwUoKWZY+vwn1gFw9IvxqVCmIJ
K4AxBx0AirpGNusBOxDK7ZlTu9hfNsuOdZbzdFmLXfRCQ30R81/Q/nhIWaOFJm3p
SLvO79SVcZ1zYMh9m9m7PXtSqrX9jvJOFjGZ/OQFV/NbeSGX6KL6hWTh+jG91I6O
3zpdujP5ham0IYSwoTcFLJkpz4gh4NcVVyoh6IAHTByPP750h/++q3csslCrGJlq
fuzQYZiVhWltOigIHjEBYanhM7xrh3Ian/NbsZ5i+6aQuI7nQrZhjhEaTVxrm4KA
Ojhey7NImi8zC8yR5hCXh47KB2igMw9SjA4d7A2Two3dB8HjtQV+B1tIcbSZ0Obd
9y130qE+yjc4gnd8SCLPXhswH+/xeCFDBmCYtmGbU+/bAOXgfxCAc8zFHs+ojgLe
tAnCKP0Mojw/QIEmSU9FR2VO/55z4Yu8wavyJcMou3e5Cjs1IB0ODqGUr1V83r/X
PJgRyD1bnzAsGGnsbHqOJCe+KSy9/HBSIlpwTP2zbtAYWnQG73EggrkWsaE5ee6G
+5SQI9h356KC0W4+aXaPJ5xR5k7pOLv692Qr7hC153KWiMG4z/bJaf8vUG31Xm+b
178O3FKLE0IOebUYA5VPgQ9oO1cChrjzqpEAvrdGYIr3NF3gNoTPMIsLUVHWuciz
AdKSwhnCe0dzvsmB1DeEVdQl7hx7V8mT9Jhxlx6vJO+KXERe0KaYPKC3QB1I5Gne
zGwwUlGaPgyEis0zDXe+zY4hYjqIvKFlpF9lxq7W0ZStRrbfDrpIzPX9mfdRuvW0
Rw06dpvgD43KvaUpTxu9xRD3fEyqBmfqdpoEPQhunnWnjgOzEKIZQCc2PMy6GgB2
oBBwQ/WQwapzRd7kibmi0wku8/gbz5RUhGIDySUEl3/P547S2K7VL3e1A4/iDnYP
W7Znq3Ygqccr+8ACJcq9KnhyOuDAwUpCpGJW2RbPHl7+xoRB33spHZHN1qmcFgUd
sPogJ2gz+r9kX4xM/BxEz1fXWYl1bhMLkvHwnS/0WlrSDlKBMAK9stLKb9UIn5hz
cMKdGKOFUtDi5wBBXKw+f9rfXS/g7H/qjCZ3FccEmg2FYn+O750DCYZk3ZGhYUKQ
fRPDRrGzyNf30Nn2eCziapUM+f0x2kDoHH6DoGvu9l4a/T80YESjHGIUIed0Akk3
kgZE3rNgw9AZ1g+AOLHsrR9RgRPOf3bN2itsqQkRdX1aup6DAn3DdkU/7IppcyQK
GRUZEO9dxGJPBGAn0gaY5WlxQ6+rY5pHUDbkpnkzpWpt0MM1PJXXAOZTU7AD9SB9
wqziP88CPVjMBYxFyHXA5GfZW1VExvDx1hCsj6/tspOirXUnNMCyzNa6VyMc9PGf
G8TCOkUCNx4lTlAizjLsb6kD72pUNY8W8ej+cOEiKhxw6CxMd+5rKhKad6IirN69
TCZUWi9z8QNdzoDpRIFU+T5BjdOsIdS0vIER73ccbgBvHp7YW5Osnhn3mZRqQ400
cpuPiAQflKVm+EoyExvOfbcvXZ1BHin7v0odgIkP2x4WTvfYscF7UjEiP7ULoaCY
w1yMlVW4uFZpqaXX0o7GZB3T31qxVtxnrbbUv0BQb0/03979n1m3vNrne6MNSWif
+dQr2TeJLYwBjjjs1NYKEHT3HsuFXcnwTeqvIu0yIl13QYrgymGd+cAodJbsidT5
fRnVRDi5ffUDH3M801gXe5Mc54C5EuoTYg2WqEvIWo3O6NSBVLoxl60cfxxVYgJA
ER02a2KWR3zmNxJjLRiwB0Oi4XqmOTTsp0RKbJRLHf/zf/sB6aVSCq5sy2JClFdZ
agzn6XuTqjaY9g/fjw7ZkhtoGnB4+IBUSR0mXQ6SuF14G3pQz6lgssGma074Xy88
FG8nyfbcTI1lRbXcAvN/B4iBtsH0CIoDg1Jkky1YWUTuU3TOXdY8RJ4X+4TV0muw
gI9lb6UWtQy1iMWC8BzinD86Y+anpDV6mj8mwhNmwyPEAMLqUBr4yjXRR1mUJ9tr
MAOtbCs+MDNiCBfjSifBhHJC7MOot+GKrz9mOtiWWs3qDw86Q+CeENNlAhKjcNEz
dw++jFw31Us6CthI6Lr1LMLWhDVFvWhYWOe5eizULGUqAc125JunD5j7E/cAS/7B
zQqh/NB4nNATIYjc5J0Jxa1N8L7eer4BNC5MwfvcFS3nL1HvGjKg0FfHvwpO7Z73
axtgmxpDbCExTSDXix5BWhMTFMx6xvzLjEVmnMs+4PYO+MT7ofvwSzlON1F54qD6
DWBln9ZeoKMdZDjsWLhjLfai++O2/elwkvH3naMWr0GA9XLDHHHbJd6wpDnyfW0j
bKVSrKLWJIyl+/BLMfvPDkVCmEvmwiTu7NgIjkD6eaIjhaKG5mXcfYgCyXENIMN9
JNh3hUCzYvuNDXOEeELqug9v7t0QONeEEhAdEywuqAV06+5F13bH/lZN4dJn+XDz
HWIZ+sIlXqN8vChRFBk1pTZC4S8lxDMHwKFGTaRA/pkxrpkjFVUXfzdbckz/sqNd
x4GjQw7/FQLx0oIfoQkqq86woy+9lQzpwn0tTKqKglNIAuQRtm/Q9BECuPfxH+Mz
GE85jmJdVH3md1e1uG6he9BQat5ch1F6ndOaaE8bscIaRjgZ58PLkdiGCdjq4W6D
gNjqkSSUBHhud7vPQeqERAso621dz7FzYjCZ78kdqq30jtA6LzL1ME2t4+gMvB/Q
5wa09EVygtTL41MqKchWDylaVVON4C1rR9rkEHACj7f1l8/3pNXRTTAdh6I3Wc0M
hoFTPyAV8SWnKVJnsdyoReR+kV7/ThwJ1NhgumxqoRxC9smJYOOtTiLWbSdq2qls
NyPx9kW9C1sqd5pykN+aNsNUCAo7hqOWTxjzoGS+J7LyhwaRt0RetBgNbJ4pzokA
NfWr3kV80B3pJJkWyy/+IG6pBepe79PYnU5lnVCzxvjKM6JILV4ENEQ0UJseBk+D
17qdrcibwHwDBAPzNmxuf9d4v3bLqa00exdrz3VPh0Hnri+B543sqX6NRAC2JCiJ
k0dE1ll7//mtgrucD789jmUiyWUcnCNiqyC6vxz/OttE+b3V/qlDyN5j8twWQj95
K1F927hlw3bTRy4dxEcIO7UJ5A1fyTbQyoK8IM9fv9x8z9CMl6DolJbo9zi3QlYT
KfmSAxReRkgQ7cYp2Ihi8gBGlg9Q57pXn2O/OSsKzU0mTzFMZ8OpxQtOOW3el0N2
B9mnGpZWAMCrur1kZLM4Vt9zvosWNn0GXgM8OF5kzN2+jqeGJguP1d0TQnmma8PL
zLLqihn+Nxd+OMWwJ+D3kZzGvBo8TqaYM4oRwlbmd1zQmbDyK8/BhBjEbz6HDZOK
eUgtHSQ9cLZi1V5Q1qOu46I1T1rQnu9W4gkw/KgPmlYrkmNfyF2glkb8S9jHl0EQ
Zv8D9SnWXT8+Xipnz6PTdFn81Egkwr+1mIg0zSPLI18QSRrJRja8sa3jNvWkCPgU
7tnD40D8Z+Oth+/J71D/qViqtcUFSTaQsjQrCIq/FxG38cgNtJkOszgt44n6oVaz
43A4h9/6Q23k7gNbUZPSNO37WEt28wnQY8W3KDAyiu4A3ivqFrfT/3qP1d55qnNy
jLFjMu3DUcAgxiD4ye1e5OF0NgtZjsrl+q0JlnfhvRWyr5Jt+aI1wNgsIfKtSaFT
4CbfVEZPbjrP8oBLeV9EFu1Nwq7aZ+KAqQ/ZokBKTK5jctCfjLDbBsmq966RvPRe
8iKrws6nR5FiV15p/raueY41mXAdhLGjSDzJZkxX4iXD0GTfWnTqX+UeVLr5Zgls
LfnXKoo0giqLkx4A3UEZFAGi2S82/ElcPwGg/eXgQknDgghEKBxuUKoOZqBXiG5x
0Av7ghmDM6CWjdBD1yMStr1rBsGkacHqwuzHNSuW5HIfSXBQdmgHQ0G2HLvurdCs
ilnhMBkrimiJpeon+hVoZVc/c3TKe7MCkidHFPcv+xlPBJeXFqJw+6yRJw5LiG7w
sykmg4G0BZNF4q+gZUddWD18R5ge9t6e8QNQfkqM2vmwXelTpJdITHsBVt+qXmeA
FX3L1u1qBhxkGcXhhvfuwiVhm6tWEyvvbdLfCVedPTKQz7nCJhEcQdoX+bva5Zxg
XGjiLMxszM1O0IbmJ94tW0eUmKZjHNgPGeZ5VbGsM+KxQ7HDhxiCxHwOe7wm2u0z
yM2LW/xFN3gGl0rCZohE1a2C9k69it3/HkdgDxVtN5QyThkuhqJKnSmAzJB5SRSA
4CetUfAiTcLgVs3qEN1VYzkYuooqketbhtuXoxLX5CdLDNanAk8ej74LxT/p4Ma8
r1g6cTrWN5GaSdpHGf0E5X8R66WEFsPd/GZ4XDMA2jMNN5TmXbM7DNzrIqJrz3OZ
W5eZydbIYqBwvWcY1V9/SYproWzYw6GZ+t28Gdvqrm338n7B2Lk8SiAxWVGT1+4K
s6MhdD25XggBrjt6p/CNpxwYXOePXJUfTtAo+RfC6rwHmsdfyMVi+SqoKV2fBtKx
W/F1lvnYFbfexBK0d5NVuleMG5bfpXJRoBvceAqMJ91z4bLBjTOChSE+kU0lmth/
dhBIoJbaVIlvtgvNi4erHXyXnBaQpYfOWJ1v/Gjttc9hmb7L5VmjfSUxxGYn3hJv
uKnB3delOnc96pA575eHo+PUUy89SUOMjhWM49CuIFIMO5Y0Lge7JdnC6jEe1crA
RhqZefL8UJu7G8goEN95JRgjYlmAXKLtupK5aveAJ18Hg9qBQ9+PUxHSVq6DJEZW
OBOgNPvhvjP9P5kanCYxpGqxNDTQRcAlDV8hoMxqGLgWx/4hdSGFe0X6cGxmmJyn
6N0WtaEJO1mmQpYfGyvPJZeo5b0M7rGTfh363Dlcjw9zfHDmsuq9mSffTeOQufBZ
dGBIMd7EmJ4I7IPUzhhYstiUyOA4J8kNMN9Wt1gCPuwE0hbrlAhI4pcmMrJuOkuR
6FX2b9Pd3NKwYZThdCbg3+er9JLlpZcFK7XX0TQhpkU38ESj1IgyVgKAkH3x5lEd
X5sdhAhWMWZOuEES7qG3WwNwYquk3U3ImVXh9TaBvv6DphN9IjRKj5/BNamqIgs5
nuMf9XTYDpDYTCrLLV9gH4N9I0gIgXB3g1bms8weZYgwAMqo5rGx2fZzy9+rms5G
wq0GE0XVFjWepmmreZpd831EpUJkcYEK8TKi9Hzgn4vM0u6pV0YH7lvoMm3NZWK3
6Jba3nwBka5Qaf1wUdkXsBZCafEMOckIgQg5If5wMysu70+7tiXDH3bz7DZ5P93P
4wA1cucYqfr7NsiFR+VphtkRTx5SAMu/T6gyrjAX9L3TfyB4pFNw2gReQaN9G5fX
VdiZsujENMEp0xbiljpcHdyQLalSp908etD3JM7h+Cd8YD5vWkcU4NCFLNFdCAEG
gJcWoLebX6Iiw+lMUYWPtSoKFmIhazzO/157++6SW79wYtRT7dFs8vlM3hm2Eenr
sdOgZcF/uokzH6c/Mxsha7J81r7Yncuel9eKVpZYsiyqK4I/CG3jL/k14v0lk5cd
e12s6R9bZ8AZ/iOe/pUAkw3G+JphaC4ARELk7vI8LKKSh8CqvZskqegvy0IeYTsU
pAfe/+k67Trp6ghx9Z8RzKIqFi4feCzypCJKkWESI7XLMhkt2yzETwPWZ32hWgoj
JUBJNLVL1+52/sjf9alJ5/fkWeHsfROa1bYbpRkq0hCpG6wcPd0mRgWfQVWPj2yT
MnKbV57uuMPQv5kTdnDtMQrWG2rnDeqZE3+xl1IREZxAO11+AmzI8/U9JAlWReQu
KjhShloGZQ5ZzmtbgHm4UFR9ypP/zrNhIk83Sh63f0BAenarCbwBGIHeGyKT42IH
KR6jrnvK5mP+ewOJFx10zgVMdifUMKJeqeoOotlgF2qZSVFBblyR0WRP+gemUaGV
q1TOmrd09riA9wv3xd32qiiUKgzycv+mMeQQP+bf+bHLNOIXMFsHI5BSLFEi0Cq7
g0p543ZxwGpTImUDhzue7Jq4ADiC+vOU0OD4Yp7mqY8qYZljlCatIvTYXmf+b3wo
T60TGIm5FGzNULM7y4COE5HpbV38nAfOubtcx3dkGRbq8m+s4Jo+fXH7gRF/QTyq
rU0AsmIUMmZwjvg6yp1zMHA6rTGXTkEh9/OA9OjTSzAamZFAtXy1wfSgAqzx3mxQ
mnhaYZOfI6vO0iZFaV4h9SHwZ8chGobKYzvkdd4XPYtm5trgnx+NyS13kZ/inbwn
1HjcLP5a/Zw229ghQeOOAUll/QBBFPuiYJVmrKcI3jZP+BhTgaVwgiqE+hbr+gnw
eRgGv2a8z1jpm84ycQUvHPRm+i6FZd863iobLTWUBHUPwbVEq7C+Y3sNx3iyPUv5
5xXHe/SJ4Qy9kWLaYaJ9mJ8+7iIOszdQufiAytFfJVESweB3ijairBTsj1d3Sbfw
RejPeur/5bgHqrMp4HzpkpmZNJLIJF5NP1dyizzNHe6TLEf0k+g5rNQRzLQ643Uw
d7gskKn5J/3DxzTkqG30VDCQ4LD7X8uAxbXPu0IWq04Yeq1zvQtr2NLjNwyO3BtY
8CkmlA7jftL6Yx4jPQZiFlpN7C6nq5EXN1hCCJ0Cofo5/qW/Jb7IV/s9+lgErBMF
HlOiDvCyrnH/jIjVb4MijQU0VPxjL8NPZXnyxIanH0ryy3CjwOLX03S5ruBI7rXi
TLfAIhmmtbwb3Dlb3YY6myM/ES79XbqA/oKz9O1cKFAIrDtxJ/TRBBOelPJXVj7N
SI0L0rmv9Ss5QJ50vmRO5UJ/ZYP8zGdANt5hSQv/4Mk1oWsOemGs85csxGRhJ9oB
w9aEgcqHxbpGP93thZgpnYvCEVJumYV1eRS5oGvJS6FSQdq6+COBWa8z4mQJX2uM
Pqedpjj8swD6LX01lIeBVbs7aO6wzNXBH5SzdNYFQiSeBV33+fRywYIrvN/pjPXJ
vl7T10qaeGqQ2C8CJnTbt6/WNCEIYk+wF6yN8ydGtqjXC93YWgKG3IF9XMS5ZhwB
5g5iT9tzF+uNgATRF2KTgwGTsgs2AfPr6nzlRclIdtReSIH7/77UWwSLdJlvvatX
UxE2spSnqzGYlCBfkxqF/YCBMZ5t9UZ2np1nTvBG4bnakHl6jsBQXGtuf7BuFTn8
OjO/b5isM2a/CJkw9Qfh5umKI7uVBCLwnMgt+z+VlFmFTTjGgu7TZ6ftZRF8Zzap
wy3eB22W3RixbpWL1mWABLE4PjsggI0e8sofvTIfOeAcey9HqJhwB40UJbhFL2kD
i7kaHrxbCmdOZl+OEWMLDBPwBEzMFAu1qsDS0qhvE4LPgGdf3mAJ3THflMgoV6zu
WB5yPlP77dgcqtSQkswHLSKf0HqWTSPyvmL2C5ntNPKKUt24Gly5I1HvSVQGahvB
xRn7e9ICISHGMUNT6LC9M6RqIMWy4/0GoCZXss7xlrSnhv4jO3gomJJUfQJpXa27
GPuCkFDWrULIXXmhkUGdJHm34UMq/qy6DjGtJzWush/HVYEkht2VJbb+aAxNNwU8
7PepvmP0X2gbcT/6fipRWbzqMCeAdeP+4F2CX/0eXaumevPumI3so/5PZYk6PmdY
9djqxDfScGHOdE8L5+jnwJjVxcj8oxCaCdPT/HFk4n8FoAfVve85n3pPS3edfFsS
dJHS/bbbehGg80tm6ts/K5RT97WEZFNuNOAxi3dJtGPsHJ+qw3v1Db2cqnD4EjC5
if2m3wsKMtlmuSgzMEcXRPKCL4TfQRU0AeGsiCgpjFTxfqCPCsV+xDJU/g5ssYiy
V4QMYs0XV1yuZn1zendYSXImcQTD6Ab7LOE2hzF6hBM8+Rc3nLPoRx3zj+Fuptrc
KjZxIcRyLlrl+qukQst5mXrzPj8uzl87/QVtdF8M+VOUkO1ZetwLpM/J5gJHs0ws
4em/vzH4gPIpvt/b8yeywJhH3tnylg+7Y5GCQ3C0ayrZ4YqF1HDER3PGHS/FaDnF
5h2I+n3iI6Xu6Wx8Haj/hUYNvU49dNDzdq0vrc0i5Td0ohuzF9U7Gqk8enQ1HFRs
QOPO666G3yCpvujsTY0H8icx/n6ABd3YAtlezEZd+QJ55VQ9YcExsxPUlT5ONHhW
jWF5anOoONdsfNQw4705v/Z823kxHFrHEeK3YKS6GzUAF559ZILAUexf4nYL3cUa
nTuzBcgmNpOYyFTCqGEgjyu2Kk7acgwPsZQiuv14LWeNPx9nkb1Pf71EDcUJ5+Qr
YNQPCqHZLEYyZyP8LcHltdnnappNkGJzVOcTA8ccWTCB2y3LvqWiPKiINeADdW4y
Y2FWsUgxVcMr2jGMMvwLzxoaMKKBH+qbpmyJcw14VnBpQF0zM2vadFjk325m7jql
NCy0BGgPt8obH10Luy6MgZjkWY5x9813WVopVKJ7oNo8H3/xkVewBDI4ETTr/3Sa
PyF0UYE+0KiNQaD7rYXXy5EggqtjWi5SQIabQ8ILRn7q8R+fhFagzsBhviU+gT6M
rj9c3b4La2J+c5HQez8UpH88H4wfiIMTLAIyjKET5pZtE/tdbueudHXUorNGiag4
K6rmHii8SvIpECkJpyJmLv9XHIRIdzuh2RRGoD0dz1zTR5JxYzccvxFH8rW5cPSs
sZS6Hz/gQAZIkboiPORw5iWZjabRgNnnMGrKWjHtaAQDc7cUUMhtuKFUlfEowSHr
JLsgMTQd9DL2MrWZ0MScJ4a9FxyweUH/ZspI0Wo5VDphUOIkACH+Mlm3ez45Lle2
RPb/nL2txsn77sQtS+uVcIurPrnbOmAUPl4cSqLLPbdUQCk7L2fghb/sTBM1TBZO
KOaSswklV5+NGYtu4sZM+bb5sfrqH7adjo0FiTALfTT8Ew+BHr8aT2idED8sUdQu
uP66jzm+aNolq6WlxNJjzeS5m9O64Ph6FmpkvjRVUzRyHZVqucsbOvxqymou6UNL
YQu5d6rH/xV7nzneLn4CjnyBXtDvNFHuiYZVfSfFtKs15ocU1KWjOXEV3nQuk0qV
1KDK8dXT/hckU8IBoTiTtxXQ5VabMxVCoZA3YKYjXPWptJmTiMVfRD7VOsJu8yvI
sk1B+MCdde9eHOTac04KSjR5dwQ4pF8EBLt9PBeRy4JY3rjRhfN3fU05UJghsQDW
BiiI4/XcNjcXXMIgI7CaJhXwrqUlrYcvhoJQ33TG8f5IoiGvbCq5YiYqdk7g1ZI/
CDBz9jpKww/M4a7TeDL91jmp4aNLowL+5jrCQ4Cp2UtKK1UC1QE9qrgcdJsBYL19
KXMjGaJgSRlc5C7kvdD1UKkDjtUrw54lJQ4zTz2r0QTHmv4BeJFgOTiACMhGUtBI
sBGwDpeyxJpbcJgqS8lifd7Tr+vQOu3wQbXTk1lOfv94WEYk8sWcoRsSLpBDd93Q
uPmPiOGN0RwIlt/l+of6psOoN9InzAJc+V2Fd+/OS9ej37tYD5ZeVpQ3hByIZjlG
v64LXbFCXaysRMZrgHu00ZdJ7tQsYAJmSVXDh8grkWGfpYdhsSzMQhDQGSz+8Tor
AyXg171MmhryHH8aGw/0nsEJPi9BBjjd+UcrwpwF+1NZImqEGR+WsxLo/M2b+qNZ
82sHbnek3vs0/XD607c1IYc1XGDC5VGdbcKUfJfOyuhhV1k/4xSgyBmgAAG3lq+I
3eHcQ7hu+OSy/eBBMzr4b48iQiQSgRWhgRFiRUCZ1GkgowGlOBg/SkonxPtAskd2
Zq+1MkGRkFiMH6b40BcH8G1E58Nnwn/oEyfO7AugJup5x6kFPwBHOfco7uHdutKh
wTYZ6z0Fx6NbBUjjYv3P36wL0uG8RwFdYMQnigAdb4sohrQ14xJqd1NH98tHFTJu
QxSF6+Ck/70A/KwntpKfoUF9CwYU6rHmL9NZfOkzDBCpgAaHGcAwj8uN1dvCqQM/
p6pMIUGvm79XCNz8HVMmsJfDcvliOcf2Qw4HrycCXHDc227z6rciUPdeelzUwln0
babU31zQyqgFEvadwP/NE8mpd53SCbUR7gZfmvIQ/773+UQw3/65osLV9MPCgvS+
r1JBfMJA6+R2lynDLLUQm3l0H9CzBd5zdTQaRDyQYllYG3OaanaMkd26z9kW8FwP
9DAfeVDpNXsgAWKWOxTODU7rGYJ8V3W14FSuWatwlGgU4GI7nlNf/MfIxnrvsHoG
CgkmufxKfaty2wCTgBVU2ahoyn5RakOa2O43/z4AeMGRnbomg6xagd20mLMN7Ic1
6GVznkLC5O1R80uJLSFmhVrtS6um+k4FkZSidqQszDuY4JMDcQYybYz3vfAUXte5
ApophIFKjP5sXxa9fGsctfU639Q/LpdAdPYqoyQdtxnI+S7vvN/yAin8QSt94E9k
Pk3TruK6fJUKeFhwOpIFfh2qG+CrjQPTbp2buxb0NqhZSNrlUZs4WTeUQ9QoY/9u
hmmzG2zl7mJaN6RCSaWWX0R3baLjt2AhFKEDV3CxctsbvdV7D3BrHn5rYJZAdaMA
W6Z1mJjkcHN5l8EIhsKBhoYsTZEsVpK5hiTcKnNmbu2XDbiTfkJinYcwuzrtBEpn
r9tY02e5Mrwf4Rk2Fow0pNy6CPzNGpduHZ5CG+FA0G28YIh0cA4jBDA49YIAuQPm
hIkHZC7j45HL1JcsPQUOVdEWPgY5oOM+zwb0Uo+HeaaNIqsRt3GKI6Rg1bn8Vyog
RcYSdOBJF6HvlEiYt+OM2j0egTa20lvW4tdQwXn0gwX4cZFGyco5ESx1WVWO+X8k
nv+3ZGHrhc8xILBcHnlVOKwCabYCBBrbW1DjvMGYGmfxXZbMYOGPoTjrH35eugyF
EqiyXelyXbN29H4s9+n4Xc4bzet2V/ViNEoaBzM2/QfbpBE7xmppy43/t8rm7cCk
YQrvdIlxKqb2xLmKlILBGiMTTlgp3CZ83wafeguMo3mpQhqWqTPs6Yh3BeG0XJyx
AbL2iDAlrlR5er1BMG8gG6BKG6dXdoXZhd0HP3m11dka56RnzqLug5CiFoNo0Lz6
Z8ugYIDBeGDBGAQQecKQu2YP8ndR4qkUQka4AzAsxTOjESLWaV45knoEbrK/5K5V
2mzHpwOy+rXXFO8PBZDrTd1GWMJemlpK/BGH1uoISkhgYpAkRsQnzqIXp0rkE3Dz
CYYLzzREnpfHq37BJt+j4KMcC3YyYYYnti77RYUAHO7t4fdytGxvrOl+OPDwVdKF
d+HoAjOGNrWA6bXnJA6k4nj8I27bUuENAagDdMemJwbanP57ZVjCxvpY4o0XRhO1
SJNrnn5igiQNRuEkUvZyjD8S8VND410H8G8g4OyHsHtdTPmy049PGX0BEjfpdKon
PdPyWxafPCuo2VfaXqxwfY33kLII/7KOp5miB7qXCr26L7SKKA8A+3LD4d+q1Dbb
YXto2YCaRA66NkXscu63Kz3p91cf1CO4c3QS5YjoGW2LZxUENSITkNVnQkobt5A1
xDqNbBmrq/YDVpBRHm+CGo7rws3FS8PaC4WeUgvxsIi2WeTF8/DvTyTcZjBDGaIS
NYnouK/nwdEJbojsPutbXIIfQOsyku7MOu5PGFMato526FPw6K3b1+Igx9b2AWYY
5+AAo+HUoGVWTDLfOOyA8wQROHBCreiCMz4LLSmtpghPrMrgZGi3z1LFGK/pS0xT
duRs4W6d6EPYybviGYJf0R70ai+AE4ur4IGN0FRvn41gwg6/wZq9ru/QX/knMTEH
tYbheD7hu4UTEWY8j+Bd/CKeOSqhwKgAAaVD1DDNrhSz2yVr9cxwX4YBXtZ17s/d
6/USB+Dsf00kTTz/PSDdlYeTcr0sNRbqRZFEMcx+Cr5q2f7PdbIaAYX7Ot7lvIr2
5noW/OepI2dGmSqZKRm+saUwhGwStx116Mcjk4KTIIdbJiXxOTmVcaetd3Vu6c1R
hsCUYz4ydK8bIWAymFOr3h2YNeaGokwJYr5qjiOKqgTzWg2BQ6vatGupJMO+oXTb
OvcOAnrBr9P/EhXqus7CmmFqFJLpidycHRESdnq1ocBILmA9sPYbPVe+oZCZkCiQ
Pb3tEqyZ5yKZ8AWeewvDWPUcmukBBVoeQJfwTc6sKGw5TZHk95YuPeWaMIRIO32W
Hg0ndhCG9sLxbPTlijMTHxVkCEd8jJnALZ478UydlqekKM8r2QeP8qeYtp90qgnh
x6FytgL20udar+NXMVGIZP0PnTkfEcxAeHp8lRsLELRmz3/op60PZjzKWOTNWKU8
SepqTpGM3mY/sUgRRDTs/nLS09pfBX5CI7nSR+uEeqLqlHhgTtLJRoFZ0L8k8MjP
T0wmofZlohJ4+a1moTAgc0UoYiyRuxy1f7u1vxKD+/cEB6U+HRkCsz/UipbarIhu
0/XZTTIFfcUpe+r2+IbMXfo3iM/tE6q4ZW70yauNUb+93fCItx/Nd9lr0Ou1Dxwp
Tr4yCd3wYnFYPJ1eNMvthH5rJGYQ2FLD+E6dLnwju9UehK3F16NHpU83tFvoQlv5
HrpUDObPRMsCtBVE02yBiYTkcZ6kPwfBPvDa1rYlydbdnbZdX0HWL4SPxqNI+cNv
rBVaSxPhdgF+Spdp4E3dFCjn5n8S7SB2M3MarBn5ohsqmqbcewYHa1/PPNpBotBv
XtW34MGms5ZGRUQd7rec4qgFRNV27rh37HC1cgBI35qouKRO8HGm46mA5ERNqcjQ
z0imF3bqDhzVqSI0BjT7NNhVHAWZ/XNGDIkE98d/2/BJAN+4RTAqqDdo+TsuJgd8
moxBwcFCLLJm4PY9tbZel+k4GqEC5xGPxhi+bfyms38hQIMuD3QRNtpz1OgBRtcH
/6sQ3kHTclRjrAg7y9Zdfi7mh9WdIILfdoUmy9f6Q804THNnqhveMPX+blj0Z0WH
YEvNfigx7+GWsg8Cy7VrHvRBMnbGUCyGGByW4FWsvMt+hY2dDcXBj9FcyEbb1sTz
n/sb7+XHRB+ybjkwZc3Q3UNckjXfZyMYwnSD39iROu8s6XECPNF/GsHPe5C7b3vS
2UqByZPv4m8KjKJkZ80wyqAY7DQ3jp2rKavRRWKBIRKLp+3uL2/tDqKV1OwRbCln
TclXPZWH0Oo1Bjd3ZtcUiXYxVSI5Ty+CCQyCM8mGHtoKsykD5drMd/9oX/PKFV/Q
iELC2klP1NdVzzbM7uMouIpajj2TRfkqHXt7Y7CzN6tAzwssnxbkZT5v4FwraTVW
7Ib20BsQo0lMQQskohBjW1IK9kMwzrmUsnHT9YIyxomFAHMyo5giIonrwkIWnLjb
SOYOEthwTdqy0TE7FJp5U6tNiMMpOHZVmudSeoQ4P4gA0y5YZozzTcXH1KczOq66
h1QuVJzvslDuILg1nPJSZbitB72cJVoF7b7JV0YQn+OLg8iplozc7ExT4eFTebpc
t66phG7yYz4cIaYALqqYK+PEqBNl8xOIaVAG32oVaYoFF7iHUOrnUubjVgnrz3P8
x6JA0nEknVhsttMRO7ncd3zU3xt6QSAaufWFcIruKYLO2wkmU69PV66uSPdj1SYd
tif2LZchin5efu3O0sZfhcgT0yscYdXwaPQ5wpWSDB/MN6BJDD+39VmmHWM2NQWL
TOpa6BHwd0/pjhaZlIBe5lFCyEhDMRAgp+bs+E1atS7Us0fwTKcjwStadL9Mnhqp
pfMBpsue8zY+glPeI+sgSDL+Wccq9hM1WpfRGCOVRFbTC/NshBrb3Y+GuEJc1xCC
lTKB2jkf+nA/a8++9qtNShikwGbK5UISFbvj0hlBLFE8rQz6hax9ZIsZH+TW7ox+
u4qHaEWLpg+T6/P/DqCgyfBNUlDaIqfeM0UuFKY8BcARf5j69yFzPmvtinwFzAiA
Z8bKxI0pNnQMbPmgHHEDeL471RzO3OYkGSinVAI9tF1TNw91P4c0gMeZkpwSuBbM
UfLJP3QMycgOUa34zqR/Xqz1GpcfD5yEHV1YLvHmIhFyG86oUkllol0Y4e1fpXG3
1ZLgjghDZ85PSY+JdAPpsnH5mlP/aPZlvChoVolPrglvWx3x4U3qW/c5b4svjhfW
dt3oID7ioi9gV2rAehQ9kSvMpLov4/K3mnxSOj7scl8S7NibDD4F77+QBKkTH+mv
E0/GQ/g4xVKUYcDp4w2zeRTn01F2ec4ZslKNG0+oLyfGIp0G2+Hnx8lCDKh+h9R5
SjBcjoHbk2gVA3gWadNvg15DgU4qL8VlgsFQ+4QKVLxnY11gXdFMrM8uPomvHyg9
It+/YGAMkDvPC+/v7pZHbpvEfnjAkJnlPmgf95M8UzzDGok9UeMpFfwtNpR8RE67
dUdImYlLvKAdNjO2YdWIhBVbOoRk0/fkA9q5kJxZfvK2CzQrWrpZB5yNJVrqcTE+
xNRi3APBbVtSafSUbvFfxAnVufACXhwMCBrSzt0V995cQlKoYGo+Ajb8WOL8I+oZ
mtt33tdG1TfHjGszFxKdBO+uVRzlO8e3ATYcjPm2sP4tpY/JwfDID/+DGSW1HOmv
wPg/ckMyrUFBDIP0ml4Pgeb3D7WNkjaEUVHXnnBFW+U11u4tg7L2Nqms4Z89X0UV
/2h6MbEnPXz+0MFIeldco8sngp0GyqotP2DYHEuA6dPbWtHw9ZNZOuj45zQqff23
Vk4ANbLy3oD33xbby7tyLyCUZCCwVlc7uCJGukxWjnnB9l9FjYlTMNBrvmNDFqCk
HHL1PCDHN7fD2SpMJOqWUPZJhSQbWGfTirZfNmo5ZE+oMWRmF12qoOhTMMyYSzCq
N5bjvRtg0uaB5yh48rvOv5iS4ngWMJ7EvyjNJwQdKsNELwC/9SzO22wLGngc7MmH
tg3K5NK7eWXYw9ErzSn15J1+Gk81G7QcCDtSWPgz2lZ+TaZsZxGyw+NBLeoUfKcs
cJODT9hJGRzNJbY7jzsIu8ycIicarzo52cDRWyRwP4Kl/o8BOQQE0b2IOV8+TTIR
c7z2WXWVBkBmsL8/x4QCX7xgiKUPQt/uJusGGC/DX3YaiQ7ZM+hi9c57Huerleuf
Bo0ScbdA3x6wYNFO3OvymJnr2PBr4GV+1kdu2/0+23MrZOkoeLCfj4da9dA5hBo/
02EBR4p+5lO0/ecwlf1HV+VMvomIz+yqzWsoxpqEyeD08HTLpTdZ4iNbySaSucZR
W0o+gndWT9xdjH9wupsPe+0fT6YOFPyRsWzxiLQeIYAYl76BJD6mtsKIGva03Ish
PUnhRHLXR9+gdpoMe3gmB6ehfUS7HOqMezmnZK5sNJ147xBaj1uz2LhoqkR2kXiH
uozrQTOEEyYMogio4BU7UnZKbCEQ0BENHaPxwmUZ7Tj9z57GO9EdFb/LdmMe4szT
1HvFN6gN6M5REy7pni44lPleRZm5jk/4lepB4/4RZz/CPVyx5SDafXclLcOGeuTp
zVEyGvfkIe/pyaRo67ITWtdMCSqZQW02TEXsm3Ys27HfslbMF6RtZq4q72uTX0da
UWuuARdYJi7XeV6v6p5x8OjMy6z+SsF25B3VGyQzYgjzmOtq6eh6g3Sa4arlQR2+
bK3z03xWSxxVhdm+LYUjKom5g6jjxs3whyYFJO79zohRIfMjh7lQ4UCWkXqX5vJF
Rclzis/PJbDey6xfaGSqSKPwJG466u6eQ+1d6VUc0Y37HSpmPnvXZNDIFyyxr+2J
fG9k6DfVxRxwlNQ8prxAB+jQZtyqOQkguzziGdIcK6uxszoRep23GFy/jApWnuaC
NeRKZhIMzZMoGo3N0V4dCHWB3kCyL833BoE4r/o9Dv+j6ej4a9vZ6my3km7iYoRG
0GLaiyb+ILr3xJFPVRrXy5lzNCYk/9e/nQQdSmW4Cs3dMdk0YLw9AePIzM8FvdH2
C+OpkOJB13NbIMfuLTTvEcsJ3EPegJreVpMqBP9kGQj4O/ovlMcSj/a5uG5LlxEu
R8Gl0txnfvov07KISC4Y3GsLHNz8CeflHi3j9LXV8HFgx9bs2BFPbvSga7lNk1BI
lr1xv2jvRrHP2YFlJvvHNM48RnS/XrmNSAEe8QbbJ+/81/dS2WXNhlixOGWr4QW7
NEcnXFZT7FR8EROQtLKEVEFniqYr99uhKx6Vw6OtnS5jeaEaSe/t+zaqETrY/fMZ
4swuXJL8drOBJ6d3QeD8908nd26gQbMRZ9blSLII2sq9NuZaKXGcaq2MmcHdJzR1
MIH+r0sZnW+BJQAs/EUds41J3RCAojnd3HYlF5/KTzWCph0NeZVzLULEXJZyeygL
QmMJlD+Zc3y5EYloLEmxJLqFwEquSiypfZSxsRh84uMQTIpEAmaCSdV7Xvy9wu9K
3OuWogFYW0srgSgq+3DnkgG1j16FhLVHZoVZwFC+XYbT/x4J/ykBvM0rtfBKiJq8
pg+qpJuhfqEhFgSsCXd0cFd+duldOqphdbBBxomp+mZ/Rh48p1GppYeFzR2RPIMY
VCgh5b0mo1ferMQfaclXs5p9lDve8BmjauQzTPg768xzxAFsnKBeh1zgoZnfny1s
NdEXGF01Qk+MxzDayoS7KLJCKY9KyXdGdSP+ZMmw76IYsW5R7hg/Y/Z7VJnafQdT
e+r42IaVXap8kg6ASMr0sYvc7yO2jWXf76keVCQmHKm0Nniuvs3DnvMVSauJ4PBU
3JWKFKpM49D/4xkHaweIg+Bao2AiZJkDE1XempB0Cb1f+qAiCicRgtlDkGhwAwFb
xfgEBuFMBNC+rJTy2D/IcJEBRXnm3SIWr5QXeJJGlDwcUTRrtmlF9nLNQD+UlV4u
u83uxRUaJ8U9YDp/xCVB1pb6EgJLpTgV9VjLEjq/zo7zOhBG0TFN+33Ir8+lADY7
LtDayuopwcx8zYKZpVuEQj2KEnTatb6226aMP13YyuCYj0rFKDfo2g6uLLiuh6Je
MDGoT7ivq30FCjvqhi+tT2TlZpFa5m0HM+3i27yE23wg+u/WprUBPj0I1q/wYMcv
jcDoMoq3MosisVTY3sqwisIaMl/VD8F+I5MaXgHp9XhkAYTsq/8KVa9Mgi7617Xn
/safEJPe4VJY/OMSCa2V9i8nQP90IZT41/y9jLOhUtUxEdc1pcuxD5Wvu8qojGdU
yU9pJgj0PWhsDXiB2Pdwe16jZfc1Mhix3CtFtBnFNf0iU9LREpifRR86H1NJ8ZPn
2RybeuTc2XQcerv2DNX8LBx65uM0Z5vO13XMflKxu2bDtxoToKYkaIgh0EW/8UE9
Lwds3yW1POP2eUzrxgUZrHBXvJUYUA+0M4gmsrPlTp07rV2B/DE20e4WEPKvaE7J
Hg0EAToBOSU+gtgCsMw6GVW5mBv+hRbANCh3Dqr/2NDm5k6/daNZ56CGqvyLw9PT
fItblgVDO9UyF3EFXKXpcqCu6T1YHpmcMSMQbGsZp1pFWfRaKYlT2NRhlNRd2h1l
TOEc2d7YIpR19/fLpdUzn6aKT0WejFl96FTamDzBpCaHfQOzyG+y15T8W8PDGw8G
n+WQDg7F6RgyS9Pb8TvlHtnco+V0ltlsNML9Hq5Q8ugm3NNhj+5/MmApXT4IjoeX
CyR4YIvI9G+GbASmZfkK4FxFc/Z/grZVlcCw4OfEQZ9ToMjJqyCFs80E/qwGrZLy
1OX/AaVJ5JrUevaRCG9Dj/TdvbhUu1c+mmF2zftTvTFnwhfycIJ8gBYBtSJ3mne7
d+5ww4iUK8PuyMIOtHeuojZAcTxLga0AyubMbkP581yXAnSOzUuxRDocZbq/WkJK
PmSxfqsBdarIA8Hm+MIOEHEk+rfd6XwKARCy1UARMqdMlov/0eiyFb1yyMIFjTvw
f3p+TlI/3nU0dX1nPHst70znlJiY4eaS3VbLXzg+E7R7VCTp1+UTi+Af9uESGeNS
2Rky40NM7eJxc/5Ota9wl4ZETrNK0pLzzwlCVTUy3s0HyVofstWIWONGTUXpk5b6
uNrT7YkXjbOGLusu8ANsdEQHYsAKvxcSONKYdZ4xD2B3q0iyXqD4ukm8gE2VrI1o
IkXBryd92v6FM0dl+mO5iQfhBOwyIw6XnD+lXMbjgA8vP5jIawkNfUC49pyLvnMK
z+XU7R0l+ZpifKZAxT6rJym39G9EQ3ucwQXQIBnUlU6SqUeA1qjQg4LrOx1khmBa
5DZa0mEHRC5y/MzvXPKBJLsy8iF/1a/VZ4Rb4ulZdRoe6Bi9kUwbRoI97huLnPnm
IqUj7rCxY+zAvB/DFMi7VShPvOAakhupNivQZbir9czPTXnzFfrxAnJsRYAWSa9k
dReEKrBWpALdd81IJoQwlBXpng3OANBxlWxz7w8jiXTvvg3VhQ5Id1OBM3fheV19
hjOtwlCXFmZfRQhgyh+vbzxWLKRRE8SKfIOKJ6LfXVHe7aJlQoDoAjhFYW8SZe15
1tdTuYGlCzQWY+Ye4HR32CgJL6iH2W6OUSsP6Mxp1qlaPURYRSdsGqGgBA6tGC3Y
V9b9d34+cIH1rAAEs80GIUFhMThSGb8/hXxZj8r/9fRSQX6CmShAY+imz7ztOB1P
meoowMWhriadIU/5zJxgSc9DBVGnmdNCvqrlrv/ZK075iI5vKIG/z3IdpKR95G1p
iZus6xY+xIySGc7FC/vUlu7duSgQ2KS6JDn0x2KStZXVbK+gxDTJIGw1mfA43KCy
OPLLex9SSLigUnpQRhdlQr7DpYxn9fEH3qAX712pji4k0ha759zkYVaqFTotoL8A
p59RNllt3vnpQqNx2FbnLrjUZV/2cJJ2P9IpH+4hAkvFtJ6LLeSnReiT3TmYojek
WaFwOBrSJoLMNdPMt6BzDEeLFVCpoqNsDUO/dZ0Ou0B6CbRrRxeKtIgPYvYWrtQz
AQ1B6MBrGhT+tlLmztfkMTJNIHzl2jILthHx+9KaOk7yp4A0DK62DQt23AxDVBU1
ogScKwxVZ9S8MSYmSmUDFKaQ9uLGo/9cgsExHbmvnRHG62bHGUs2dxUyhqvEocFr
O6zrlzQEd946OkZLXyvFJhQLSYvObbl5UqdNL5O52Tzqz2AsRm74l08SfdrZT8ZY
MzomfMTX7ESjGvlTnd8ff9Oef0drwY7Z2fiXZO2iDoX5uzVerb/GLcS5tdV32x6a
hrLpIeMdKVKx67s0T4s+ieIosYh9FPmu7qV3fbUoEV7h6bnf4U6QacYLWEC/MxZH
7grsDwKmp4484A5hZDDOQybAzYfT5A5LR/CLkHCf1Q5wM7QHLWP82NwCHGBos7H3
YDaAh4m3UvG5f832QdpcHFhCVIojHHz8NJZyt4SQ5uGk/CdeQfEy8tFvbNJ+KQ1t
jz5gzCcPOwD6VHPETqqY4ECFh6hfCZ9FzzzPzNleLeOD/KM2uOneK7lLbLbS/TOg
ERuX/Y5+tOWsIvAEGtDmD1AHqCux1McZiNQHBt0SSFS5vQwUFA55FRviTEzZ2P3R
zPCNPvhYZLf5Ar8Tgl2fEWVUZvHJ3Aol2yp3sis0plekb1JLEra/3FuSgYwiV43d
I19qKiUDwt2Faa05MQH+hkhrxXySH2sGAmMVtVIYE4YmwZImduLC5P4yAoPYrwd0
acKwrCrEewGqydSFygLiHOVoX64A2BSuGt8d3oOfG5Ie2Y2sLD0vwqSuKyDpfk0L
xSDHnlBOpnTs2MtXN2OaGEFWbO0XS/IM1iv2owS1odL/IUx/Wtb7J/recfi0JzPd
3O/rZvtr8XZZYNYsKs0f/e7S/NBPO2RC47An1OUdELL8OJSG9hE/m9pE4V1/Ijnf
6F/Y8EKDEVI+zZ6M3pCv8YCy7EbxBVY7h6K5/xvqjutq2lgsz2TDGhb6x8eNK+sc
SC/OaYH0T7CnfGGf2moUrNDzGaoVzqZpl+a6HSPbjoazBrzsB/0DgnI3XLuxMkjg
t9lYWQPy+TplEpdcKliXXwUiIOKsnWiikcXb4GqKbEJRWqvu2jjdVp0P+fb3R4ec
HbgfaYCISGZ6aNwq2MgFbT+0O6BevlllrSR9G65t1QdchrxJ9yIhsSJ3WfY2cv1R
AtNcasLV9oWly44OrGO7jX3Jwf5FuuR49RZJsM5JXnG+lCBdiQk4iuHTHMIMAFXD
1fIeJZDZLWD4oePucQnQ4ZiETEtX8r809Y1DXAoac0mmBsaFCeHOYN7tkplGgf07
VKE1x/LY9919xcCrtS5/221MMCtpeRR4Pciw0Cc/MzWvuVbxFsx01UhbOvF9A5r2
f3C66ZGTwTlqQ6mPetAFUQV2ud9xJKgPkFgaumEUfIiXq+seh2E1pJX96QC8VqqJ
CD5Z4d0VNSTVDj+ixjC53oQm6/4RjUJy24GVbZhtWU1RSxIPH8mQZYrWACShsB8A
E1Tfg2LAh7OU6W8jcM0t+NsxgoNiYtNeq1M81Ok1Bk1UHXTvlNbuvK5CXHbKn461
UavZUp7kRJPFEUOlwTeHuzqLd+CA7jU5XXxyPppV3DLP7HKopRVYYWdYN3AamBkO
a124Ly+dMh7r64zvAI0851CwRlZddL5+T03eo/HEXULxMAC+64PUKj0Dg1Y0eIEc
0vV6ehtJlz9aUVGIjTLOVTGdDxECwO+vP8aYV/yd5zAeBWFp0nN47l+G5ylJEqY8
7xEvHtdPtTHBlLlTsnvYebqtSg0bVM3cGplpPJrh9Aoq7A+VVvCa9/eKDq1CC+Hv
oRcfGHWgGmDjiEFnrsACVbkoY2f9v6Lsj5t2+UL72zDmlGb1gH+5f112NbDeueHT
9PT4c+pSGJHvvcIV+gfSAbsn8z2zgPMft34mPiJdeToH/cLfeP8fd7Mrpesd9mJk
Gt08Dnv2lqG08vpP+FDFk94m9DazWY51SbdsJro87u5/f12HBSAxJqWLVsZl9wZF
FUFG9W5O+rVP94Yj9yrilOHVa5O3GaJQwo49SfeEnfQ6aJagU91nABMRQnFZdx3q
s5tWVOzd8PwQoATVnEQkPLtY4MbEk3C/A0jGj8Lm6ofBG4ip7fioTMCWJXEZZQR4
SxUPQyv37lrrMF8fG+gS13vLlIPOpE773rnXsywCXp28OFiNTRcZ2NXVwWhaI3NH
HCnmmNd4IZyFGqgVnBtR1eWJOaz1P6a0yEFrGm83uctXzSUgIjJ4HBf0MPHbqH7q
2R2nsjFgpNtOsKOUGPeXy/0JuFirhq7a7o8t9XnwzGjMi0Loy66biMT5aM8pDfJZ
+S1NREGnippyeymvWITyNyc27kDUK5OjlKOvRGHCxlc0NABxeR7XQrPJEdmor2XW
DXqHL2TuqfsGVoN5U98nqyRuZkwqWRR2fzXFwcJbzBPp11huDA8lOdq0APOdrKxb
ur7Q+0PBtJtqgchb2oCOR9DmzTgbaOW1hoRO8ZdgvUU1JYjKs3Ii8o3N6yF/8xa9
bfA1MjaGRXzEwzn4nayj2GWIb77w2HqqydOJB29rkB1rispL+wYhiuD23GeiGrEt
wTaW5XWoRtYUqfZjSBJEeHwN8jWft9jPTFG6BVhyr7mCgxiLKgLnGnrwmIQvR0bx
JSTwQlj8PVlUKOzSHKbVYyNG7yyQplbc7Bb4HXWaPp83suVKerxd0jHng9qmF0gm
yoRwKeqnL9XWVdArLu2fiPIpU3A+2n8ZPUCWqqrUABrKkG8nLmjPZXosnJHLdnyW
BRsrmGsv/JhpQldmOSrC6d+TsmdBEoslV9PjYps+CNcaCV3kryqyRFyvrHp7JK8x
9KMgcXt2Q74yrjCVTo5NaGwdJqcBJT4HGj+dLM5tx5JiomN5a/n99/evgJkNC83K
3rFliQMAPrUoq4jggXVCBjfLfcbQXaBAKHBYTGu1VwLzIM8wEunuJhNFyPT3hQlB
W7+cY71jXg5UInsJvlsuLC/6zQpy7rSk5B96YEIgyB1qSy991UQfTpKSytJk/5WS
rLtJB13S94RaQ+frVTFPEuHjE3xZ4BTGHSeFUhatlh2eSk5GsqK3lCIxFiY2oRhE
h5I1CJL1d7USt3mBFepu0aY3FRHnThTA5wsb7Y3Lj4Pp+UKAVqd599A3c1W5D5br
4W/RvljD2TGt/2fP81zBqS0fmlwyuJVmvk/XedsZnUr1+CmYHpBclSd0CEZSO52+
66WfqaOFCMdFU9TSTPcSgd0ukmzgtREdgokPpLPy6wkJlGGuQHsxLh2pW5qbY5y/
qs1iHSEW8kDWS9IW1Lx2QNP3Xz4A22aUc19UuFmbdRZV0SIrs24iGRgxwbJDMJrj
NRIVheangqmKO4iBWah2yqnTNbpfLnplLKuelZu+y8KN9VWDUFBOLfGU+7iwklu8
P+KZk1xIt6PP0pdODP2e+iDCushpppUB/YGENzxIBS7xv4PnCs4Y9sy83SC6kir/
li0BLZYoIOLo9kXkKeigXnieVQ4oRtwfrlurkm/P6sPlCwuEjccGsV0dao3wb+i6
e4E+HkITLyFzPJECJGvkJEvTQKAUW+1I+fEVJ5K68dhdk2SxTvnwNVFjL63n/KD2
KNsEmVWJ7+6I9Zou+QNeN4rdq168XW55EdgG2QkqsCepTay7kY+r9CoorksTb8EZ
SRJx3BsLp7YFEaBJENWyMVjUjc7J8iH8xaVsRDPv5l/CV5tnbippPtJjDO6UmQfN
CWULSeQyhzcHvsR8m8nou6GfHVC8Ejj+TPbthHQjBQOATFIEjfb7YT0Yu9tvCIEg
Rd+HB5pz+POpDg0oIBZsTeoLr1g5D+VMXqSrzssWLhH4cN4Rq3gUU6rZjs+sUC8h
53kUOk5pmwEkS6ie0nbnFzSz8Rbufe//5w/Fy2jgD51mqGy6gU8a5qtFySHb+VvW
jcBbHA4IHJhV6mQcPcJN/EELYmbkfvjdQly6kv4h6i80IcoxZUflhPMPH8vmyRkN
20CK0NBz8us2me9YgKAHcvTiXPqyNBATy7PvZIByyQIQEeDkM3nAbK2lGcygkpRo
HNJBetPZjSkQksvytkLICfTGh4HJ0x9JFWQT8mOhSxKF6OIrUWHLxA2/NQ0SAYEY
TEh6g6CvV8iTABHsZhrwdFTUfv/6JxFIloUnY5KP3rBW/2XZerUK9XRJDzRm/F0u
WirtyMr+a/2JGlDO0eAV8/p2tSeMh0ryLmIT8id2MFJ1NZmjSm0j20iFmWeh+2gW
JDjuiQPyHpqjiZk1FzQiZsWvYIkBqh50/89M8NuDEqzzr3DozFFL1RPqiLu5fpRU
6ZNJFy3r8Fq1iFF+SDi37BnzEYhA7vWFX9aGiVi6aEt0LgYO78WyFs/+4yG9N51D
ElHeQo/pKuKjQ/E5FlndnEteUsAk0PFpPc7xruiwQVzgZgh0LeNmRW6POtDTudgZ
ATodAE2myP2WGQDe+IcY17t0MdvmLGkzVRftAsdXtJyQMZjjm1Oae00tADcgkvkI
pKDOpeEHMyY4xsGQJJgFgTCr0qpGF/VglpORXXpb4/v2FH8s0Z4d704osmmVUu0M
RdEs632fE8dmQYTDSldo7ASq9kXFk2NzKcNQWa48pUgMtRF/Qkm7ycGghUf4Nfld
k6s+fFJzQMxh6+SGJqmIDdFhoCcbXHQL6kJitR6x8b7VAX18epvCZPD9rvVtBgGI
46INPDnop3XkdMpY+osCjgDk+u7hVMv1OY0ifNY9RoKRzdFmR1KCvktVTuwwwJq0
YM+9dTj/DVUqdfw8sg9IXPpbujqKbqVditWp3K333kB8Z2ZlFk+KsO7fgs80fKJM
4Yxeg739NAEcjR3VHQBNbp4j0OYNhxgDvl51WYJTmgJSevUV9T4hv5OdSBgy3lWW
QnJrcJiQ4ur0JnkaRbJ9Ug9wk0zcLllf1Eq7o+znJkziGtz5agVoj6d55Iw0MyLY
USv22G2I5aOxR+uD+3rSSXLoUOvVfw+lVVMaIPB+9YVdsVCNITq1G7kFZKrXPKh+
1RpjnRm8w8Zb/DpORniE6HrKpvpWim2WYtriMm/jq5eM5ZSl0fqXGZt7IfL+z7wK
QcHcowl0Ac+dc+668zqC69PLhxQ6Ko5gf6/lyb7zV19x50usUYyoUCgKG+2IE8DB
dgR73C29jPCpP6sqbYTnPFZmzyOJl9QCmOc3n4cZ437C0biLaNAGIM9g7j37u1Hj
Qs+6l6o6eL4nMml0k1d4RF2E/pqeVv7kXP79aTT8py/hFpPcRSiN5VPSCTTEdKUT
sv7rEUVa5mnnt3iOo/wo9nSMzcmWB+RNIhpU6fkRsJ2IMjMJV0OjTXboSktn5FUt
+3jGCgmnTuVGW5VSJIbVw076+yAriBtWuh721SFuASZiE8XP9OK3b9Y23yq74P1f
iTk1PKsMaGke8fiZ7ueihvKn7XOUPH8qbp1NsDLZpRY93ErkPzgcUljd/AmpgABu
wWxKV20nFJ8zpoPCConuCa1QMKi7/10G5UWr7xRP9TecXHng3NhsnfxXMGDeCuGy
V1HCfyh9VeN7oam+OZqKaOrge46tli/OXKbMVr013UVJm4oH4vDuGhFtYlQjt1uP
Ri0arfAmpaw1PSx8cKcLhIZJIrNU1bQEy3idZYi6SKWFiLR/aWYwFAFKSqg0TstM
Nx6roLspjcTwA3HVfOUU6YWPbZzGOErZ5KB+eT6cnkK6QgvDznhgp0jDI8U5JL+W
yv/h9+ie79U9ORitit5XNcnVhI3VkH6wKLDPEL70/+gj8iCLf7HUUPU0f9Zc7Qln
SBMV5s9vtSONGpFe5da949Y5QjA6t9XSZFQkz3ik7ZEMQIcqhFQXcyEOmXOnhFXI
BpExN2jVEd84XqfUn0kShiL/OocQiCJTll5RQlih8TRrNVLygGqDh27LnYz+jRyJ
qJSdK8Z4wj/XWTJDXjfcEDHyVqOlNEDglcilNiztNpK5AlLQp7q592sQdWHhzy9S
i6Nx8CNOjzoHcIYu6X9K8hYnN2zTt6GWG9LCpLJ2OUGb2DQP4/6kRrj6vPy6FbjX
9oSpEYI4p4TLr0p9uzadqeKypCIf/T7Hzv2lZvfDeqU4x1D+ge9wO4ZOQL4w9rQ1
ogxKiwaS5tzA4JVrzjepxMR5RJUvzzaQ6+eRP0mQ6yWqm8fPLofkHcSPE7mGoN+G
c7C6ujn07Vxg7mhw7WSaKeYaLE35wr5HYIF/le4gadgnPAUWaIZGKr7lAR6+687g
HpqsUaEigRuSaFMvjlitO3eihgdXuhseeX4dBUi1TemjgklUiD6NXqBllz7V2ZW6
MjwcPu0UCG/toDK4yvDSNn5HGJAwH+BmZ76/dhizdXckGMxu3d+bBvMbpvcFvvuK
deJkXGn6bvALwz2SZALT8YbOAaudrxcPnNCVLppncYQw2G1Tu1adnU3LXkfBpWmc
kgkqbpb9nJJx0jgNUPYiEy05xBuDrYvLkOEEiy95V9/DXBaocOUrb4U8+H0do9BE
Ba8/m7KO2pEhdXR7PmQi8/6cBjM6qNA14DnmaXG7XIFxgFcbzT4pyt4Pkx9qnp5C
f9ExbWP3GRROMcFbYpc56Mce2RWRXvyokE+c3lmG6FAVStrOJhT3OUs6Mk33IN2q
BY18TKhGBrRNJo3GKaW7+TKBl9YBgtID1uO/7RgyHoExVmgJMsnjKZAiGemYLedE
COZCwW8DUs0kcBkffSvoGLjaSv9NgjtovBrXjxAYjpfZxk7L2KNwuYPh6otqqeI9
RypI+/4hDHSvjSybVL88cuQJeKCeI1fAMFGIVByKYqRZuJ90DZwJgjDp3CfCmlaf
1wH3zvVTI80p3VMrE9Olc9ok6BreyzQy8uC20uhynRCl3F+fiCVv1bKLkmDkJXNS
LlWIjD2ImYun8sRK6xAae07r+IJ0605cSVWpywCjNmhOz3PUCm85KgPOvvE0UHG0
L3kPvbe/oJlEL9N1vDerOkIzBlb+hpkC5BHWGcNbSynhhB4jIb63J03HvbzbfIDo
RNq1chbvMRaMVTmoZFsqfQLXECDZpNdwFPn0CNSimiDlA7axWFA4jl/rS3j1/08H
XpxR2aVRHIksJEyjQ0w5dhLYd1mh463add73bo4iKuNIY2GVBntZxSCiaJwCM9sc
3PFmjrzsiBrATLj2hCOKyef4hLFeunDu2NOFCsivHc9SLWvfnEZh/pAwNjB6RHHo
WWIzPZTdwMQL20kOWxryQuxehj7HMtFlqvkSQLc98gXwJQv4b8SGm4ohgSN0LdO0
k8Oqa/vme6DH9TXqIDHn8BAwvlCQt4zv6eaKlUjzc9PPycVKJOv2gSF8ow5ogLZJ
tbxypygJAdHNg3Adinvce9OoDW+9J6NA4VLAnyDfw72RwOuBGcGJXHz8iC5uBOIN
hgmkTNZKFlmM5uPxatr6Gew4dPtBVaGLpg5r0jAjLpwfacN8XOthGkQzMfgg1tUm
SVI17fwmq8lJRIL8upk6JdSIF4/wBZoPXI5+D+8axG5MSCbc6QsS3XznB5I0vXMo
HJWaRwOIeLgiLTEx6BlR6+C5ZXy/45NDqGrTnNGHMI3jaC4w9VR43RWD8xUvLR3b
s8+incf2OqWqBSEdg17k3GjG+BZrWhiASjc5Cwe5WTaLy6R2/8CLdh82/qQx/3Y+
3WNSQ9TGur7o74AdMP+hWQRtCkNRjhLzaYeoT545jjEawIhPzeHnENG2d0CBVWtF
kWwmdgjAaf5LU3Eu2KDcKYVvKwo1R/CLAngXR1gFKqcgw7g9keUZ/tINEpyqATrm
fKTa5Z7yeVdWGtuW56pLQNomf8v6q2INy08/IfS9oYAcD+4UhdN4QnOvq1CwRGQz
o4GJYCGFlKFJA9iWqNiLOvzuwdwtaSJX91ZnLQi1QLpwUx9uLuwa2gC+WjvIXW9y
4MegFg+UYULHzGYmDD6taRyIXsbbpFfJ1sH2plQSWrh+4hLRf35snfULqvck3U+T
oIA925WpV1hFlIwaotJKHsvsJGsk2OfAC34XFXzS3TWsqhx4sfS0yO4YUlsL7X6O
MXEyMQ2/VTGT9yetRpvaLjdaIoUVvbWUZzDL0d8JtGQSiLT8CYsRbejvTNaFTmVE
+NicwVg/+H6K94A7OjFuHAjJHsjSbY9jpSDZSnwkdzpBclM5DIEekOAgHel2imLL
Ra/wbOng8qsFs2KHj23mGoliBGmRMm0gJd6EBH0SCY7HJFoi6ZKS1PQcrO5iLSKh
dtwkEXA1Xy8GY6t0IPas6PCE38B3Wx8ZdomGTBLT7eveFH0kS3IsecEgQWQB5hN9
mvsMoNtpOvfPGgVC4ZYmsVU6fmhEoA+EGxr7UZc7oPUcTAr1w24+hKAUPRyW5HtD
F9ZAC+WgK4BTfdooEjZJnuqotIKDWBiJy7JULwGh+WW6J8Wgr5+8bqhCJ1c50C0I
KkA4JrsmoP4uL9rcYhmD7kt4C1MKW5RRP8KbbaimRP+FFl8u8Qkm5AVSD1bNweVL
1ngDwimFDwydlrzaUYeWciT3kh4VfqKIgJXzZkf66di+z/wCGzSoHROxybYyof0P
c63ekHdaJjzW3RxU4o2eN0rGMxtjK3RhP96aIzCxl/oIMDASHqAgt5LYJ0Ff9f5N
lgDDonUyK6N+p4qCNvLpBUgWmxG3wzZ6MtdNwJOGVE3IAvThC+3S8WH1MrrV/sod
L4ViPm3cpBa46Xw+Ip7n2wJfhBA+jsZS99uifhlXDyVz2mL7ZEXzL5CH+mkZud1S
SF6OiSu81JaprJNq4mRhS/30wH3i7DRAt4BqN0rjVf1I2UlAgi+znuaBzLaSz77R
kQ1pd1BA1ErIuArDJibt/+R26vgaQMLpLFx7PyoW/GUYy34fspqYp4Cc6mpucAHc
LeCxnP1VPYsy2qxtzIQFuKhXr5EUj+j5r7fbtnGBN776iL6ctYJ037HEinPQ/wrw
7eUFhP+nvzM7Pnp+3VbYp1B9G8bARGt+f4C0pP0F7W/br4RD3hRdAHSUr8yOS5UU
KcAZpgTr/Xttj/8JQljv3COkOCtrc4lgC3v2QxN5AcGYGpEcVgoEfK9/ueNY2cW/
Yt1YmQR916I16ZHy48B3zEZ8ijqsKWNKc0yd58Uxw7NO7PBPSKR2L9ASmYecxbkD
0uJ95guworqNi9BpUof+abp2b6dRgZVRBg2toF/s7JnhqTK6zDinEtFPuPOBmxzm
ETjlQeAMfSZXIa7CUI7yeakx2T4K7J69x1KJDHnrueEletbZVUwPsqv0DhMEzqGh
G4Q/D0uJuaMl9Lmz3zQZQs+qE8qB50nfhc+lZ5C288E9+9f1hLYUvmLCrG3Adcrr
chEMrAYSeFgq60MCJZzLe4vT5Tcq89jYsH+AjtEQMWCjIPU0Mm/vDbTvtr0O7VMr
pceCc7b8ru0ESAoesT7kcJfkKSuPR3Lx2oRNw1x67+Fr+sllYPymrQhs0x8qJQIs
OSrpHHKKkiZeQRoirZRgGrY/KZ6f6i3PxOCR1rwKtGcmnl7b1P/8qOl7Ta16ggiJ
cqeRXAFDz3vSGPMHrKsr5NNTcDrs/VC2p88qWUu2dSTvNTAQ+/eZDNFSdCGD0QEO
dfCTpz7nNSegJQqU0uKwFT8igsZpkBDllHfWap5IrMjjzU9HTggavHL6EAkfHAvQ
b3TCCJkeqoUbbfrd68b11u+VWlh9w0YuI6nFPOpYLrqOWIYGW5QeFSoBfoLnmJk1
TCdwO+DzWuTQy87AT4qSrJpSmo3h4ViLHbROHq9jsOU4SCI6Aw7BMud+LO8LUjK/
FeRn/wR0cHDLNYAprsvGETi/n+681+xAhIADKDUjMN6ekm9stDx8rjq9wwi19z0r
OV+X9kROCeBfZeyDjSe5v4a5OyA3/K2jCjFTQkSX8u09Ui6qaQX16DevkvyWPTEa
RMjjpODV6dBQrwnFUoGrKsdGde3ovFWXDZ+TvHtHFsYJ16MIw1Q5YV5qFMeaibxX
GjHurKgmJik17Bv7j7F4FsVjcdfYRf/71DO9kEpdhQQV1xLZwCx1XTQVFi0v3xu3
SBvhHKnb2UsE44b9WpnhWLjKBeBgK8Q5RqJdnaqejsH0+6baZh95y0ejSjsvRXeq
4qp/OWueccv3OGoKsbPIXGcDhF+r9UEYaTDOP+5lRrjOTvcLst+NKKwsgiq4+jPs
V/zvkvh1m+rsxJpIbtpx2Q7+U/2WvAFeIAykqnMan7T8RlF68TIPa5lVYsLyDk+f
Q7+01lj9X/oGhl7jWdIG7JP/+1I8h4fpKUaJoby/k1BMuxnKj/0W2e7nWsBTC+d3
oesIwlWW9zIAgJ0yWVv1/lgXsYqwX4FUQbK149cyf0z2+tXSRbUtSyfGNdzRxYIb
Xf/y8jnp72xR4UUxVzfiesfM9/yoQDlDhq5uaZaa8QxL8WCPgCd0STz+aneWzUfd
QliWMQDvKGGiCa//JxbC7pRB+bxhNM88DsX/kukINHk8RRE0rrNOoexSIBSIkhUq
irOolcz6RlYM3iJ0C+ScYD7R1Or8vYRlFLmoND5EiBBpfWXhGDqsQ0Mz0N4DL03D
zIlnKRaSFb4P4DNHzE0s7s0B04hj7WVxHcelBmCv1AgK3i0LOnQ4B7yuggGtsLaJ
alQD/6pm8GXURoQ2TXBFp2wgoe+M0TexF399t2AUWFI2rAANZnCTOGObvcY0Gb3v
5h8+svaPcNzmvyKLcwdUi2P8/iX03oM8DhFyrXntcGjer2zfHWqtGTjBdUa7LK3E
6YXD90xtEpJQmFCKeeWqKcp8f9Pv3KHdkkdDfUfxvVYFQergb2EaTh/8/RrYVyjO
JDL/1YDfVwScRSJcqMALPLBv6/bLb0wmMMWShr2UrTE34Ul2P5WIw6EUVWenEom9
KaltxO75w0YfehRxWatWBUN4Dh8KJ2QqDD25rXylWKZAOv3egdbNA1XznI0CEHOt
Mf1gCXuSQyVTY+WsP1y1DtElJ73iEnHnwkwb9vmUnGM5JD3YMq0IGKawwnxZPr+X
41wevYPpT0dEjtIfOiDRfgnJwi+cHkSTxrfyV2LUyZQKZ4XNcMdk/4lolXDsh0vP
CzyRBw0hMaSzFsYFUXluWIUeFmKVBmAKbsQ1kLap3OMuYAuB4bRUyWAG1R25/I+Z
pCaweS0rIVJ5iL9omFQ/zzDSce27CRrQVrG3vfA1UMW4wTA4ZDCI6tz+RSRZHdYp
8yf63e+NXXh/wL1GYifDxGpxRnOxG8SF/Qb7GyPlbQIGjyc1zQ/ZU0IkLloziksb
tMdP6p6qe1r2FjYyM7iX0YhVVjeJaiBR1DXPB2VFkJJLejzrgTYiJ++Dv44Cx+vG
92dcyoG1b/asgM2FQrLr8PYZoFWHYF//OkPee0R4y+IRWsyY/ejNSHyNBBT29qRy
iSaHAn3fSQT02gEV9HhSFPYRSB0hhiFSRJnUi8n+vihgyObk5XEsWx7YEaxjaulk
ivyTOJPEH6/IPwlyU28xlFlwFPYxxXLvPYyCiWqyvEiwjthBJPIhXhb6BrAh0GfS
YWigB00UrKT6yOJ8Dkhvx4oZzr17cXyT+yGBH6PS3CM57lzaoydKdJQyodwMI8lo
pgLkKC6wLtTDnp59ZFmhZExbarXrkT3PHUdmn+5qB4UnLXeGN1XHsFgfEjRcmgZ3
vYvOvaXTkKqZmRPLmNjFUPlmsPdAgnbQI7bKIDl/vz67WQnjUYA5lK8SQmFtYUoi
PX9cfTvTGr4h3kAuoW1luTXWDnu4vQRxB8f0MlN+T27tlJ1aHnquoUq+A7MXJu6R
8pBv++Qi7JQmnoyTzezyLRMg6SSKr2MZ6H+87J3yFcKWMQVXGPHvjFNu5A24omxP
GQcEM4uc/7x75YWBtC5hK1vLQ5XGEKxqrGH1CA0B70XDAwoWM3/WzxOS207rESZO
7z5adXRgAfR8Nf9NqewDCszGzLNV+Md92jsJQXA8EDodWkmbS5Io0eiSDqlCpa3u
bRLFqY7gYF7I/JJVaPj4AoShGi1Xo+1hJOoMEuB3DXGR9tEro7NRVq2s0tMOwsIW
fYsv1Gc7xUdAVX7zvXDBg+8xpKZsNw0Ku6RIvG5SMSZs9AWp3AfazVHZxLnjDFqU
igHxIxxU0oHyTGpgekWlLKMhx++Cq8+L1AANHauFCBzNgWEKUkbB5bhO8LyM8geW
WCntMs18BFKXz61YZ8IwTTN/NaWtR7fFpYRynhCD7hG8/U+Oa8MD/qfB2YijLZ2v
Z4q6qhtzOAvGM/HbVwwjqXREH01ZWMUVYIvjH5nm8FsCwZu20wYC4204aZx5Jl5V
bV4TrPkGhcBMMlKVR22EgnG3x4MABhe+H7Lpdvw6gfeeLwJwCLMfkvN2+TeQxhvd
W86W5LHuC4WSteSIYRpqz0LkBq+MkM1CYIjDNmBpmQpce8kl1ZuhmT8s5coOwOKt
SuZRHfvtUkbV/xAsI/VVJPPsNrTCm51qi7GWdfkZvaYDPVWlXnwPzvzOLregs5Wv
+3RHl4PNk0mv1VfsyDTYr4I3DNftnrJmuBWtykuwneXS1vCyvZjoOipUsGphXonk
0RZ5RY/cYHcDop6C9sjE8/joaizp+e+WPStNkKHF2fQDb8+r6g8UuLixWvko3u2s
wwlT8m+V0xbaTC8tqrNAUJMBgzFdFGNynUd6MUzamqPtHRsjLBPEzvgPCuJOcfHT
JDo3QKgqBllGkzSFSO9giw1vunwwq/XGf2lRga2Pcy7aecs/VbfICaJXW/qgD9iv
+xUntgftvOucjB/Yc/4MYRYuQg+oYQzwxyDV8ZcrhqmXNR88FVNzJA6seZmdZBpD
PZjEjMgc6TWKh7ZDexsGYNcNuowdZzIoUSPaA00aRd5bDzKF11rAjxa52qml+vBf
0p9hyZotpBmZuP5PX2e+LrU6hCtp9OiucryViJIg2uaSebqs4gCiL+QtAZy1nClT
7c/H7Cdem9ELEfM/sUwW2A0B+d1q/SEKrgR/IjcLPpRZfCt+zmTrve6jMfrpvTeX
/od16g+jDRF5I84616wQZrd0FcteWcvlLZDfz3DzuMqQOh2DmMEok9rk7gAfr5We
EoqOvKAhr7ahzKmBNIhNvpqdEVrKtY0Lbdm+XGGzNhBpg2NQFtdlT84nA3C3z5xq
o8rtBGPSqgDgyUA6t7agUQndHcNW1oTy9mbAmaFFgD4aKsdSYO1nOsGIqIVQ+ljd
+nCYXoXTErbccNCaIxHc6s2AcoJFw5R8618KezYh2Ezz+onrfV8rsx3vLXkfjcjN
nKwAGxgUND5jXTwSO9RKA9Av4J2DDD4q0wVM08QfRpaf0RmsmDHAyv6R+U54rq66
jFAU9iLm3wbECRi8rqzpzwsJUzAweIDiSNOdqAERJGISO87CogZeNJVvPHritn6s
YZxpn5PNDdM5/M+aQSIpFZYFdeYr56RwfXsP+qPqhu4xPTtv4FQF2MZ5hSovuxid
Rorv1cSc6C9vr01LKsT/Ggwt8YYCsKJ6ELtA4xvgTDfnoo8uZ41V5jmsjp2Zw8YO
4y7YwVziLOvl3floPHHqxlO5ywJn1OpO6fiVtHHeNpieQfAD3Z/KMIN8h3/h5ulT
aBNCLZTNb08oGPuki1dqwVpbUkm6sVQcFnYI0sBZuWqyR2fLlC9Yj/J7OFQLI+Rh
nNRr28VWaFoVtv6OuuOxG0cDUAdlMCStNOeL6tuHzSPNDtzXyCz49/8RnL/SeN6s
QdJJx2MCNbmk18BNCc5Gv65/bsADefwiQwbSrgoEEAEAp/EbMmhr7vQb1McwR4ic
bEyK/ys+7ddd+jux794sPBp9y8Q7edJXGAkiG1KOwBIEAiowur1wXFfz3U23p6Tw
50kBeJ00KM7oGXh/0m9EBX5joivOt9EU0+wS/UCUUXVgzEC0DAMawWlfzGEKEG4Z
Df8fiPyA91qMjsi+hKE8xX6VBC/3lSuYdCQLEtrWInOVPBeueg1CU+5qwrBTCnga
pa7kir89KrGrPrtzbvd/7It+G3l7luwFv4Yyp6h87GPYoS+1ncjUN8FJCFXd/sLM
GGZb8PFQ5UVFXGc6hlZb8foTOs3IzrCNt+evzaYo5VCysJLVeo4g81VWHxsYdRqf
lP3WYqBdsVyAiQyfGA17QAciO+L3wjAhN7lcwFv0Oj3SJKz+5a0cacCOKUOnfiHE
BvdLv0ENU2/NGNZSdlnRqMB2hdRsPKUQCuAGDQBegF4HwM7bbOjOChA7aRbDQ6Cw
EpYseuS36VpdfwUtFKV33K/X7tKa4ppMB7/mvSYI2Juz00IKQkeLbwvIOkBInM3E
RFmH7C/ouiTpcZW9gmBxY/kSClIKgG/GUCqhGG6QxUQa8ujx9zOyvywnKYydxXba
ObOVuxTItFaRqYK7CBaPjkyuBiX7LjMSjVgXLLnZgHe3uegTbXxu8Xf9AYUbpowj
dFZfDslz4631yLMjLAyo9rqJ0R0C2JupEb64x3kAXxyPNcxOJ8MicMscWbLZdMTQ
atXuqC42W4z1RED/3gMlAYwKgBDgMZNFM94SoWAEm9rIqNIImeBNXJuzUjbQ5VQS
FXTKlh4XiDCcgQ0Z27k1wDkdO69gEpPY3LKM/h2H4DEtb4yl0UJMvDYbb31a3Ttx
q3Dg4btr/iNl/ufDyb+76gYjpR5fOrFg+SZh5BTGE+fGmGdBTHiMieCur/RgSTR1
TqvczuG0isEVTcR1M/8c8S2bFLwemWuRM61PjXGQmYMoVR+3ruC7iNeJs/AgIjdC
ddhGvS/yLfGjK3YV9Sqo1ZnhTflmns23KlKSEkaZcdHQPfDXj8Fj2Pp19Pr31MIo
+huD1gO9W2su6FFpx6V/7fCwyomLiv3jdg/CnbyNiaT8CMcCb99IOLClBRV4yM/6
aZXQmZJlL3nWLLdxRuZny23wF40T+f98FyxiinzRt6EEiZZiMoFuz/rQ8+RRmLiL
gVZufScDA13NBl4LwmxqRAWlTj4w9Q2zWi4KQA4H7wmUKAEOm1FQr9O7ISmGxjI2
b4z84xPPOsRUTnmYk9gcWI9FOfvB2i9TIDEsZqAz+HosOysLvUl0vYsyZpdxjjJ2
DlVWdW4/MO/HxWoCM8B8NWpiOtBheh1r4MbZpgv03AU2MPAx/pVKGHxUn1i9rHNM
MXCZcYCCgfWSfmGjfSk7e5/OWaoCwhEbyS9jULNa024xcHhYmgx9bj28OnsAG7ob
+EJvBoEgR/ILPdNRW3Y6da+o9uTP16zmHaacaVACugnIiIYhfpdfKmJuEkvoxvTA
khVus8Hlj7QoYgjO71KSTDrdU4tT5v/akjv2iQTDg7XoZRsTJ5ovOxba1PAPfvfa
R+kR2o4aBoXOOaD5U1Tzz7WO3oRsltB2VphaNojxZoGCmere3bU2LHMmygLiirIU
HqYSBByqK7wdrQFSy4QBmhc68uUaxsJdXlfnfuquumpGbI5fHNik5AOSwKyv4LbU
uE0Qm7Ah7rh7kzn3OLEkRiQXtNw8An564bizM34ChEUDKJ5rnEan2NhhNV/Is5BH
Haf5Vp5IgMZL2x8bGSltzQkUJrDutKt+xq8sLUzQ6Fp0f7pGL7OX8tiEbinRLF9F
p5uCBXdlwR1gO59+IzXNmEWpoCGW27ye5stn7sjpoDLQOA5c5/JdMveQg95luBWr
NBOjZfFcTjnc1shwZik1kmj0fi5IgFmB2g9URW0Clf0eyZwGqL96iHzwCR5UWTmR
ZONjHqYPZ0j81vq0E73XCAPnmzaP35pmZPNc3e10Mz8vDLB1Uy7uwFssUQAg+dKO
3zdP1busmCm01tdpBU2z6DSXFId+B6hEN6idA3AHMb+p23CoQY45raJP8lkAh9bq
4qZnVrfVCA3SblaG55lDAYHwQ4SoBIR0PAD37IVOStzxiqcVr+ifSO4oGDJGGU66
vSIGHHGcRp3AdRrwv+JvDmOWgox4PGOlHIPRNHxI3F4zq2mESz5qfEQk2N+4z3Ws
8QXfh2jkDkcso/21HtHFz8ipxGxIUP/3tA1DiSVgUMyz3TmaHo5gKvsQFiqzIrv5
eo5nKPIc5BR4hvUl56fN5YjUqVA1VQ08HDURtThs9w2wG5TeVrHBAwyHeip7JiI2
sId+cN28M+Tb6Achgu5cucfwmZ+dWcN0sYYY3sa56v/KN/ZHhCPzQLgqQjdK1qPa
ftRhweeA1WSvP0suQJBd3AFQ5HMHrK/94p9nUJ9GKgynYYmzQ4ATNV8caI0rfcyG
/YJ9tCtBDhKBeupnjkNFVfDaKjunABcFSMXSTy1BE98+YIuBjcw5ekbOZwD86GyM
oaBJuza18SxfRNE3oyXqjhPtmR1JPAnNqDTle/QmIQXKaWQJuR/yM/yiJmL1NDaV
0zEQ5iJsYOgVErOVBJTJv7jjLNV2X1wG2GEXeuivwirytiV9VI08qpiMwVCedGdN
1p9zGt1bRzEPfZGmnzIniCtFhWvkiCq4hFGvUa+ZLkrWCp2CiRVJPqnQQavwZ67A
uJen/6wy6Wtt3/L1PSwP4FJNiK9AC98TPgWnVDB0cFFDL/rmIQIRUm/6f0UGHMpH
0x5+VLbQW7O1dYxIo881S1D/PtAc7KhSkR1cFYs/E4n+Gz+KZfky2RKBDdTsIqmA
OubZcpy+Ri5uqQg0dmhNtu6fMhYfG//WpOmgGc76IbFh1Rs+HXdHF1SzMArieQIY
5Qg7zfo1X2cWw6CZ/GGHgxNTpBpGtLfoU38S6u9G01VCuFzyEjkcYDq4BdrZ5vAY
/y5zGuB7EphOfLQ7HH/PTZACCqtalODI4sralUItLpN6onTN/EsYQ0OY6AVdkl0s
dZW9+rykJFJcYtmy8xMhmSsuAnemi9WDnY84xmFFArkUpMYwsZLhWHLUesPP3kVw
nQlMqlOGehZHR9MVId3JoYlu4b9IXD9cY4fjq87y8SeeXpw8KqTzHl0ArZdoGG36
NL1CoHCIjumA4jV8t0vkaMsZhJ/cenqMj61hyAhXabOw97GR9GYJVpJsCBxZvTzC
DtQtIEGEkiFO0KIeRp0zSv/ohbTNmFPWc+ekGijOcmy03Jlwjx7lR4rkmK1Hwfhp
zlkWivbmCpKDEETiFv1iRIkTaPXhLGCR9+tCXzSbNI5RaFRwu+lojzZ9h9D3QFIN
UG6EZryhPqXCiE/ckWRDm3j2uwX01Uw7nxMmsnwIHkNMLo7AoeevGakOqWcaNAV1
zqq3TIHsvAiDK4b4J4iVIQrtyMr3CJqRKiDu2ThodSmBRbztFRQunBZNYbwAbdhc
VXjbaLIyKpyq3ySFpFpHO6kJonWTmUXGaeF4pw4xC1DzinW2MoiJtUkHrQuatcAF
NWfFHXre77gGGlSiuslC9C1kKjfD21jztCONL0LFPjWTvo1FMCUVNd9HlzOsPfTo
UuycVRgyibneaxG3MNJdzB8qSZL3UjB6Qkup7JwkUNueMqimnli5W1lrDAc/WB9F
SFWcJI+p23csLVKyFCv/3cRLPPlKJ0TJkLOyYACjZoL8U886+1UAXT6NMyj4FvbX
zln6uhlsmsmPC2Aw4TlWNKA5KI4x/IaIw7TzbErSfXPOuw6JF8hWRKtOa9lGulXo
rJwYjECVFho+ggUSP0+9XMDNhzoOfBviCxz7XvyDM6ZE3K4o0uNy7BFEssoFPrWd
QwQNcL0mDjcoKupkr0n9a+bIzKw2ePVQ8e7sobbxJbAQ+AfQfywtoR2oFHw4ujOK
NMw4WNRUVQZVRKMPIlnciWUhRXxM3qLcAGbGtxJY0fB58rl5VzeVyHzupBPR8X9B
W/hp1qeus4oOrwCzHV93fCoQPgmOMzHTdNEHe04nVBIVdyQEkpjTrVe7I5TLhgv/
yKAMsg5zr80KclgN8MZNo5zOONE/+wTao+ZjxQitJjMS7EArdcnamgHJ5HhpMrCj
LbfXIvbml+uOb2QSl0kJ0D6oSLuFbbTW9m3pGL+Gp2kGrHCe89wJc8E+dTEtaIin
pWnm9gpPSr7VRnJ37wxBW+sZ49WvRSrNcnbeMZ0gFlh+Fv4r9+1M2DY6ov5aQFe0
s5XF7G6sYz34qzMuEAGQl3lbZcrUvhAoz8uI/dx3YD8nhD3nrVwH10nw6ykwn8ON
juPPezSydfjPKbRl5RMgRUypOnP+gdqPD9I4OT060h/aAZ41Jf3aYS8xy6KaCU+D
JWh4zJhciwY5Tf4XpqudRbOT15I9ONivD4aqG94hxW1oBEG5IVlC1Nyk2ze8qcHG
9KmEeWVK0W1M777W/bQJVDJG0am5bLCIQlfjGhZMiSP7Z4msc3OA9ywLcX4fTDkT
TW3C5YWOGi2pno6l2AUWu+hpco75/C+Ut2WMV2O2xaHdCVk3/NGwI8q7LRc3mSHw
GDEsZ54hHWfxjfDW8/6i8WD6mU3xoHanBmSyo0CksnBCYCT8ondUVY326XKSv3nK
x3DdHshRqsyaiDn2+agVqHCQL4PuKzpm1C7A05NxWZJWtcnElPpLpi9fqhcDdUq8
mtwoIw+kvQKaKJrvGVPilZZCji7a3qiRro7YZyCSpo/KEPc7TZ6md+KbACFwbIKp
4p2xQjZpU4Boe4+XEpEYdxCDlWdCCOQKT0EPtLTRXZllqCo6FW87Z6GjQ7//p17q
gvSjp1B3iNmg4shJ3C9crYwPM8QcPOXPTFjeeD3v588MhfeUuP50PPAhyZ9S7n0U
fYRBbpwDQMJWFHZv8CaFKg4MZ+ag4L3Y16HBpJs3ZsIMA4zfQ22vBjTA3YuOzKdt
GUX4w0WV9TrpkAX01fcw5tO78ApM+Uoapm5/mgTaFmWrRfPpgS74/i1scFdgUBzL
9+TzYp7iPEZFgdex6sbMnbnom6BLvaF9hHHXbNdKG4SV9k3gTW9jMTUPWdqTgUqr
M99LflJZ0beFoiG5HpBFz0l0bBo8V33vGKPl9JP3ia1/pTQ+LbxcMblwSo3Dv+/7
trVSQ4iumdQcoC1FRhWWj65ZNycL6Ibdn41wxO9oIcZ6VtJUjZxioPfeu81uK4wm
b2lyalaI2WmkcPZPmxGAGNG4AgmrWc+ZiPrZKdTYyRfGZ1SOX4waVIVdqE43Y7gc
BSQhsKxjwqyvRLhsIJ663gAb1UUuQSwzILM3+BVpLLzJuBks2hKuP8z7F/BKdOfD
Qo5NyVAYiD77+LtesU4gYR4XCC66eWggGs5hOO6f9BVyrrgv5dneIzMxNV+IX8KT
catCLXu/P6zPqdEFl7kv7abQzOQe9Oa+YkXBFMUnk+MyvZvgQwo151knj2ZmI+lr
eP+q3GfA9rGDJi17r9EUmnkRNNY4Ab3B6wT/kSW9Jk1JOGTEghjJWro96Fg6I/aY
o6SC/yc3KxGOKmCBPE/ywO94qJLRMbrfh1bnmH35K+3hdTn33rDxzUQ+CxKkERcL
rq3wo1PimtFZG/+/fxqy8XK85i7lHtNIMJVJlm9mPBLQXJDAt6JbjsJIrgLpAmhe
x/f/XEpkDX72FoZsLt8vz48ad6H6wlbglKvPuvr1UskYj9i+4a4BE9B0Rt8L1xYu
MBuPZGy5Pa2UN3tjd9giBAoGjM54jkKbtENWTjAZNtxV33Lzp10e6VB22O7wmPFg
eZ9woIaplJtjNH2nymKJbDiwFtDrBdbEwH0H/BeafoAocQvbFA6Hobarme4lV2P+
rSnwNPvpFoKCwCb69YGeJdHuTGfiNbq+yBwtHEnmlv2VAHmzipbJrSRkQvHvD8Ol
pzTtNh+/flg7101LE0mk7wRl6KW7iYCwWKRt5851QcLgnko6QUGXj4UKhpHwF1en
CuugwwGR7p1bogOQL8ADbSCL84Gog1QrMYPf7xknRUPITv1WLM/+SQrvMbTWFzqt
wG7zxQL6jl3DHPAhejiljYeSrZvMs4Iy+qOdxOV7iLdskIsmDSiAW5F6VulDZl4B
1MbfgzR8fPVko5TJ6+blP9cDDdMvGz5qWdUWCqJ+TRw2UCqI0ODNpabr/tr0uUJd
m/5aFm+SjXUmt+cKYRv/TuSrosZ/PVi1Gp9iAFUDSytai0hsR3FyAQQrcaim5SlT
GHdDw1lzAXZRli6YxW5U6/Y2Hzh3I2SncMnp71HMSs6itPFOFyPJ97YBCzsYmzcU
9ipByn2mBpc5zbCmTU9rPWI1dc3VVqjRU/zrxOWJU2pN+bxX2T1qYrpTlH3UxT6S
9hYJMn/TXC6UrXuDIgaVN4bjcr31+VgwOhm06mrOpgAz84E7AYK/iKp86t28LbnI
UIWN8lOw2ZF8fvoA8Yu+LI2St2WnlUC4pSA4iqC1bEqmzgWARgs6X8a221IhtvFo
icVug8X9wu+gOM0AM5Cx3vXRz0BHIvPHjQLNxcMOWRKGxQOJalEAXuGCEA3osF9S
nsAxYiQxSWYPXdZSNkGOhC4FjImLrCEdCeJ7ofU1zeUvNH4N6CQZy7oJBHMdnDiX
EYXLcCvfBbQqqVn31+jiDUFSeKWZez5peizSIwPgAN1XdiMrdZwdR6mkbj90F1su
YJnEYO+KCmCi3uNNAddYjyEidB+4pW+G+UGhOCRJ34BYrHg/J5qAKun1JwGUde4/
MzHyqX8cL4rpS2XGvkeOjcP+SLNelIPNB0FBpI3c12MLFredrbvbNEIsjdUn66a6
ydrx0XP784HSlTIWu0peHnSX2SRKxP1tD/pulJzzcIz73oMuTkA08dO4pKcWv/HZ
5OxbEv0E3mboJaMGS09r1Buh2/osx89UxNb01TycYUElMlKfNkeB/0UD5FH9VKiX
boEgXbaF5C4s10KfxWDB2aNz+KHnB3+xHuhf4Tqfr93QTxMr5YzBVrQnsT9Tk/IH
WSXiYxpbS/A7tTrSopprpJbOf6dni+dA8BV6sOYA0GX0yGPyr2QzxRE5cDmXFiMk
MBm1AsBP8MnYbSsRGxC46rSl7aQUnZLpA7EwB0ICrM+qumBK3qQoARy50Hqon+aQ
uMMWawxFBM7aDDhQrg7hEILURKXAIpUfJknLgdyUwB2fW+MOK6nBrJt/9llMA/Cz
U977JL75Hm/DmSdWCf7VxeiO992jtQOYTnqiphW2fXM7DZt2w9j3h//d2nXIBsFP
MNpT+mK0XHdnxokhPJfosjEWacPF6+PSw0y9EqqMVMzIHRFjsHMFPLxrkHYyGODA
r2v1Tkwi6VcntOOHok2s74dl1QJxiHwHVA7CPBkdu5AH6scbXWA1yeEI4HCBth/A
aPZT3oVZZrexuCtpXi1y4Mx9OW7bUx8lk3eovAkTPa5z7GHoFqQ0kotbWePlAF37
OYj8pJt6hlxCC1+0NScibc5oFqSiKtC5YCkd8VBCpsQcwOYTuGE/N3HKHmEcNwYd
MnNFmtNM7ZW/69JM7PDeGAo+D5T3K3bepR23Db4pvuaMGc697XXRKpJquAtbNFtn
OmG0Pdj2kBLjXmt11hEdn9PBH5mrzh3POFJXC1IYgKyVn1ywWIedUmfTF+R5KOTi
Wn3/apmJ5TGQv0yREnoGitmYDQfWKSdHaZRfJDgQsrQbY04Z/gElgZrr46bXIYjh
FrbDyTxdWMIqzTasQGKRY8ZIubvTbga+Y5Uaa/UaC7FtxMbLgedpkYztIhKDZFiE
snTnfWTwZA7/gNzRbQ7QX8iILqRHxcOb778NnlYCO+IRNykIFaDZ1UUqDfU0zuQO
MgquE/HZdMe6hlps0HhAz/K8SQjhp7TFUiCItnW34A6cj2roGqhnRhTrVgV7fwO7
SK0lBYuTkDfXgB01EmvbLo9L02xlAlzmmGg2ZyIDOZpUh1muM4mWQ0RPHI7gBT/h
hNQrrXKtrlw2KtcwKfhdsMLgsSz3zCnsiSfV2Z6CPQWOfv06OIURPHQjoxafeJMB
8dq0IuyDyscGrJeLTeNtQ+fKhGt1U8SExz6gTxczZv80hUWf+ft9emoLdpx3cq0z
ONqnaTsrByo3XB+/i8/78kPwx6bP7ymCjDUIyB3ZCnZQeUnFSQDZsBg9CFG3HiBc
fDJLunIOPGw++7XxLHRQ2aCGzB6xKJPFMhwMNqYqCrqb7JCmxrf9/k+nmrLP8vWe
U1BL5MdDzRRbHCIBxPr3WawRnBL4m/ALW7a/UYk07izfYIWQCncs0boQH6nwv1Hh
HGg84JCrFgDoq6Pei60NehtbkFDztej/VNaYYNWN941dCMyYgXDpZm5h6/U9Y9Pv
r+bDsCa7j2E3+v/6+x3d/pzqBXMEKpbwl+NIlB0QIKpN+TscpmcMx3MztK7eg0st
fZ4NbmOZtUMDKLCnASeaqqPg6v3aw9amWCUHYjtDt59TKnutv1mttwsG6wszcs1d
awqPB1TvluXlfsNJWczDH8WHC96Z9w9ZAUdZqAvf9YCbS4lP+Q0xf55tvAZBg0EQ
QNpuzLuJfK3HA1yJ96bn6enxBgjUj5o7+9sPNqZyiNdqY0+Jq+2sUfoJfuHZgq1E
RpP30QWm+h00KYdIRDj/gdbkdQCo5vJgU2uFZWA6/iugTpxKexh/k1W4OgKWAzOs
noEewn3CrgfhqVygmArZZT27HbPLN/9NPJJsrkjegjxJK2mo8+THC2J6HZgQgn4k
ONRD4rmrlgYqj3W3Q7jEhh3jBLJetQCOUYfA0x8K5Wx8o3EatXtko6BbwDfJpKJb
jdtoVDaYTxfc4/t4SqERTdkZHaSqd+ac3aMWLoE0gSZuavfO3bA3Ilh24GbKQh63
JC45D1JvWxe2ct/TZ1W4+Z8BDYx7Sa567SCFH+zMfLfw7zsYU2Gdsd9IRIvPd0aa
TT1fS9RzIFDGMQ0HpigYST8gA8LYKCAxjspE9IANu/mBavBJ65DPvBlUUizvaLpb
mDuadiU38lsWsvbokKeUhpNbmDCL1tmr2eMcxVEEFoOjcPfsiKmzKbQlMEyTXJE1
tYPCL7BhAoPzAAiUGz6Yx+7ED1nqFUs/S4H3JmmKubpjfrPOnL+GrcF6nlaN1q7p
WPWk1KNQ8drYLQI6J/Q1/g+2+TsrDMpxLOviuCSXQC3LPm2R/UClYZhLH49CrsDl
6t3IUyo1Bho3XijR6t30JAQupwdPF3WW3tQz9xHZJ5BznlSzX7xQFpgD63ZTIwOJ
1UOJbNY7X2V+j2AgzB6Ure4yFz2V4VrRzZwv+br7+Uiu93yIiuSMVEcuV14WLqk5
MWsH2oNEpaP9OCr9tl2bYQSwoqnWytszsNH8SXt89dDaW2hQujyLoFJSzafDEl92
GtOluww+/gqqiZNWYBxCZTAlEDTiv00yTRufxng0ZgEAhU1mmJZd3IChV9DlCW7G
TEon3neTigmbb0X45aZ94bog70bWf4eGjKg2lOR2o5/XVGvmK02isyHouW920C/z
oqBCc6Nto4hFR07Kt57d3lngvJi58CidziVHs3YYyScgMO/HkNuTD2thrl0aXiba
Yuh79XKeG0XuSwL22RIJZ7cDHs5c3qBcrXCnbRFEW4qll+uHgq48yNSCKpwmuFL/
dwl0GQRI+qvc6YBixGf8VA0ho7oze9xyOX99IvZx6M3wboOKKhCrYA8QxvgFvO3h
o9q7GFyUJ3JT1xTpuYfwxiRTXXAhlUAF9ad+fuaYi5N5bmfKtpgYKVgX9E8zPwbb
QKKOZKIVqkzPY2Esa2f09DuzOPpSHvojibmxD2l6B81v619kL5Z4JvN14ekKLeLB
oxRhXaPmXP8r01lXzPHYmuBJzFL70ocJmmLxB8kOmlULiGzI1vCemNVgiBj8HivE
iJgNs1CT2oclycF13sJtWS7htBqRZVUfybeJ9n35jEQTlYICUREWKP3GZfKI9hSN
wZgbDp7CqDMU4bnfYkYdccsWTUYH3kKnMZqfZeMMoUWPIl0TWlVOo7LFHA5S4DDt
x2moSO0qrL4Fil4GB1V8JkMIH4VQ1pMU88A3lfzFDZy1ctLMPNxI3tygYpL68rdE
Gwm82Fw5lNzJ26E7l66hqM7bfdv/SJdBJZ05X0z9AKcCCawG1IamTiciyMkNbqpd
CHhHK8k3Xh1tktFZc1+E0v46s4theJCI31oOLZRJ0GdYz+LjAp2Y6d3ktTv7Jd4E
THjhKONemfVGzNy6PnmmcRlGm1lzMD2rPCCLaVDNAyozC7CUsKXDR2ICJGrBsd2A
/DT0IaUh2i6hvEVIK6qg6Dc7sNucj/CCacRdIzHe4ODSy04DHgTu/0GVdvF7Oj7A
mlhF3+W3h9lmm+MB+ckPHqXauvTzZRuwuuyYZWlPwDmgjWj2hA7+bN3htAYiAxHB
51ETeFlTp/JMrS6FSA1I4SJR0bjL6ChVGVh9Xkw6MqIyBEg5RcKEP7AC+C0Bn1o6
+WZqQabtlijZd+hf83YUeGDgSwc5MswVyc271sMPS+t9FqVISymOU/e7PnzezGE5
4k0vby0Z4fXHBmNiF0LZGGIPudnWVcAE9REwo6EgaZkmmfE1fgo4R9qcs3r2dWsp
jAdlE95P6qvht10dRy5QOrEg8oBqNUN6kr02lOK647xLnpoIUoyIeKN2XAvWf/VQ
xRE4QEGZwngzALu+z7gFt1l7PDNR89XljuRylh3PqqO5hha+eWClW39VQxNxPaN7
FyRJo1ZK/YptGhGhfxZGKgWZAZt08ER2/l+BUfZftqnZiXf05WdEY7qut1D8O+0A
MkbCoA89clkIp2wJfgUT0wWd0OL1kqtZRqQXmzRQfOjj805WNak4zBwoVErz8MbB
RCI5Q+78YglwFfmUuKiu4gtkXvFIL274d23nwN7XbNuBWgeSPY1s/C2Bza2RDHUh
+UYTGOCTVqOYBsNfE0Hu8nAo9b0ZppuTjIENdv1GIqPPDfass2JvY5GotXn79Gn2
rQ0JT7UspTI1mHRZ1eC7iJSLJgsq6uj5IXd9UPSTR7xXZKQUMxwaTmLtNLDUb8Lq
LG6W3LMaw6XZDf7qPntl/aIf1n5ytYE/Dmy0BB/XHbuSEo0fx+Srg9jx4Mrv19Ve
OsRgrkvtZdzKNOvPnaS6x6LBt8nEmEDPDEagFvqKGuGfAPWoYJZgOA2/LXgC5MUd
PZCZSg1AG1oA+iYCTT7ttWR9YBInPqmpS7nQ6I5Z+KEYub0/ROP4uTaAEPxBXm/h
zyGhDR8Ozpr4TIR99EqNxNhYmRsuSgVy1/zi7dLHCLZo9xae3U/DdcmRqVK6s2Nj
t8/GYwtfr82YC6ZCAAzKBhkssMKFYC7Sq8pSocClqrOTXt7T3XITvYfxCZCf/Lax
0iQhjnWC7kyqF13s89vCgbYck7vD/obQ4xfIrAfFcwGAv7yTxNDqbKAn4sC40uA8
hauuMNYtBKV5JM9aVwro31vKawj3cWGXCpO9kRifSxUbiVpLwmPJehce3PGY91vy
fGYt1ejcshjxZX2mlJqZCEsoeoGG4/0tb7Ls3bvYTCxZf251KYmRWIeG5IyD22JE
qOGMvDesqb474x/WhzbSRoMBwic9wI1xyH+HYj07xQeSDMZcopCEDzLbouO3XOO2
EV7+tvhhM2wIx3UsoTTnS4N+e7U3TA3i98QJnBerCGyk+8adqqeSuVvCd+4wz/rF
oksDwi5hLiA6Nku2CAPvvMCA/G/76iUIjOOmBUolv9iakqo5EXOkilouIqY9B5nv
qPGgx+OhkvGdfCfCU+w/AEu/XC069rC0LRcS7gFWztDZQL8nEnQ0PQoJeEkflR0+
gSV0Qi/+MbbNmnMeB1PmSuK4YkKaCy8WDQBScTkeJGZUB3pbG7GnoXZVqXnDfScd
/6eZDy2qq9PGdG4EnSyTuGqsqHRcJlsFJG7SSXhTi26ILHUbEwDw2Qcc9Di+nmv5
1up7WEQpmYFshsK3Ky0fGUEgbInmKxrgmgDqdsUlzwNcklQy73S4loenyO3pypvT
scIL4FLUUm2o4pTqBZrI8E/734uZAGO8svKos0VzWrXLM4aknJajl50vdxHtDAPo
/cPwUhSVTXCT/23AMq8VCT4wdS+j/i6dNXCdg5a/NvkrD74CyBUfIEUs5cF+U0XH
Efi3ix1eQLkiRYrNVLnFPHVR3qcONO2aJFIF41kephbbi6AyH6VVnxJoXkeHR+YX
7Nki3pygozm8nldBrj8/5youz7izi/1BuR5QgkmnSsPXYUxYSV6mBkGGHCveyOHN
bzDiu+F89B2dN02sVsvGD+IQ8LccJTd7xMQt/q8ro/vZyopMHiDOAzdRI98nokFt
2w3eN2AegBN6lfw7ZjrnYwaMm4JI2w3j2gcE1/RVAamPIhNpvlCSj+grtot/hfN2
AITaIH+bIWasv3khJ592SpWULecaxck9gsTQsuvCkny8HRqzPByC/59/ojk2R+cI
I80EkV1baAAwYRBzsXDfxMGRnva/mEoIVlRPcH1bux1IyOZP+KqgRU/rkPZh1ei9
xklOUJ/9qShHJLFJ8Hy9pDhTlqKziqxGctvaFweXZco6prz5Rchvt8uSLVpR7tPM
Q0VRL8HkvLCIiBtkMleNO3/OHMCKFElGv6LDR+SYlaQIEmCej6nOq6ko31PK10qH
xeJKiCelyIecgsYGYbVnvGLx1S7o/JTPfe8gFX06xMCYs7np2EoBT4EEGf79/TCd
cOCWyCS5kGm3mpRd6708pRVQFLlRa7Le20vTKLUx1qkt5hQoUvUARjtpDGaF8hXT
s8ImGO3KUVkywWnfZJOGpTUITcJ91NKi9neICaWR1ErDEvRkZcU2Nrmg0ywWhJBd
9+1TfbgRyD3N+q0kc2a6TdTueY5xQEpbkC8efEmB/YfPiYQVx1nNqunyxUY0ANJp
9GbTwI0rYmvrN2rUwBqZrPiLfWrZ4pawKX4ayrsbs0J8PWYlntxxCrBCBOgeD0dj
hJPRyeGh0noBPAIe/Ra9tcqz016WTJ5WUwLZ7bTr+ACqQ5X1Sp123PKHvAZl82jt
llQfhi5iT3jugX7tPfL6rYB5doHEAMmVTdyQSzbpPpRatBgVg/SjBq/EHRj1xPkm
Gv4a1V8O9dhyjy5fmCn2DGcg9RiXv0ZOeNAxH3T3f+NuvT8KTy4j4ywFzKHIbMgH
BDvfqmTBoZ6IS/igQHHKBS5/Ofny6fTFP+675+3X4ogU/5Ygkh6HqZ2cWeNr7fGu
rPl4TxmKF5g2+SqvzTgOl5yEzRzxvGvxBn+B5zLq8jcZlcGhsQHqN7KylPQ+24Z6
G296tTjKpiG5gieUykA6ZNZzUbDHjD+bZcNfoplQeYMeXjmByE7ATDtQfAGlh3L0
ScRwNkqeUjSLb866sOkLsKQ1Gp7I9bibhtm5myIGCNp8y8eo5gpyJRe73GouNCEd
5IJKSTv48CDP9fGZd5LaENhnKBQdgCDMFzeGlvLJYPKaDe+r1seRrGeVn9ylhNxP
heJi6e/vwvFWcfFoUuN7cWYkRq21BvgfeXBZQfbZ70Dc9Pbrv0iRiR0j+9Yufxds
5OG9WejeONHJIm9dC7R6aRlyAC04fmL+GcNhoOn3QbPp5ggQBdHmbM7hwmxfyOs1
lEGXxpmPiIYvQJB3kn8yjZ6FW/iQK9oFEODLb0H6Y26vOOOaah1sa8tUZtDSiNoL
mEh++uBOwYhx/PRrUlSS2Xa8RP+QKN7b8OeFySz7SwkSqW4LEpPmPDaFaPESMl/B
6Pq+/TCa94T6A4GyIlr2EpW9svw/Xa6FlVxIEZ+yjQrGMp+B6RKLJn27V7AALBm8
4gKllmIRBMa+qQm2gPzBO/vYnfj7hKxQFTptR4zz7hTYUMuIx18MfNCBdXHOr2dW
XSYOrjzvWj4tdYaGFXr5mzQkCLaW5AsMFYtE/p/yyJuauRaqQWEqhkuvfxX9ptEC
nOb0O+oLavqA0wYbVz3UGvmwLxHo3lmdrmsnzBswMbsXi1QZeybJT3v9Vgvn72HQ
RMKp4jF9Kfh1xezNCFbSSL1xcEPKSzMKEyLjZQL84Omtjx1ahNaSe6+utJ1K28x3
HRMsMnMvbXeMHb3o1MPtwsv8uv5iuZeaWx4ZLtQctBEhQhIooH5Na6/qaDvz9lAn
qeoSSRqRnYCzUtFq23gIZBi+DmlVcfy4eSK3P6eJYF9MJfPy7XZYEBhaSrACVkcx
YTuE2K+AUVlT8T0x+63d/8RqdiPVrbSXQRwWGRN/dxMHXfzQU7MlYiwXhqYvH5MK
K6BlsaspMVpPF1sPUhd2wfAr9AHPER+/AJZzE/q4DJ9nqIeDj7OD7XOdRNdF87+u
18sMfl9/FO8l9TWiiKw+Kj/593D9lyheLJsA4wakNE+Iz4gGuHTjB0XzC4UsCnAn
gCbx2NFEJuYy5BzcjxFWFL6KzoPAtgGUZ3fCfMH1hMFUc+FrSm7AfinFfPe0UWOD
uwNxnf0SjBhUD7UQ148XSJzFd9+ba1ehylzhgbD+xEn+5KjRAqUNS/lP2Ygt/BwX
EIxj+WdpcAjN8qHRRrOVdOurfp2J57n85ysC2dkcUMWyXa9wU45a2Iiz9Hh+e30z
09Ut25ebHmK+WCLnBSipodoLCLObPagnkU9O8xtPn6GwAsSKCP3DOv4hAwLRcFH0
EBq2ycCiNa75Q7dxKWufCXXaoPVHXFq4RbdnLxqdUVdls9LYrOni2EYkM207qruQ
eCU+/gVQEPR3TfU/HlqocYMlInVwXV5kOhxgsTE+aYFr3ExhuSc1LPjhjJOWQ3x2
2xQYP4uWOpxDkL7wsQgHP5tiTOLgZ4WqOuHJV3yqIVX4ktBAdei4iCEz148oStGs
WasOMHhwTXqmPtECJpTgY93V0oHIOAomxBv4QLKyhzxzJczTe3mVo5MBN1Elg6I4
QNN8/cdFzsamRAl9iKDjQcDkubmLWXY/RHlgB1NWrZK/bY5pgZCZBhBuXJzpt9Ff
+peRNW0y6Q1PKMdlCe++qj+O1BEAEAdnEmWahYgJolY/uIiAozmUZ0e01bSJi2o3
Ta527xUgvBVqZo7T0qzNJxtg33DtJOCzn+UG6sKsoe5cQDuw1Qftqq4dz9sSSa98
bX2YwV1P1zzom7yXNXl2ji0u9VAhkkeyLlcCA1eC+7BZTZGUnaeaY14qozwf+voV
ymLU3SdjEHCb2W3oP7RR+vjX0p4bAQnTNGuxjHHdp7vdwMjSeHguJ3NgSPOqMqq0
BO/SBTGqMwFdJAPgD/dZF9jp+FxG4HKdVGMgtuiK6PFljlgyAE/uaE2ZGAVKFtc6
Wd0JKnIBxnSEgUhRXbQ/xzF6yJd+1LltyzzS9UhpP5tuJJoj22zzkDli67+OUN1+
Opwbysa91fx576cYcEujoVIx/4h0J2K2VyKgJmjG0xNqWBZ55DuP5UBAa2nsJLfn
oT3ZgGM17t6LGOrwA2l/RpnxNfOVVQLk9iVkd2TB+oymPEVRxodcf5XZB6Tnjswa
4ytUeR4jCRhTIJsy6cFDpoJIRBppYWL4RJESkj2w6cC29JUvbo3o+NqBRyA8d7q6
SizrYa76CJxLkHJshCFcJmQFsnNy4325LGvZXp0JjyvhT/6vjj+0lT/1uP8DQS7M
UqNP+BXR7YKetNBUk1BJiwFr/1C4YV8othn5unpBQ/JmTkqXcudwcxc+XeIC5owc
PVR3bgZcQ6PNrpMXkWx3IfsEHmEpYePoUk+mpVWLM8mRVvW920MLqdIbGsJMhjk9
69MSdKfeMTKMBU558Egs8nEoIYr4tX9Ogj5u7I5EDP4+AXfSfGQZmKW2mn9ZDYYQ
peMUAjSTMAqSg82ZnNQo7HYU7OUPk2O4qS5A6QgoXRuDp6XRchnm2jNaK9kKnKsM
`protect END_PROTECTED
