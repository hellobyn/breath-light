`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSqGxbr1ewmW/Y1kjGkXpTY/igMgnP3l3BZkBBfa5zM3+fhQqbDQZ4MYK/VcBI3t
Pjrd0JtHZi7TZQbKfZTjNCYXsf9F4Rf5rQE2a0YjwGNz9WgP+DIWHd5Mh9IiM5Av
9toi5r5uiT6m1pcXOk/kYFIBCedxbYlG6U1hPr4jZisyvdETetbiNMo++x9rdCqj
BjjU+z6bdHPJkkycBAX5lJCBSrC9wkFwvWJc4T1Q+WHAqtCG3n7UGJzL4UKDAitz
SIDHXemI5itiKmHKz4QZjW46Gp7eJMZd1hLH1TYAmugAhfiHWmC4rIvczNbMHwgC
OjjIibHcFlTrZyvKkrI2QwMJ3sAR2tBs0JWXn1bO2+xSq62WbnfZV5PiZHS1NIf9
irdnQ2ttrG6YM+ZoGUz0aew0uI2/9/AX1xzAUQKXWtubQgIAqF2XuDJEwxYlHk54
Yb9wKBQOIIfQmICikRKpMYmuk3snq5ED5l2CJsmOKWgougIKLBHQOWTGAbicP2Lz
Cv75W3wm9vMzBmWsvkdFVozgP8C3+rY0NQO/3pfVaQp8NHsauozt2Obb/eUlv69i
GI0TaDdoTbNr+vmojGkqtni2Ui3/ClsiSfn3P1QSt70fDBnmeV0+xQrvgGdZULgP
ItcbnebUwei72HLEjlP2tQXOM9gdou2jUXLElMad6VZsuSJHdMFLQBLqSxd5vANM
lJKSh8m/M0Ub991GqSKjvUdKUlEfwuH0/fiR5K8XPVE6gW352LUpczoqfnxk3cWL
L/9TrY2PXD+N7BU+E+Etkas2zu7l61qmka5N5TUTZxEEQjlUtqr2tNMmKg5GKU6o
Kjz10ULzj3KUlUc3sDVp8Ci3+U4BgiN7jFrc+J54f9A6ZZy+YqiNKXzpkKM+G1bQ
nSiWqexXu1OKpQ/TCZ0fEBhziW4nt7vV5rTdmzUbFf31tXCRQ1J5LjOI05QQ0g88
0q4Dr+DrPLgZbUhukAFUN3zOFrI/7yOWVAbEWkeTsPmPTgfkI2K7UqNicWW6EcOS
21pNznflpgHGK7y2UqGPXSFy0D8yu5jelzOwOejGnOyy2bEI3tcKTYYwkAQ4/xyi
I6WE/aBV7DC6ZylCoYI4QNXyCu8eWu/GIrYQ7YIEersltdAnK21S+Q6eyYeuOdRW
+WjGHwQIzoGbz/Ck4zh7Qgx4IFYTEgTWvThYTlecXi5kuJoV+ONz7/KeFoEqdKn1
r/dlt7Mds2VRIhwTEhGjG5K+iLOcYAJjkdvsw5dYm2zuzzAOc0s54ciJm+FzdAJF
5FYi8Fc5QOQPS4HIqf9iC/EpyO4XoUkD1n6ivaXjth7g/VJBNz1IA74mwtbAg/Jf
4TplPiqKUQzQtPX8elty5ye7GycyqmKwsAJ2dx9He7qZdC/iOB98+p883+7LjdBR
/T07VbJQVUxUe8YtJPUnOUI2tInZowDJYg9OKjE7hyIDQCv6bZKSQcDhqnwsi2KR
FM961SWcBCsjEt7BQbni8SSx7PNv4qi1h+ROsfnzeQdkLtoorlU7fJbdpwMz54q4
4NQkC8VX/oluF7L73+oKgE3tdIxJuc4fwIjv7ABsCNjQCoTaLb7TKyFlU/ZhLr56
FIm6Q/kPU9fIK1rtWzchC1RnDmhCYdpJ1fimVhnPeU6DEgkS63kB76qVNbGSKQld
mlhHBcnD7ZFzWUSyfZTnKcqqEuOkpbbGHaKJvTptEyT1TeCTxBUtubZojd64Z3WX
Qed1do03B5wfcab9Cq0y6aNLlRd4GBQILva1N4xGmPgBgx+dGsE1Jrdh3hDI+OZA
PnwYLTqYHKh59zzVE79XPE76B4aqgHtR8xMImtIOzKoGjmn2VkKEFks7pSNDTS8N
5iwUIIzlTQ/c82uP8iRwewhmfVbeyjtrZc/BazbV5630ec6xxNYquG9p8B0zKk4K
kCah772SV6aRylKW05buXr05cvf+quh8XVEgloLt8Tyb1bzXrViVgtdPgi6mBZlY
oDhdmI9gA1g80YF+qZF5rb85vLtyMrZtdvRzGdkacIJMSPb9ZBxvQ/Lq365HgX9o
ZjhSB/0giBGJppZcJY9QNPY8V6mfq2/DKZiVL/zDzr669jnUHB+tJ0QTCnomcwfB
AVcNQGgSo+x7rxmmVjgQQy7ss8EMSWl0/u6MQuAtJ41KOtgf14jx9TqanBlLYYmG
XoSSvRtqH87hK0wSaOtAaC0gaUQbEf1jYLeJ9nrP0VqMyE7BZzk8Asa+CPruDAVV
mDlAXacculOTpdes/VwUsbo94y1Y1LjDk+AQvmC7HJxdhHlSz1184P8usJLeJGvb
RL6tXiniinbcgFRIXA0xQ3z4qpdAYNldjpjdTdEkt5tNaa40WQQsHioDegdCTcGr
IAFL6X3LcbxAztJF1stK3uJw+B+QnCRhjW99pIbv6vcprgdWjpOOfAQGp3kHXV4V
wFgklU3rWku/smuMIbKKvsQEkTSZo5ZYsMSP0oZKDdQqa/HKPKFPPsBlw7Gke668
3HSN2FSj+y5ExlBpnIsT8M61vRy0Gu3n9/ru+t9R9JgnqWitcocx6Mjh5KVnZuss
OW9u9PdM26hYiTqxZzA9c8sblx3zJdIt8c7DbfbWZmN8i3U02uYXYnVt88mDz2Hp
UlT8Nk8eFinEVL1xUvQ+5QY1feu1gQlOw1Ur4HWupJNTe2r8qZFgKRzlztH3lRYD
TYFyUkUzK3M0S7Ppq5l0XNVjjQ8EuwdJgsGR4MUCE68dzzS4LMDwabTJjCfp0LgJ
A8E/JfWWJA0REFuAqRFDjZV8HY1T3sVy926MEJsf7d+ShEvK6uMwi2+qgFTdTHfD
Q7khS9c1wSWQxc5FEOr0eK35CHh57CXpk3vPV1tH7hMxXz7Gs3D3ty9wIK/q9IXb
Pve90Xa9STRBhwYthpo7YeDs0dgOs6aJRv74cjGWdUBcr+yQZvJsTW1tXKTN+1hy
mg0e/9Z/f3OW9LOVBsjAGKJhQTftIXYkJPMLqtaPKnV+rpZrXu63xNRUdNs6j3g3
F+FIqa6ywb3dxgeoPnMCGGDtv1Y5n1hVRSypEH4/ey4rfXte1o9GmPLoUXkdbao9
bSusmFZslY/IyPE+hSuGrz9JZVcqeo1EgHs+DfiBEDfqMTT+tH+3v9chOBLfno3w
bN+l3Ir9BRA95vG0YtCclgZAT6NNzuLovZtfBJ0ST8ZrLOIs2/1LluN5+Ik+qR3v
vPTC201xyTCFwGRi66bG9uzAlDGaKs1NSAZanSxFgLxnljT1DRbgRKLjXTujFtrp
ZBuqIZdbNsBapWHPoK8/Uz6y2Bg2CZXzM+6/uUxdaXMAmObuCxcnsLqrSuQcoFbO
KVf1l3jIKmD3M3gyHh2u80PXEToU8XFZHfKOrnOEfmf+kzNBuqlzr10mI+yxIFUX
KuULuoEEjkeAiHgYjf1yDNHzap95Wk3+1+YNWh7cZZL8AYpt1DWYi/baU64g1cXN
k0DbxpBhVTUxb9KkxOnKLQ9msMZ3w8W0P7mBnfZfxN1u0+vu4DNu8cZxi1myIfwF
LqIKafe6Ts77DIme9tJQZzKyAQ2t8TTJdxmVi8xcumRqleehnLfmHdG5lNUhyNXY
4TcJJNeL5XR7N6Li5ATIqo+D2PEXd1CL1qQOq45i0PKa21dEzTX3SgRiRwYlTvUd
v2UHHcRJvTjnsYcmWhOYYnVb6FbI9F/YHNdD9dt40oHnIHFaMulv1TzVBEyPyCP9
RcWYvM4ZJEJPpWIGV+h49wxpebaN0T4fcA8HCt/TisOlkhxI5gJcAFavqBj8kngx
2KwBNgfVUUIUgaxg+xaNpw0JQNS7p4e4Nad8iV4usM/z5x75gCMsOumne8bANYr6
4yYWDGfXPOf1fepd7faWfgXwaXCchx2a2XTmIXj4cFuGZgPps7SmmNcbEvE46sRN
AQDmcXoub/+5if6MOEoIwHvfnNBHTMyaH8RrRk92PjlB2C3SUfO1m74jrFnA3IcR
K4SYpc69oKcMyAaV3OYiLDXdqGjq3o6WEp6HBy122DvsCQZZMxtNcr3u0z7ypbXH
VohNYB76bFHUxxF9lFER2VTjoTaw5LprTvJV6aDvAWb3offRZKZglhJ02f5JlQkS
XB+Z/R24ne3ouMvdykLndNtYLMxVYPsqZ6rO8gsukkuxYejAs75Wpl8N6ypTCtgu
xeMz3rB6yeHZx8OBAV0yvlhn/b9xHwPuwENM9GbVkz5jQJbP37IAX4OL2wU1BLM3
gCjIEq2qQn4r2MVvmq6RdNFCusP6vEeZ81mqWvbpX/s2ZUehJNVotT2twLXKfj2Z
znm6JVpsi/IFjhHT3QNa3RUAVJ1LlgVbfIjbwY0HhLuUe4CSJhsgRr2AQR6VYdqb
RVdNeGwx8Tuzcgf8gPj3KtA8sDvn+1JCOnuMHOdsB9kzf0StmPnb8pWsu5Kl2Oky
SRsCCzZpDVlBLetHfxJ1JIcMRZ627fVU5zuKkH0/MxCzRmgDQHmUeU0DYzN/YTU/
kl7vpcUCm9DV9uzqAye7Fhzw95Q3STA3p78ArbzhySPKPWdM/ygu08xN2oIWFCHq
q53fDydeQ6F8VM/zAInFKz4/0jNdodqrJ8/5ZBwElrAZme54aMvxpt9UXE92026f
Q94kX9UjJ6HOvRyBlgCZfoMmgPfj9CxRZerzWySSd4DnpjhuLx1ryG/h6mxOE+w0
Eiv8BjYr5QqbbhmeN3/i9CTZmrjXSIwpTH2j2RUh8uk5Mt1ksf8AmTUd+4TDfMBh
+MV8YvY0elHBUe8PV9N0tpJpczabr+wdzcTIVyYmgBJGuxk8uhntz6O3bRcYV9UN
zBdIzFwBFbzGPJnz7yxKdlCmufMahu3V5TpBDFO4HnN7ZRa/NnNdVn9KZIDW1Qv+
/PM3H9CUEib38J5Kh7DcHIVUDC//O6zpKA+whO/Ds9uS+h9+l49Zzo/iS8g4B+7r
xbJQOeglWT/0y8T5Pxs+T/sX4VWTjs5oBuLnhRpokPLg+QY0fKeH4VqODeOPjvV+
niopXQENZ03SQnoWt11sKKgqveOK4ndB4Y5p1uk4ueWm73JceJxcmlBqXb8zQpDF
0F3LGzKMM1VZpdZrkWFwbq6G9VfS8HzXn2Cx2D8a3TolRJe7MRUtaB05Jgw9ipSb
AYsCG4vEa7yS7HDeqSw02sQ28UKz+4xe8+JyH71PLs6xe7DgHSRLOLiUGhkfRq4G
ZJYFesWGpVCbpnTeYz4l8ephWu3+pH/U0+wkx73wkIETUSy0plnyhWeM94w3gR1c
8lYQYTV0WtKqtKqWxmE+SdqpR+udxBXIEdGsDXtGUumWL781NnhcOrnEwxmFP+20
uTmZDVp5EMIGXnNL1MNQ9EkEzqeaoVamvYFKHVmyduWdjba1hl+BxXhqNBy7l44d
+0VejnqOQljZbhxf3NHqW8bWWiiASb9ma9XMzEBF56NslIz3tIB5JwmPJC+/Qks9
KC/yiMI+gr1aspZtcOWQ24m4U0WrxAJCwo+NxkVXSs3jeh6fa+v1+0IZn+72BK9G
4FcVWd6D7Sc/t7KVok4sF+p9obTWMifqT7ewILz71AVq+JXgJn9H8QJWbwkhHV2q
j7XaXUxhgFQESDiADbwpss1ZRshPw1hdiwPCwei+XYLIPC59eH14+4rtq4s6ZeV8
akKLSPxglBGHo//yer0FM4dbhd4VFwz1hpE8nrD2IKkTHnFGbMRKxVRNJC+SlYGV
7SH+TfJh/WEpJcQ/ZDf34JC6wV1kucqFGisbwLAz92eMTFGaIMoZWyGSXTz26+W8
itIjAaQfDzY4og3bgt3krdijAusORMeOn204nEErqFSkh6VkXYTBJOmJPor+93u4
R1xJ3/glOsOySGiKB2zeQQBMZ/OAqvkG6ZghBV5xECwg4K8tY3fnhhcNKGeJqnYQ
LrOZ8Nx7ZnjMVrrtqdEBOQe5iWHvy6xEg6erir/sK6NKVlyWEzhMInVj/uX+ye07
R/ap81Ji/bR+6vTZ1BmPV22kAOmXbV8YmiPlWun0BQpZuGSlMHw5CQKr1SPNX8HB
dkvaucAUkDGcr2Y5M6/zluPjDEccqR9CykNFfL9sZg/3dg2Sw09g5hIZ+EtczKQl
FBlfBTZ8tEO4gAJz3QZkMzIYJdOQ9xbFF+2JphBj+fpxULvGwSlUUxwzLlFGHVDP
lWiqqzT5G0aGv4oYwjZfRiFeZjzyXpHreQGdaFTbbeMGZfr5SwOK1xAWs0QErwMS
5sKsH/Q9mEl4XGd+Q8H4ORo5rMPVfnCENr7Vo2Yw/AI8x4oAZyD47OHzrCQtj0Np
aLyjX4wJJgR4sFO/7uBeUFRe5kryPnlmgVwaIuUbuYEfVOWDGv7vieyemW2ug/ph
nnh+T/gAdFsMWb2JhogmKJ+iiyjTBLZwQDvPnwEnPXLl7cOKTijgWZW18pPgtdai
IADuXOphSw/0wf8UT20fYzMYcGaRS5UTDMKnEx5gbDAG6CZO/zzit5MTsKJFA/Pp
4hNq553x+it4sGJgVA9EtG/eEry7SaGvjs8EG0MTpdG7yfbrNj8c6WPl55Wm2Cb1
+yAUikXOF6q1w62mzCpFVGyyvlAa37yKGa3aHuQFUrlVqSQVXQJzYgxG+PCNPRIT
JQZgDpxU9hS5q//mT9NYPpIRvmMpC8NulWPAi+Nr/U9LAvxoSYBJ8hvyX54YJvvP
qlaQJ6TFWVPgEhGLf/546LS9hTiueHjY2HLiUf17Speo9fCoTN6InVwIkFU6IILx
Tj/WegKSX80/vuRFyqE7/mCzECs7krt0qu6+5xni84+BrNcgGFcLDaN0SjpzxmzX
j6LKJ4wF+325Cd8d2BRhZABVnHgyz1ikeslbFhNtUcvq3mpUcG8YJOQYfJ3Z2Wtb
q4Ll39XsD74hwjOyW6wuuTEgswp/dMBb0ge1/rv8VCPLAHDZhwP6WnShP+v61cvE
fzYkG5idzBJJLGREtLjZUMaDO2rlV7liyc2HeRmijlCwzz+jUvG7QhfmvZABF8ub
ZGkbeFCOLQTOIPidOHbHvbK96j/UcqCF/8C+ayfdIEL+xyCW5LjLeH36lhzdWyHE
Vn0cmbfbKZqDO/EBMzeSMVvdSzlTYoVDgZYifpeQ01EsWRVSUfaDFqFPSO77VrNt
Vnibtb7Q0BtunsdeKd1bq2MnSNvokOOcVrjYbjO51hUakCqXr14KiUv+n18KRgnI
RjDr3rBv4FB7kpnIlTUlZ86verkOEv6FW9WSCuByu8f3c0exJQl1pTl8QhTjQcrg
L/70tPiLyYv1j3hETqy9dJQBGxxAfzNTzFeLz8Sc7P6FII2oUdSlTByx+baaUvFS
N8unIF+E146MkORqVL+PU8JadVQEEWqi07KG25q3vPx5Hfya1Y5nMzEUEXgzg5jA
8XnANCIhztJP4zghnWGyqJCWWW3/ndwh81Lb3WpNpJNXM0n8mC/Dd7crL5LvRI9x
Qui+sX+8bqzD51diqJQ5tBXDnHsoKhUjmP2Hn1PIJNDbXERvxlOV/YaSEz67MkFo
9lZUue6QGAzgsFLIezsjoqsBt01e66NvSX8mRTZHSiHrrx++h1CconhinTXL4zod
1mZpXVUG7/cSRhnfCh2RIRFabjnfv3KdjnfAbZZFf6f5J7Dn1yRXdsre1j33locc
T7drj5tluMcHVw3tv2nOJLbxsaNqEDi92ERh6IbRseFWyGOv4Fyi3UNL07vwpZv+
ySJZoLISsmQG1KN0VKEpe7OPKCp7dX36WJCFK6C+tGDvxWD7A9Grk34VvNThcqnb
WE1AlFH2rEp0Y45greSFDphurbdxw9DSuY8+sbmIwKCorHejKVBH3DPH9OWw6R5u
NwfhjAsaEXKHodxRjmhRBtFs5fHSRX+JrlV7MC/Hb1uTyRhsik0D2eyOby0O2cV5
+XpNXg8tAzsC9x8//0KqzqGN74q/XCRx2GZdNNDTXsrIOwiXh4UwYt958mZJnF4a
5XIU+acRY/oue6XP5BW2i+yIVlvEd4/MpuePiXM7bcJkXEFYe4fGqqxmQy2KH0Ba
/l91RLriIKQ+jaro4GRMLhesEVEvjLn9fXlSNmuqy541XRo4+C0I7BxScQTptOAo
4U7O3S5ZcSba1GC+29Q34+ZjGkl0JUpyNQtXLTPbDrjd+2udVSevQmjiltKq0Zxn
8X7f0dnkoA2FmcoNDjgagqewjj7RIDb3P8P85H9z33EG/gwbXbI3hEZ0Jgd+0ngH
DpWqhbYq9LL3bGgYRCd3JRJWJQYmwsWpVtt7YgNa3p4MER/u/Jutxn+TPEQc6WLs
Egp6b5xUJteaGU/nvfmcHESPHCKom9qgTL9/tyRIz9/sQiAPr7RK0+AdJQEQt39u
uYV+Ba2X+mbz5uNgiowEmo01U1Wb3CaO7nXbj4n5KD00YmjxZEaPqAzITZfc3vqg
Q0J9VN8Qs60t7i/5soeeQb/zHjZ1h9Yt53bStwsRmRTEGiGYxuGP6oBvnXMuEHD5
q9kVEsJjZ+NZGGZ8BRT3TuXvAF9C2OnfgwoRJ/xYQbk6hZikiNRDZd01Mhz8Mjok
L+DACx+/EREd36F7zMCB0nM8XO5YaCnt5dY6OxThgcr6+42g+qZ20iF5eik5PH07
+x0l/1kqWHft9G8QZnZItp0SzrXhJEcqGNC0svD51m/Uoh9zcs/UOde5Yyvta47Q
VauDVSZOtlrxH76RZDKCKR0ufvV9QiVdywKWY8Fpifzs0MYYxrZxwWjFQ8QJs+3P
V5ptKMyRC2/fscPN3Iz8JtAUR57Yt7Ul4BoB6JIo1fJNyPrYbG1t+r27NlId8eHz
hBmjXHTZaXRZCMlyqarEcBK/wLA5Y8OiZO/LKvLpIDLDj7KLuxt1dLS56eLdMlDm
t6/SegxwchP3ElzenlRRENaEH9vugajADLAwuoAzucUl14nOs/vyWvfrVHqVmV/w
afZ68d5LZVBmHzPsnr0SBz7WTqXEiJXmrILUOprZ7YUeisXzFfxndyKoKkRoxByX
ZJRxmrWpmGjB/8a3TA5asmCO2PFdUFiEdsJyRRuaaMEfyeAuazvGoyrG81ATcikg
br+H0O30W26V+YYtWtgGI5zJ2l8d6QEO3qhlSvdwVdkD7zBTSpShqTpHMvdKtRET
1Hz+JlvZwTgIvguXiRQjIkT9kQc/A1CoPoQVov+FaV42Wfd28FxRaY3NLAsq0gie
6wf6rbOCjpbMJkZU+MK4j4423YuOBW02+Cu2D/o/T1mySUOB4yJQLNQGo4jkv0u9
H3CnNmrtheUNjygsuhh3ImVqngxseRStF9kRlnj/SV41A1nRvc00h/hwCe0rNRt5
RpHEvPYhKJgEkRBywD7hXxWaTiUKOIxXeU1iuePaAXUTPENhfRROMIpQrxNRrEi4
lF0h+C+ZaFtoHWyOeOHpuse3ja2Wj+rbzXAkrTEPnL18knR4ezvsNO+mpOINZPfA
9z6HdZx9mAQPvcvAtHS7EP9dGDLeopBNVbr6TttmSBAsffT4/10Rf2J9HICKjx0A
uLRqfg9lm8d4mcTON3NDxcvDeiVVR9jZyd9o9k1SVId+XXiGfFd9P9q1PlQiJaKx
ZjY0nVhCshAShvl7frv5R+hQx6ywMd4PLHisMBdXFCUgWFHmetj6/W+StAAh8MOq
B9U4MmhBsihFKNZrqFxDraTYw14BPUWfJYzzxLgz04Eyx/N8pyO5TMrbOwdoJiLQ
QV6Vo8F6ChyPBObpu4d5BL3KOHAt8BvR5zdZwRhGaJgAfFUlToEwt//T9B/dppjJ
1CZTKEU85DPz2E67ojRGqz4dkxS0kQNNQzCuIkrODdfR3AAvWEXHD79sQ/pKBIjG
51Tfej1UY6WUp0LT5a9c4dp4iP1sloRZ+BjdaKxMUIsxy2ZTZAGGFssfE7q2FvNQ
62t6EKGrzlpDoS4QRAX0Ly9elK9c/o4JMX0ZmhAYGvRHvoglPGtvs/YIK5DP4VEt
kQMtZv+XoHCrkUIUFM0QgAjG94EyAmkS0Ium5GQ5nGwYtk7fhxrE0IMaKT+dc4mf
nMBhMSLdbVMiroDTtkW58+mpbVz3I0KeX4vLPW2OQw74T47tkwZjEHjm1QeffJI/
izBmsOkXXDcgL9vHyana0Q5wjh7o78P7Q8W1mqWdm1IyUsNQAIMmgX+AwtITZWw2
6/TVpv4OFgMJX9REKtbly70bAog8tnGhw+D92s6rklRDskvzi3T1vAKku0ZFVPjD
JyZ6SGGtV7wWz3QlE18aSLhynEu94KZq0WQxDVajneCScI6ktG/erDnCua4UO4FV
mXYdidAB4ATvLFaQEsuzEU57JdLeEK35nN4HA60thWSXsdoOVPh5Do756SuQIZ4u
fGdou4vL00aJt/1MWYkXq1G52tQftzJIxCUyDalYjPj8W+8/GNp6aOI6D2afXG3g
+gDo8yhfEbRs56mpjRMt7mwrPOiW0Zzu8ws50FjPzc8r3/jTEJyBMR0ZJTCgkxOa
UUSjbkcZidqlt8DIUwpyd0wUeprFN2CcU3T+ekVWvUuU0i0/iI/BxGms6olEt9HV
XsnsR8OHZ5ZmaGbbWRBcFMcnz9VqSXt5h93QH3eW8w7jcaavQRjxwpCUYg9rGA7P
JOXcKoNZduuw0snxQj+NpLr7n1HCWFxnq33yPH7pvf4xWVTDWwiwbf9E+byZ05DD
vbqiAbCHhnFFzaPKpVjAXbF1pdnOevyfVpjpQD0b/YoXxIuT2tAO4LtVNKK6VBc9
fyY8dlbrYj4Q235x/z3iiKMJ4CJ5AgsxnyHT7UUEX4Aj17phWZukkWAiGEzSlq9W
M4oKevsX8ZR0f2NCPgirpCEUz9NSTrD6WOEi5vagZvNyIN+q/myFL+fC3QPFnQHw
6tBpfHZonX1MxXHFB2S8HIS+kxI5xCkeWNSnX5KeRdRCQPZwaGcQBL5uzlH8hHJ/
mnzN5LqKm2F3P+KIuazoLaFLAGp9JGNt4IgomFnD6r8Rc3Yqt3nSL4Eo3EfB0lCs
/vCYn6mCxkstYlest6guJ3R85Pf+SEIHIA2iGQU3ldoCAa5P+7AgIPRZh6a+bBnj
Ksxplm+ZQPy5x1YV3XzDHW20LjpT46e5XHK62bP4WeBqMHrmnaFViE1n5EabIx3A
D7pikG5qre88EfpFm9/IhAvc7L1MBq6zuWDHlC6nzMAwi1rk4SGnw1bcSbySYlkw
YXzytK4kSm1iaET5BbCZ6944/mEyuzR1e0jsf8pJ6gEx9y6YDYu3PQJZ4DrcizbZ
XSaxgzVaTFDFMXal2KW3eRi5rI26eh0iWdZli3Xd5Vp7MiDl88vxp6reHTK/Abfw
2wJ+ka7YTwu0Zj3SMW2cbpmT35M1WWQuCuHYO1HlJ/ePbT/TPdJuPEgYGaIAklvD
wsOyO62LM9MwKEsCQ9QtphNEvyR8U+IOM4jE2fLyS4Omj8iJDpK9mEQdk1xeFym9
rw4sS2FMI2P9e0EDpF1p3YupSH9ZBN2fzUvB7poHTvB3/QPHEXCEbxVrV7gdvVh4
VIbAcVdkP9I3VWgPD6lZMP1s79Cz7v9vqwGm0HtdfkPQCsw1Oooi1jSZCrlpdLsm
eqscy4xKUEqeqqzkMPVwWUuBEMBH6UGMKeXHkkZQc6wucBRr1LM0jMV6N/dzxrZg
KkPoRk4TqyNUPU/9Vil1G/dfmdEFR3EjT5Nfpwdz2JeMrzPIgYEql+kegRmNXc6z
IlGq7vD0VrcvWcwFuNsE5nY7RfkbpoEYVPBc/NKiAFv5u33whrePooPFN6zoD7gv
A6loNU+irvgDlTqSkrvQuMLfVa+Aee6t3GD5PoR539wMnSFN9Gzw9+5tnl4x1ywH
EZnlO40jvDUyFLe/9vdPUJ5XwxUPQhVPWMAmnRBinZfVZKvqnQLZvUSkeNPixFYL
+xwkfzB72DZCOaVixH9V7s4S8txMx+lb6sP9IavqI9Juw5yD02ZTy3BFmcjh7sAs
fMisSV7niFZrSLChh+i4v7nu9DYpVN0Nb8NBQM3z7UvS20Mtz+HfpPrk6DIFcVJw
1pNRmfuU5S8am2Z5PRXuO7MJvwxcGKUIO9L4kqL6KKlLMyTdorAGfTcvQu0ELo+2
PH3TXX4bj3ae4IwkjMsXSX2qwTwsu9gu/vPuti8c2CUAK1mYq5KXd+pBTVPyQ1j/
88yTmyrz0j1AUY1UrUDiKXYjd+a1GVLuV1QHOqR6QImILpSTlkxWpn0vJZJkGRUp
cF2fOoEHmbM8XljLaLZrG+0mMDcwVDf0SFArkgRttaDJgLxd5ibzDwpNLjj/bUyb
oJSBIyA2PmlFowbNWcSnARIj9v3cV1dicRTbBKbUlTpR9+e3ChYSXdinc/b7gyKB
IWR4IWPBfGnQeXBPzAWJRts7hEvwpJtaA5pPFv5w9g0VvElWVVniDT56YmjgydaJ
p/SvSH+1ZoQ9IgQBfzfUXAYlz+R6R++vOIhKSQjvsBtI5K3LyP7Gpwwzc9y5J+Co
ZSX1b/E6s8xe+xw+su6vIZwpvohapPVxJ6adXFfJ9Akv+sk9R0b3fiHqmemF1o3f
sRb1bCd0o3AsDTdKCIc20/bbXOA585AJIO4peaarBrRXJUJMIwaL8R7ZejWHvFJr
cj0Xq1ATw2pxOBNklFQtkhS15/tTe9ryhDLenEbzimin59DICJUehHt56AYS6VVT
UCTpmixSsGisyUv1dTnPmjdO4j02zZLkw+YWDilmMnfYm3h3xBcHAsYWwgf8yS5r
NLPk2aJMQnEspPjV10iqbtv6emNoiGVqI8BI2UfJ0fCczngl5GY621GLkP2kdU8+
bfr8dwItpEXqJ7r4E4UFXASI8w+4u4OI6w1QsskOrbPmY/fXXB6VWoQtGWQz4eOt
2SSl8y74GM2rAKb9j3/N3CNjP5WIS66umsHFhFr5Bp8WYcsF4BZ/UavLh5NYG6ii
7zlM4Sw94QDMcax7+bTzRVVtxvyHn4SwoVou2T6dTL1XpxBh3Cy9qvbB0cbiFuNU
+VT24wXYP62c9r7GN6ZgJ0BPyCiTIw1dC6QTR4u14lCPQJU5yNaH5ocDnveDgEzg
l9C9vpFoagSW9JWIDqE/Tspl5QT0PIUkX0uKnwMVa9tnC7QxPT+jLT01G651UOBA
dw1q1tLukwkjRI4AZ08j3dl2CYkbbBDTq+tsFx2/Qte1gCnn9lhAsWVhC0T7oUZi
3+bNVTfk9ncBje2zCIOoYtKa9moEjlR6yuIeDkuJMfSFmjcqdoWe9OK/qyW2cZqA
VHEEOEci+5wnUL/E9f4OkHvWgTv8yrhIGOZUno84zcyXn3p3S2HO4o04/+PyqOSM
0TXp1QepwWNhm6wBa8vDcbsN4B2Ox+CjhaLZSbHOKbbN99kaF8raQrmyL97Q+ZJy
zjmcU7bbm4XoMyO4+xePX0kRuATCcXu5hhV5WNxrWpKin/WyCywz+s+ACWOGWuDp
yEkZBRfEroPsoQlHzH8maOeL9GYNvtncLLDYirVWWE5o8XuSp3rIU8b/otam9XQT
0JrJMHOvrRVda3Rc133zA7BMsxJpmnGGsBg1dC6tpSdspdb4GCTD3WnfsfDdWHe3
pGT5/xsBfigfs9GlBtePz8lMyHKfR7s8gmP7nKXCdxIbKNw4/CLPNKgW6rNcSkXm
D2F8R+lBPXQ7v6VpQcmN1SRvdJR5zYywfF7yAy1HdUXo0B/lxBmjJ66EMREixAXK
tCbXhtl5vzEHt5rf5OGXbamNOM/PFkaBCtBgSgQ2KSA5NsXP5uYOMvHFiahcOG4M
O5d4kzprC+UFKzSnyEckQHNzhFGkmKiyK4ALiMjvSGJccMbmqB71ArM3/kMYwimt
xCyBjD9W5mMRx8iyNTvb4VKb55U8dl3TT8OpL4J91RaEro43NLRgD/RIfAhLNVm7
GLw7y4qcP1ijIfXRTHyNNjfPkRCBPI4CZB2A6Vh7+3UbKbzq5MDQIzGkv0JUiUqq
jyW8kd4UtA/AKGYE0KCFYgko3H0LEtaDuQj62GA6h/Mgj8HaWs1h3qBwVXslXSaS
CD6ch+rROAQUV5r02fzmCliTALp7ylipp7I6Vk3AwBX9OXy7RSxdwuIXp98oczHf
aFAVcPjQ0lag7NGNMC4bSVWt0dBq0z3Dx7iXET9Vzpk2H7v4g731smWSY+WAGocb
e6lQ7FyKSpAoBylL9K7hpyhwOePYmxCNN7l7Ud8YgE+SuRKRf70mLaaDZ/94Q9/B
qw5mwpm4k/jgHLGkFsgGL9CIddENlcwaLJZKRuegP7SpGrBcirQUljfrhxLtv3tx
3D0roIHsaJgiQduLRYQ577rEgYAV4+lr+WWv9gq0ZBW8GKoX6gEHtV3b9cdkJPvJ
vHhHd0kDjIt97mHKXt0OKpNO6DXnM60MH2yERLLz+f1Yy3ISytTo45uZ7ubaOAgJ
qLTSUc/BXIf2RHVUEUlLFYfPPEF/RN8oi6OC0I9tPoC9ly1baUJy9Eb/DcqzNDn4
I6+oZWq/Fuwhd8FzirHV0Nul7QFzL5BYvlYfOIeD1cRb6H26guC0qjEfIfYYrjHZ
3HI50RcI7E2og6jrbnPQ8w555flHIkuYuDsx0g36IF9KjGO9G1yngiq3LhaXngwg
MafavT9LADLV/TLyOAvlQfIXGpd2HuXPtb81ZZ7UAdZCl/TEnWIr2/CDzEU+3L43
NxILd8F+oS4fnwBRLqQSuuR4Rsh8tCCL/yCkPpOBVSuDmjfiTQZb5+P53CD9/qxg
mXC6e/MT/a3hiRxBxCR0R6p2FwppCgQPOVU5W46u49YlUpl18m6y7BsOKeZ1nWCL
t6hP4PBTeD5C81HAEHK8IVWrYbu6fJqj1lzTJDkC1VejxARO/KfZq4cIhnyWG+u0
HrI21hUxpKRNnWbrNHtKphyD8xo37T4pvsEfJHSSqfCfvfdoXxErJPZhwsLWQ2od
eWG/HIZfrOM6p/dO3Wj4N9SNQcROrjMvxvjP8Zsdns26SLL77JfVlc17b+kCMpOl
O6jnyQr4z6lg7OJbpiy6HeSDFrIPIFRv3xXlyW2Lb6qSGwJS1vARREV8ZvUsEatf
v95TuN8VPFsRZV4Tw+hAf5yBo4LSD7OjIbrkilHLKtVQyqzdFuSPCvpkmuYu0tgd
EJ4ecNqNSzuBlLiwxbr/5TbAc6PUXeFlvwzV90WaR2bPv0cVIANwmPDNwoyM5XQv
LOFrHtDM95K04QZt9RHYaunpjUGSq1KTmIie9UsQ6GUL8oFiGeAQJz3b1Mhiv4a8
b0lcllx0u0zFkOe5FB5Q0qHlCn0iqTGSFLOakcPWGaMtOspcD7oAtUjrkzUxYnQf
BhT4Q/pmNe0TCjcGpXI5I1n9EOiSDNEfdmM31ji+YhtdmSlLEJpiFKMmCOEeMpfD
z8J0KrgFqjYV/A/INFNuVBnRSpQC+yTXFhui5z7KWwY8eGYRXliT+Jn98c7lzpoQ
UIUjugTx4EBFG5zFcQ1s3ZAS2jvgq5dWJyHu7OYrHLZSuqWzVWA2V/FKlfrHplZd
hfba9WQPb3/bpnm6jY7CHo/q015m1+r6qoe1MXZ7S+dtSelsM2qrhuXRsrPjsfXm
hHvxfMDcD0CPGMEZTXEU+99T/X4Pcil0aDDf46P3BzEp7OM1hAeERU4dqrKkLx4/
FvyrEfgqT/nVvmJZJZlOPQRAk7S12cuEY3GR6vaslTRSbdjX1ACPsDHwRBMANre6
73HEofFMCiHMOhButqZoRwNZY5Tq580JEKkbmzWIh8PD/c7TOMOMhiDAEu4AsX9x
FlNqJjKgVkSjr4jVjRblznPm0V9c3vaQwEkdt376VlnqiionUU2itnUrqyjUTYgP
1VLIT8GcDYeXC3nI1DctiZapyTN/CyzyUJWhxUJSqBM5fTxeBmDHeTDaqFKdDLZS
lYW60A8vphAqN2/Rj1ZV2t5qVYB1sd2pJheCKOIZIy32IYgqhJ4AkLJpB0aMuXF1
D3Xnj1ms3TiJzgw0z/9qj0W3wOIPYVc1QaDsf3kq/l35nHtSCwTYBgTyZMGBfqpD
dNzDDsOtJyXfLM1pJ8j04S4hiEKq4WPGyfiohHpt6Kv1DDMScym1T8Tm4YfZN2gD
aw1yAvyh2JgAROZbaYS8Fnlm5E0xphTBws+TYooMPKtHyLgzgtYxoR4Nsd04jSpP
HuroWX38Ia4hQQVxTW2RvvkakSyFhDPbgBhiJdXLeB+yKgB6nJgoQKSS5WZTr3T3
sVqfUZLFkDCDGGEe5Og0xjxTsu307g6Hk3z6RulzgoMS+bwkSye5JLFUky+3Ut7o
qu53nc2yRBW7c5lxahdUWPlq1VweK2uiqidSB0TVcb6Ba1nA/wgT2PShIkNVKw11
m9re9G0ANRnktv4WmGS2jnwPh773d87B52Bl5dys8EjhUNBJMsibA2/9MH1i+EPD
JRsRRDQ+fPoRgp4EgXIFEoCwDQ+B3akQ+djQgHt8zFlOlJWzuS58CfoRaa1nTPNG
nZ0T2kNzf7S7A1aVVjvQpdUCg+QFZ9UdVqhGeqjik58Kb2Ve/U4LXYTJqxUgFKkv
j53eH4LpwRR7mJRWiful83yL2dQ7rluWvM3gLO0lz90sBpNXpDNWzw9R9VsOWa8l
8vYIbS8kBvhsMCCiIbaSExrQ/mqWJ8S69xt3CsQA8HzptKk7tJcdZrpJP0GZa+Uy
C9Db0rtzPAQma1hEHCw5MTZdkhrV3HRl9ealHPobjjc9FIk4npcFEgcWON/oBK7a
E8ssF3TPI1+MGMRSFpIyb9FuU9mJwesPmOGWmm3efOIKrgTp4xH7y/OXckBg6RI6
0TvL7g12r4uZ5k8T3f4dhx9Wk7s1VAjxUjC2/hfircoqOcr1U0ERfmbcCUHx7Ygp
ECIe4alDeaURgTpw0teSRLyv14885j982HTz+2pCJMPYzWQqsrvFvY6irQB/A3Ua
KoMI9O5EGW778qbT/4nOeN+VG9NnSPUbvFLZc8u+WE6pF2QoMl47QKrB2Cjc67os
Nthr/Hq34dMsWZXCZan+6Ayzfp8msC7+RM+Y79rfsyGGnHEAX/X6sSwnkShjzZ0e
X6jj/VMHN+qBSefS2Py+tUeEP82D7p336pOsZXs45W45VwH1UKhaDLumItik9MZ1
cT1sMOKMS/AvuG/LmEuSlLk9AdZEBv4MLeB4CikKa6vx/Qh3coduhkJk47T3xQbE
oDNTEa6pzmMh5PNBLj57qnOPJJq6eR0Y9ymM4rwgv62kEzOmArhAMfaG3aKglpWH
AEhTkqXBh2pKffyq5TDOhRDDgMXd1DCp8ie1G0lIBfQ4zjRJtnaIq26iNWKnHYhn
rpOO+pC6BKBu7jK/GCQ81nTaq8rmqfct5AsyWxx0fiB85/U2/XRBCTB8G5ny6VS4
Ke27xP+6uLzf14WkKoaxIlYuWjYquZqrrRDK5UMG8h/vs96il/xLuZxtdRVVX8jh
nZ2r1JCahEkOsK87mOxSKxjpr/GakYDvu98h8/yP4dynqrTJrv0HfGuZPDnZB/W5
HbWhw/DVhORo2GC+ypWQ+Oygcbk7BDfj3Wabh3kCFHTjJWqkiFsLhNftGz7OGLEY
mvWDdhmliv4rD3L2Zmiuk+QN5juYYkkfvhc41VVgb2IJwAH1TKoodtk2nt/gR+F5
IkDW1Ofom/4LJm6PSz3NuODVbC4ZW9yTOXrrBLUB9HMTGgmcL/VktwOkuZVUvplu
9u0Ne5RMkihavS5BaDB3yfCLexc4kCT9axNdUULTCtWOT3W8MeucoMi7NH1h9DIs
I7uONcr8wV1f5z5Sod3Bcf+oxqw5uFZjY9tv5yvF10Vy9Sse2mcVs7+ZzM8Iqx4h
EXnAAhZDL3lHe9/OYboEqjFqjmU+JUoG48WCXmfhaGz9wp0o35Ri17XxO4RO267y
JYbphETtAX3TC9f0VBVyQsgcuIE1Qz6FCmRqbeCo8LPhV5hrgfOFOXHpwTI4BlBk
tjay+Qv6+R6LBFpHL6VaNbLUVXccc1ACmeMQODTHNpG7BOn322vWw/HpvlAfUk1Y
AKE/5qUg0anMRvUex1Q1DI65Tod0nmizHsWQnGYkdRc3Q9uMRY3KRRdaXnbHmBtn
N9klZD/B/pBkliDRdn8PUDLmftC0xC58HDSaEknX/rgXSUhRSVDv+sm+BS5eQOzr
CCAVJ8s6h5Soyl5tJ490jNL+pIp398f84KXpnWNnFG6+ww8d0Y+MamDEoNv8Hklv
iy1lSIstnuvBvCXkkYbO3b+fmHKjAy8O+9lUDKlHagLTaPEXv9nZW3crB3grrO+a
j6Lrq+d9PItel9iWJU1wFNmRN3O9N7Rffet7b0/2h5lFDevy0nG9MFYvGm3Bc5vK
l/veJZMdtoV3ndcAkurxq4RoCKdIOk9Dk4qL/xHQoA+Mp8wf952/dpHFcZPeTyao
/797XarccRgEWax70WJ+6tejHUCevcyB40KBSTZvHIfUTYFIdZ7cXpY3qXrfjpMB
CHi1eaxH2sjMJI2jjEIHjnuT0o0VSR5XZyVlASxsf4sTYMzhnYC3QU0sPULrpWmq
oHdIB1BfAZd7e3WBdodb3QbKeYD5z5Y40qn27OS0vbqYh6hCM1vqciFP5PKWd6vu
iOEsPqULLrsIRB0yssPm3flSlpE3jnJ6La+JbkN8kVo5PlRKbGfQS/498tM1AnQ7
4kYehgTiQfJhdo0QIkObRD20zFfn82gzE6cMDGLupOScsF2NZs05T/UIdiTUT2Kx
Ay17PzK2DAwR7K7YcExUsx9LgEFwaE+r7Uq3dok24/OBE7M1AlO0T8CDqU08MQSQ
5eO/ercwjI94mDb1lqRIQcvQznwokHcyxwqcHQ4urrngdVoswgXK7m9feevEBfrO
QiAYy8guyi2N3E6OQQkC0WMP4n6drf+iPu8HX0YxohuaXQ3GE6QGiCfIDqt0OUmR
oN4kGvsvGvJ7GpVqf6zK/Llxtg41YfZoz6Prn52DkjyV3GHL/doZZPqXib4eP03b
mRCzm0jY1AOQuNkmmVW6UHgz+tebZUHioPenahjd9XakuM+gfLiPtYsy4UaUvxM5
1sig5AGDdavJRo/ANtqnDS+49QHJ/vaR9Zj5isZIv1e4byPFROALitloUIOLu92n
EBPonvYzyy23MoEqM0zYrqbl8sexdSKcHhrDRcGjhVNtFje9RIepOWBbtEyOaWmz
h8+sjkIeB53WhC3nwgAZlfOMlTS/tlqWNjEswpS+b+rkJEUjz1nGeYzDUAneO9FA
IZHtS+UkYT3+wAtRUfF8FfYiMGgaoE71GSKuHQBIWnUwRnQUmUG2mtwstz4nNErU
wZDLTjepymgpprYxgN6iYGaj728vYTo5DapLrqQyXoW7g7kWmf8nMl2vW8y76ysD
/V0XTbnCi/ieR8muB3Ibds6urvWTsCr6IstxJpGlcn0wvWtScB3D7Na+/i03TD8e
ASOFk3x11v6DOtxDNWCBL2v/OoccqDRmUHm2eoL03tPadObgxjch/Xivk3JMI0ry
DM6E5AoPimHiCVu/udKV3/WCJrqXj3HeszTNTw/1K0D/ST7hrytIJ5bWIU1Ai+x7
LPk+Q+3+3WXP3h1f4Hhoe8TpZkBm5IZa8Xa5tdJyag5F5Vd1BQS037rPy0Spa7ZG
T2VAzKuPqmEBLIchvaCxV4JzwSV4j+RU+RykW6B74AMVXtYaZhRoF7aEtRaioSjY
IQI32VB9Rkxyl/4mFG8GIV/Ilhp778Ddc9NHUWHbmvSHdDxHgVOnIOKSs0ZeeIsc
5CyqCpox4kcVvlC36XzvCFN8Y1B7V4NDynhDWT7utIW2UCM5YV8isWMeqvyKVAg2
68bi3jmehdOiWG7MucSqMN3glrLpU6BClBXnhRGO9kG5G7Uw1XA1LQkVs3AJddau
8IVmGcfeo9YEJvB54adrl75CKdTftaT3T/6d8pkZ9JUKMcqe1Jw8cRVVuzv5+yHr
AiZ0sBZtJrRls8UPW3IVd6eMSdxTCDTo/abjG2JnJx/m0NJSNhbRwFqSAFVm8luP
5GGIpHAABKP5w3lY0ZyzK/ER7soxBi2qCqIOwTFmP5t7TJ8WhmZuPBsOACabk0Ry
mQom1X+ZpjeSXB7M+yRcHHkg2ZJqRtIocO3jS+YX/YuZWFg48gCPxZXG37Ulouua
Wo+CcYFD1AwdqhJFeTd5gccsI5mRdRKZ20wVqsSOMUJO3KRrL2OiljrQO/t+xEpG
ROrUnx5KieHz3zCnj1XRGu198hiPwW4xxFC8ZQzIhO56OVJE+3Ne+zOntwC/kCMo
DrKP/oIcN99Bkc9+GutMpWJBUnrIR7CIFxIyHquH/0H74Rvpj0ZRJg+5Ux+5weuV
XAlq1W4bBT0J0GOJc02IKshv1bxPlJgy7g22/c7WgVRYWf28j1m+G1FNkwCZn3Ff
AxEvgZSO2SS2UFHnhh849kuXNnQyHNly2YvSoXb2D0XXWHITGKZqMl7LSdeDWwvH
+yERYV2oJU4e/ntlhQUIR0TaZCK+bJIEhUAVjXzPdtpwQpIaO14fPpeWU3X55oFR
7/qLsD6VBSTpWhEswmlSdQ2ohQE9ISbSkdECbplZOuKVUAYVSluI3zbkCc3a+80Z
GCblE+6Nt0yfWGn3xR/JBloJKcT84O2jNh3Kk7N/YVg5zJonCyMqak4QjtmKg3AE
8Oof6ClXZfiXu/1WMz4IngfZaIayQW2JrK0RZqTTWNg+SuD8Ji8tyi8lMWbdSWqH
3G0uaFMjJbbiBEFduLaDYmycKSdVm5kTMYmBmak2JCiV+EN3jdiFHjQZwk1Mewr+
GCnnCLdpVf57d4OtVoQGQeFclYQ8wyZrLPgEeNUYfFAlLCJJCpska3h3EF37uU3Y
4+Ei1ti9wpPOCwG+vcQWeAtBpEgMBO7HSLVk1T2BKlWTOlouMS2GWQPVFWyjCR/S
k3G+M0XjSXVytMtTX7Zw1DmXOcTmUQu/SjmdqXJp8/bvUF7+/hsEXinJ/FuzQf3j
Xjm2mK7YKrb+tRrec+7d64aRlTTX5Yip4LU5njQHnytOBBqjBOwrpJX57sk2zIsN
Co7wjFgUDRXaymyUiqLu9y6JYUHC3rBUsL1grye+wANCJOhuYOmlYoQc18xdbrZW
P6SJCnwD9umQWt6IxLpTaLmv91ryIi+idev9jvgljiXDIN0O8YdxqJDSGqVgiv5Y
67Kamhj7yHXFEsS7AAn2ugZuBP9Y7KlqrttDTaaAEE9HNl7Xk2jAqpzk+q/rsRDV
cYORme+w92A97sjcnVtB+AXzw3wk1FX1fxJ8pvHefN2NB+jtXO3IZYmR0ZAftYZQ
y6jWYvGd//6pY8yi9xrQl2sY/SOupxxLF4HDnr1VrD33YU4zVZcgtcJY2BK8/+5p
A3+AcuAwFzznmwWg0qtdxKpYuHGPsYrCQaqkqNly/V9JS2VSnweBS8rwcqqPj4bt
pB53GdQR4q5w6IKyOU8Sy761NskTD927y0JN4i9M7k2jroYVuP+LCR3C2b7sDbpz
jLJsH1r6qcOxEqlaMDTQA7g8Ti5y9VarSCPCZOxr1g5euC8rrjio2EFdkb+3bFu8
mmC7k6zjfh8VWao7V8ZUpOKhrUnrtztywWIHOQ+1cidZYPXArXgNdUR692qibG7x
n7OfhagwhIQN/BUZOtw1cZmgg+BtFuG1j9Ov/kEcMR2VX1H/cd4YvNUU0P7cBtxF
cof3dm6b7YVJmEQ/utMVqVEUTI9Io3U18f4WG0zp1YQnxup72WJcD9xex8vKQmzE
RJryVyWOM6JkoB6WYGCQtsbDuAUqr+uAPsKlxgtBbPV1j71aGJ5Gyg3YuTvAT1ud
T72luKqgrC1MHE2/X2iSEVVpH2KjOBCFm8Cb7u19dX+0aInIBb+SAnnHFhQulCbe
U3JaE43GHy04PGTkKC8pB+lqru7Y0Uq3lJitCwT4t2IcuW9hPljKqHCJvWxoScN2
JIkFgJvNsxGakDIzpDDPHE+kjhD4mKrtkOaIcMg4wEXdC9akEMqItZvtA+LFPYEb
D6WZx111LwahDR+OoOCu9ipfhGp71uer2O6WhFZYJzJsDo3l6bvd0kMbcoyBYqyX
HUAI5uUTinKqp9NrW//RN5klrex9KZze/i+OaPAhjYSeRWZX2+Uam8EAarsRxEWk
fz/Q0P3dA08DUoKFApZepKYhK2x90lNnUdf+l/FzJl/aHC+DAgxLlFHIO5OV9tBw
PmMWUU3bO4nJUhvD2leYLrwoSrGi+A4rg3Gx9JXRmGPx7JyEEidtGF1sN0s3koMi
GX6CIsYPaGL5BwjadvXwaDXkWHlBse1iyXLp7uu8xNjeforcd9GRbRMHMpcN4y8Y
Jj6bZ6+gWGpJqXAhsKNoiLCz6ZVmeWl9IoL6tYTjtmOYgysxsOVH++/iGTOFkU3o
DMPgsHxfLmC7+SJA7KPwrM9nwGHCrAv2aI0PeF0OnwyDp1YQQWCTfyeVPMcYJTAe
EALFHn2HoaR4EBl1eoeFVpWNxiswPIeJI3GyqSHIKpe8y+ag/Dox2FQI+E2nP9eO
WmpLX8RPaH0nRtresveIHEoDXgZJMWhogQsF4Gn2Bk/WC0luyjXmYqT5sI8QCqtS
uUoTO2jmxXL5FJ813TDvGoeRw7riJWLevTTEaFfNGhEB+AxaeGlZhmSh4dt67ftx
bFf0pX/6h0WKpgdMxe37vATYl4L3aRj9AlO5BonZGFtehgaIAAgqB3yTl4NWpTmp
If/Rx2r47d6j4eNJ3s7bxrz7/OwFxtv0iq+2nuyHsWXvw9B5Caz1ErEGWRNhVTvg
SN2iCFdFL6GbcGXggn2pqde1rrMThOJbK8p2Ii+YaUaLAgex9pSM6igN2qq2s6xP
+jzOmpBDezsPxXJNs5cbur9jCbkQ9kpLb3w+sK1yl7UPsOwtk6NH5OnTOHpjiBp9
CsTTDq9eFLXUBeC3Mp6JSOoYuorILLsoDr7VepK90hGCESdYzn09obOGotfPwR38
4DciVboTYxQTDughmq6LsGF2R0rBKd5k6Z/LNHLJcAVlnfoX99paibV7FxffUVez
tiFuJC3ow3/VbsJme0ACwyzc7WYc8/zhWwl3b7LjcItpP0NfBeYhJJCjZpil8bja
MyHgAljRf/C8Ted6LJEstNCiSPdVTrxa1IT/PfM93+TaKs3wX6/HToqJF0uaBwqP
Vzli8xaTQ+KY6eB/fnvYZjoM08K/veQAESR+TM6yLCc5DjPq2AGUsgBXVv6vaOmn
OX7U3VQMHQlO6DAd5QnoTElkTkf8MblSSCne0yzGSG3k4DwTj4I0bb2tvvNltpJc
ExvCQ5hjT6nIJ4pJHV6dYsH2OX/xNphfa4G7vHSbkjaNZUPqfW86MLMixzDwXVXb
xx3JeQCJG3HYCBThMYCW5NhRQAT+lTJPQTtOn5eUdBZAM/g9E7YEzHXg0NgvV9C0
pbGMKHs38FSk1HRGUSDoi73usrWQR9aZMBubsB5I8UNpr9YA4VjAtW5g/SJOOq2l
GgBJD+2tfH4vHjKwC5/1ZiOM+RduYDWARlbvFPqrN3NkEsdQ6q1WqrljN+QXUZhS
eVZzLXrJoOZsrrlQFKZVBxBOAe7Qpk2AIM5/10EG9kgDPOyshk6aU+nx3+lzYDn4
PF2p0fUoMGrxX0KATgmNyD1Ed92BVt4G4M/eNi7COvcXmvcdSeemRuEbqtHEGKvV
KgH6mQZV25F8FFLAPCK/WJUUsyFfsaJ1Lj9wSAo/s4I1QEQRh5plmiktYAKkJcz6
5Jkq3uk3ovwz06Y6obsZZgQ+rdZnY/HGm79E3xj8YlF5jqwLVz9dVAhmPeC5WKlD
XAfyPisEK+Vl0Cr/b8l5bbN6Q8cmccdpHHNA0M1g4alXDyHED/yG+W3g+5hc7o4p
4i45VNvTy92l/44iYmqgrOoMwAEuDdjyc/4Iq5zIFe+1rVyDnn87btNYLPiIegFx
Fi6x4p4UUvE3arMUH75ULPr0yan7LoUVl/3vA4S/tETlMq798Td6LnsRoz4YJMHT
KUgIw1K6pXGt4YWwN1tKkI6ZYEs2h7TwgT3zSIhiA/NJwFmNietESTE7hOSUNp6w
1Z3jOukK6VebRVkCwtodotJDb/TDwYKeUEBJ7e/iNUbDCPQ9SL8rSdjlwCXLr1zJ
3w6+6SbM8TM4XY6w9dyfuA3idjwNYDyTMINxrn3NmHtOMqa3pBCgBVUYcbbuscq6
hou+rEJWc9h9NNsDG84wWWoJp0a39uvIgFmx2hvz9anUQs3BnIhyUj++usy2afNc
mtqBl4Pda8fjgLC/mgbWWhsr4DTUJTOIsKvKwKL07VPJVJ0VZRcpVoUexD3Jt8hx
idFHN3+0ktoryVsFEEfMPRSzNtNBspBqOZaixTCBvy1P97CWZZTu7XWELZ6FPS/K
pCcaYg8fDSDhE/dJs1E/qlolV8YSaSD16CTjcEryo0dbPH9/0L2pKsHoGDADL/D+
h0y88F2eD6B0oR9pIj+p/AyJUIfGp0hr4l3+5DLQJHlvH3DS9oitF+0NS3hPwnoK
lwiKU1wpSScMiZK1T9emnAiUN+U5Wz2iK/Xjg+2gVa1T8sS1cGZjnMHXy9Jcpjlb
0ROt+QOh/81QkpnPpwVNN4U89xi3cnblT8p7ZlbM6Zvwd1u8bw7bE3t1TC2TghCP
NMllOAhC8rsjsvuNGtkIy184LjeDsVqM7owSzlPGsjh/y+8Me8h9ZZLKeraCLeZE
ZaceVgZ+hBO2cUUrdkVvfqWAFKA0Xs+WyAs5Dh0Tj3rLOpBMz82JhPTLyysxy/EH
6vvcdFE1YrZ52ZmEEQy+g5QbwcFMybJ27ZRnR+iwZn3YxfdGLwKMmZCASz2hAnor
HXTBoR66JoMxzsxmMi0pPUJDm6aU332a/fBMNQccqQbgguMAHKvyu/cuYiGUgfKe
PUjH7yUSPpdGzW23PsfLNA7Nh7vfaRGhK6FfUS1rkJi0uRobxhjNC+ISBmaajDlr
fpcEVTXao/t8Ti6A6YzfyxEPy4rc2vtsWHgKFuvZFPLy7UNmZGJBCaIBTPAJoHni
bMibHS7yjxuSRROq2BFlIcDKqCaAmZihfpFqYwB45hgpXRXCzpOb6kcaV22MtoOE
THr7yPecInFLQIjopc5wUUXEIeNQUbZDNThS08VEbiWdYEWMEcxRus3dmuWFuLgr
p+pIGr+60pQOmqofp5cCXa61Y/OyRrYhGFLqwu4HE85e3Uo1KqTMYs1yZrRdh/Qk
7gGiMVP09KD/RbQcb0uYaSqv9NO6A71aqnJfs0U8LesxO4o9ArdUkqaLjwWMl1Qy
XJ29vxhaIyVatPMxoTpyL2grEksq/svPaMnAjl8TZILjeeV1tSYQHk7z7FDIhOGe
8HG9IS/X6XN886nOgOn5X1kAjO3MmXk6KjMw611Sea8RuWtcZoPyXNX6pqDo8ok7
h9LBMx8XJi7MmEE4TQqNt8p3CGdCAc3EfUfW1cQdu+MUH7tB9t9EiMOGR4yHWf/R
BkBNknY1hYr9DKrSuJ9A8SD3uiMDLRoG2juYIDrRyrPZVjQYYD7V9q6vm0lA1kzz
YEDiolLcC2Jiszm/2/Ub6eR9dfi8igeI/t8eo97GwS8LOh+2nAyDk4QXfkgmBt0e
FVgO8vhgajyz+zfmsY8NVAOmmQn8JxREtCzK1zHPcrrXZt3A6sCD+Bx3EXymlifZ
M//KtKEkOzG/wf1tFoXWRSKlFj9L3ROpjFiynrp3SY5TLMfp+CD1WTV0GnTMhq1W
5WFTCB8dA6n4hh5jU1+T0MW4wQDkgPqY4xuOa7c2kncNseQARvLxpuyaozFHpYPr
y317vkBKmcwMF/a3q/m2pEqVLLGPz5b7JOET6gSLaklXotOUUWDeWuIoNZq9561A
oZ39yg/bjCm8qwOYCBgbf+5/LsJNVUXN7MFRR32aFbLq+W9mtBKa7r2G/kMvhFzd
IqjhAWIFieFhczNFa+gO8SfLaLXqTg21q6VVKtGuHJRRjaATppoqpgGVRpeQgv41
a+EdGJCCzSY/W/j4KtvcL7tFNNL8aNVEdQSfzol2V7JfSs6gQayuhXUX08pPpfpu
8atwnxWmerqYD6J3nnOIGUwpuPgnTkgj9/DgNG1/iyGqn6+hCG+1jHGeNyI/4ZPG
3sxyVBc0jF13zmESpbrDMi7PnCZV6AQ+dAX+mam2OEnkrUiVlUa3td3FFDZ317FX
ZzosLocElPMQXu/gIr0wkHAf8a2cvutt9ZOD3LBPnxPKY1Vn9u+4MtwBRcLSM+pP
n6oTy4deKfTgJVc+l6tJpVWvsSHJ75a/+1rAnCLYOxmu4H/r8Ze24pY5g3W0s4LL
KdCdXsCpF8Ocnf5njBRbJfifZGPLMDNGL/sjWi4wSgirfBFVE0jn7HZi0gxv/iol
IK2dydYZLHePUWOzL5q66+QCiI0v0ZOPIP+CzYETFwvKpyRkvcjGcOcezzxNOtvd
cQVTG4RGoI4rEylmV8JRDddCuW8siOFpLLEvNM5eEWsP5PUIyxZutb3m6gFCnCXu
/YfRzPXbXMHoaDwvVkQIsJmLp20UrWzAJIl716hg2MXPPELQW4jghfiEmLsUgGzw
rabPNTAp/6lBp5JXBc7pqKFnXHI056VQ5kYOtM5uGEf+ok4Sg7coiQG8D6WJ8ZPn
qFYCdyZ615U80vY8dmJSKaREfGNZEC+qJLyp079GovZhVDuVZI+vstjrqm4Fr9NY
kmaXCF0EHxc+wx7FlUbiuR9HIX97Ni4At7jyjEIlS1LaRu0pC9/y7opS+153utBD
JCVsPE15utrkZ7GQwXngjjT1hUT6qutBVAY27TZIiJFTB07gT/92Y63NI81bWbOG
ymdzgU5tl4flkDnyg2vhcGNj2ZcggLDJrSuJZBygUzMmYPT1NMsV/Z1qd2bhJDuu
AlBWN1vro0sAQhynXVFcWtvWnKypgI0q1fWLnHx+vBz2Yh/AMMz0qqN6TGiwq/Ir
wYJs7AsGN9+/pK26ALN0zE73eRf07soMNQLmq93xgx3+3Xv+QjZupPb4/vmFQ64w
W6XOddQkXahRXVey0DDkqOK4VUTdSyw+R/MZdqUJUIr3agVyADHBCP+xRzkb0d7J
4OsNY7fWtwLV644K89UOLi7fRe1QG7bpFEsGjdu4IGcaTmN33kP9CPm0/gI5Nde4
5J8kKJYLCP44j9QBNxORwpM72qgXEk6QL+e9nPVCt6BpUecQ7gibrUr2L/KnG0y/
9HHuLIFO/4krqoi5piOvDZGTZVyVFzfF5vJo0n1Gzb3QrhVwkf2efk8oy0xaBiqu
xzFEhla8sohnaVwFW4DctlG1Yq4ptg8r71dLEwNger0iy4ZKBvlBDQPjByoxqkCh
Q2hOWWXNubmUCOzIvBpbPvEss5Pqv0HA/I/ha4L4G2kqmgIIKHX7M2FkdeSM/Lss
jIg8cfBcv6/iSX7rQzuTJeaoBn5Qk9XhYIrO2q6H9k2AxCz8oVBrxY1N/L7ahD+m
3w61FsjvZmhLLELFuKK2SLcyPPC3hOdizgjmXafW7Y3eFHnDbUizVaFZZ3s5pEES
BOj/N4MLOUxSbWw0336wNC2SHCrtBqvW4zGaZr4p1o82Z3vfJcWsTT+N8mFxpfud
3OlSC4YOJ7QspLb8+ziiuVwJ3dA5V1B0omuLqOS3Sbtn3anAhhg3OgOuBAGd9wIS
FHtDFf818yHSPDBGMdVidpiUoDii+BxVzd02sqlQlqXL0iSf48hWsZuYmLHhSIuU
xAO58oYr4NxaEbN0YXoU1B4VXe/GcnNYp6S+W2VeCW3g3EitYEnycq0nPlJuGfIx
9TDHir0jVp2qWKeKTSkyB2faYxKsBxNkotx6bB1MdyHDEO9S4woz4a7o2OKydTen
4nqjyysDHDhE5SXLLYUFpUJdO7npnJAfjamh9vx4PSfe6aA2hDZbtxE07AHEdEpx
Unm0sU4wwwsWM5ZWLt8xJBp3XLn/+q83uBUep19mmP1pJxngxsIqmt32SmGQqDk4
V74BchhTCNIi1QsLW0uXYp1wOpw4RNNhlhDLBx26BYTDJSosU/1hGc8Cy+NoDfC3
t9nEVXlMuIfVZOHbHeYeWph35XxjGVCIYJ59goo9tz0ji7XlFYNOcfyVj3JARuRS
/+bGghRTWfGZ72QQRRFBn43y5hQZbWJTeMDNW2hjRwWFL/8nfte2/nHnw1WsrCoV
xLXrve14hI4QGVtMD+AGkZ9PY+OpHhup0qbT9cXGhwIPU98uIpXvY3k+C3PHTM6Y
/SapTWFot91IFAMAhTmFHEM6FGJ0UA4uKGq/DUxSeO+CUCMYaJ2Kyr4A+N9ShVUO
+PHyCyiepfs4dv3iO6HNx4oDwsjvS2AqlRbNvj5b8kLBnZH907JlXDZZUYmVSQTU
rOapsfzmtwXzvM9F4ZJMqFcPNBTER+ltIl7Bpzp/R+cpye7cgBC6IblJG7vYc+oH
jtFJa1blJTlgDVSR2hFTBxS4wEC0xSobxn1RctTQmMf4+4XPwcJrcnE/7bDzT98q
8YIOolGgFHJG4IhLFbLwioM1YSK+NqMZSLaB+kGmwLK6UrJkrvA8BCogDGkISgtb
6DTWEr7FiGJa7qWWd7df0PDbDzn6YPoNgHw2aZcGaQDi0KRnUd27xFX1TI5hL3bF
h1QaWdqlCHT/Tsr7Y37+4tIGlwC83tE/F1EZXa66V0NXxwk0keaY7FnWqzR6ZHwL
gxG9Q0FS6sPwzUUy+GkLPDTLhs/CGgJFz3U9Z5uOe9JCsNYyCDxf9l6AOGCzvdJI
NDa6frG/0oMhYh2w47+p/bUAvHnrFtvlO2iws67wziH5PxuPE2IxfK+H02NErMbs
ea9mJAcQOqLIPKtVhX241JaZT2EJCBbdLzIi2RPS/YyzRrtmMIHv1ZHaovnhpV5i
0RgMl5xaIpUAKGqufsHAodf1U6qzKeS5vcQTP80YBShCK4qp+brbXPIzbP2b8L1d
qMpDS1ieVvggpoNt5jZdGRAaEsFhTwFFxiBggjcTL2xpWhM2hyiKzLefflFt2PLV
gyUrZfvdVLQ3eeLJnV9E+AEdc2dClGF3nlfHDqGxhsUlDCTIR+S7YQdaVhnBqPIq
g+4j25H1RftmmjB35Z56WniGsoMPDDz5FAFFyuuAOm/PxZRgzUdZZtMYDHYE0jRY
0B/iuswmgodiKzuPSkMeKpm34C99xZ8jyG/VdXGU1W5zzyT9ZUKNsaBjv4iB28iW
uJoB2xxh3U1bU5iSDw/8aVU58eWelxZSTC5N5zpeSBntdNxOHqZaMbvmHle5MAku
YB8WAIfQlJQuH/d1xYzMb4Y6/45peck+/15absXjCuoN6IUszDS0vbpTJd8v0l+C
nd68sh2I40Q+oGTr8oVHKPcN91mK2jdMGOIInQPf7UeEyt+8MEqLdKsd4dH9VmPV
WsyFXACwoQKk/guF5r09w1qkz4G33t/5R89ff11xj1Z2HuwOqcJ3VyZKLFLicFox
WTGCWubrdrZloO7GJrmAbYDPZJKTcyr9xJIgIFIzc9xi8vaGb9KTU3JroC1LrVv1
M9tWCgDjzf9lpIik5LXw1QVYRqhp2zdr3tT+ghV08J3Q9sMh8FUeAS8STiOaRfUd
Qj5Uhcu8AtN0eBHQMcbQQmhxEX81Nt+uikidZM+KIRGwr23ffuDMvQR7uaHfK2Pk
aY1PkC9m+kFFofycrwHi7qt3KHRJ+eHT4SOyDEB2QdyJRoHr0glpkLK8Ibqk0SOl
whSBCvPqHWmCrXANgDuEHUQ/q42ZX2bYKdu2QG7G3PqK17jc/H1xblaLwWkkq3Kp
Y/dc3ipSwA5004XUhgNVsAHUylFIMk1N1ZYVWONsUV+29sOQqieL4AsUMU2hjcfh
4aE3cvuUqjP/z4Ub6qPYmCK7E2jVISw003eOGwOX26mzVyuRRI7MBRqavv/6SX2V
1PD4CWyijxy9U5MUPgstpbFpsNiVZZ20KtfKcVn501v+tJOA76XdYUj315DXBN0k
cDngY+B5DY7ltylyR8q9OHt+kURIWJ12bun90YJ+NZmbaI9JOL9smgn3u7/EH8r/
BxL+QqtDsZUIr791y1DbuMVtVTViPlGSesoV/s70xPThYxuY2ZiKBtCiNyn/fJxJ
HRE6hySjKWBishr3r/HAbnLFXb6b3IL5kyK9v3yqIFGOaNwu5lTdzdihht4Er86d
5iZ8gL4UihzrgOucnSij1bL1IuZ2w0PfhNSDGfloiedROrJ4AniiRuBIIULzMPmF
s+NOGvnnYj2YcPm5k1eupbN95bRxGym27SDgMxgHO4mc1pVW9zjHhRSBfD12rEzD
XCdlVtBnXpHiOcbN1sA/UEKhVx3+qYwhcrLiKU461RtodGVd/YAAldK4eZ/mCWUX
/Uz2uQpw2xLB12fl+8Eh6CE/GeuPjsgeKwYjFoLpR/5Bm7mTlZnTY/2ZgyUOh+l+
SIEX3FoHLxnlEiM4K3X7ItKy/5VKi/VV9W5wTuLgCCg5JeckOdVGFr3KJU3flkzo
il9qGMluHdfaChrmVopnYbLTuyB2+WGk5rB2F8poY5LdBZSjUmBiHLmi18+QM2Mu
uOsPwyI0n7EhA+FEGADcqGBA5xsPHNnRyokXPIfHddj/BzpeA5MqvEsZPwCQ3XTK
j7HwczhlQZcc3PLtXzntp9/aUR9v+ZNexdWMq5YDwqWGD+IhFP1Ah8fGGmdgNwOT
mKeym2B8NF4oJxLZea+FLH51b5MzdiF1c2HuNNWg4AYAB6ouyKtN/feIIQ722AuE
HQ4FC7/mup1tJoo4eaHsunW+tophewdvroiavUrbwPOd+0sa7f1aGNeBHKynIVNH
8Ws7ykVUVjJBbRBKEvjptX2JVlwFYM8k05qDcUiglb7MtaNk+UuPEKnwu64d6FsX
wLzpyIxPr7Ke9mi2iRA++YUCV7NHTRgjIR/X5jWFRvS9bY16Pv0R6oWj24qphMco
rN+URDpuSqCfrKfx47wFGpTTuRjc1iNGF312tfAnOT8=
`protect END_PROTECTED
