`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUnfbRGTVGV4thwj05ePB+oC21aYvdxya2g7svB/AsEedIRB4Le/+03j0SnALdi2
rB/RHgj/51qMpE7UuLWDQCE5ZIWOaQk+2kei/Q+D23s6aQEOFR+IOdOma4o+pPuc
T0kRy/3ZvTGLC9cCH1QC3+O/oFZB55/ZttkUHqIWuwmjO26yDoW1Tc+thKeZZivo
DCvHZF5B0nwk0vXMnyOSTOfTB2OvofFAxR52n5wfxBKmTKAfp8ggGSVggfwbdunC
+f0H0rqNfGMRCKMuq2a1pSZw4aULW5HU4gsKjHYhYf4rucgMmEno05iFfNj4dpTG
Mzwm7UjcGqGssRJ0w8DDS7qkMluvPkI3CzoUPoxgasWcQYD7Vta9CjkpflKXNBeg
hUuM4VGCp2wwXTcu16PX1R3t4OWZ0PddeOFm1WiVXuxX7bpK1/d/8/oUgpZj4ttg
b2/UaiT9jQxenQeYqttzBPhJDXYgWQEMv2kVYwWiTvYZokuCwkrFhWXfTaAUCZYd
VOnGI1VUUCVDtYqRBgV1tKsYBnQhjUPoItIGG1yylDJ8Sdb9b2ZTb9e3ELZRvr1+
ixDmXhLCdw9aH5ny28XefrGYabnC45neBEml5wGoTldTVCbqags/P7Zpnb2H6dDh
fGOOSDvCo73l6yujHiIhcsyJrBL68n5TIlIioQXhhf4moV/aBL9kvj9RDy3llPKS
NCv5osKCHCk5swEKFCpdWofchR2qElBa54zV/vNWgxqhwJdS4D35vmQpLEywhgQS
svme6zNWVATxosnG0XEACg==
`protect END_PROTECTED
