`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQfae36bf8MtlGKhEqpHcqr7IXrofvkOb1643ldVMcvY58Ulp+aHTBas68rKE7y9
qsLdBv7aRTtYquL+U3jXZt/qjDEoSFfGtYYfhy0dn4Yt4r2UJ95o4ajPUN/wsvpA
7HlO3iWD6F89Uo8RJrvEWPDZOSBE7n3lNNuKSsX59ICwc8gxO5Zh4UZgeJbR35Tr
6c7G3X0m6HNMKWmy73+immFO9gFgukz4qv7z6pHL8oEIpg4aB/GL9mRB5p/QTw2a
4OaMNobZnWaXF0NqrMJDT1qEOoUmYcz0zXm6DLXx4+wmho+y0DEN6yQa7IWZfcpm
p+Qg0IVoOr6SQvUbeDpZbNPMksquRw1gpTuMIpIZm9gTF4hhsx9ex3l29GWbd8Ot
EBJnCGTNlaTztB3H3pgFHov3NQUW6tLEIS9x7osMA0Q+gOXAQ+7LwS8dbtqVhQC1
LzSFwyzFNcDx56w+HXaXdwAjkbIowGX9BHcK9iEL9ftCgMUv5jRfqtjpMLJRAvd7
1fi/5OSbKlCslq6W85WLip7zoocy70irHOVUpULAcNrLERuwV05gAfFYu8nrf9bm
CvBLgfmmCo57I+dqLSXAbw==
`protect END_PROTECTED
