`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NOBZwOqX9HWHpJeWXR4YtE86vhaUpLPmsibf10T72ywm9+DuSSGApv5nrj/ruCF
wYadFb2IIFkP8mPRNC0P6B3bzKw5q9CSethowBMHNOTavmn5Kn7WkPqCWTEE5RDD
51KewJFyKBOQ4Yh49+l/Dzta6ayuw9zdW2wUe3b5fBU1W9ScSPK4toNq48blf6nC
IWxrSXm0ZhhG1vt65AsIScxvDb4RqI/rlf0aVRCBtUHNPQyfPPTWXOqsbJ/rzom6
y1yLNzZjXsYQZ0wfaaqey3CnaXq+THmTyZAY49Txh7WEUzdo06Rs85AgMHBiSoaM
NNFFEbKVjrIvtwQxra9ejYEmr4roQAwiVyySJxKUGM7snMX5C5EHbWxNlDLECAbJ
`protect END_PROTECTED
