`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAFI/8o2fAu+foXK6ozy9+UV4Op1cqEmTO+oJXyYsWhVckSsl4uc8HMXXLNpHpO6
D6EQT3Q4bb2h7WqAtb7ztYHv5yCdC1HovnSfUsLCaO+fkq2CzqcL3WcsrHqjfU6j
E6zA6qWYioCVX4+9EIQ10C+Xcllend/Ruzfqw4pbjweVG1TGIUnm9y/s8AP53HIT
sEEgmywBxmEvEIhza1wToNoHHPiF5IjSxWMojoj7yxLyJrpddgo9XMZQnklNULJm
0tzVlXVIf4IkOkiLgzFT51EWf5fk1IKwq2vRLi+w+MOhsScf7seYQAgagvgxcJ3n
pjS08DDX1bt04gzenTC+I4htiM/yNHZ52CfKHJkKsBJvamTNMbMy8bTJHNF9e1lZ
y/58mY+KidUBEGxyoq0fG8SkqmnVPTjWUxW5x+2uPtGhR+I73HQHxdrpFkE06PFx
P5y0y96yjgWy/GzcURv4RmOZVeYoOe2rHrRohCnyM0GPz0Y9sTMLNA+pYmT/ChtU
IToU0AmoQpkLSJnZBIwD/qdmVv3GbkOF3HfnEG8VLk2wl/nbfsjE2csezRaHHJXX
Ut9EGNO0HQiiJdgzOEKuYhTJiyzAmH1lLmK8Pj40P5xvw2NYAemH0BON7A7gT7pz
YcTQv+cDeTboP2/mziUeCCZoh2S7oUqYHTxLn9uBmYoz37KtbJGxzXyYXoqI48xd
9cQnhkA/p/bvr89RMiwXzELiObE1KKsUqURXkwqhTQwPkc6jakaKo6wb95GIP1Fj
YUUta5E5OHEdnHxJQxNwAw==
`protect END_PROTECTED
