`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7t5TuVNdwf0z05WuaEiJGdXi+FPyjSCDVc1/TkxaZF8j4SbCet2CorQaLzBzdaIp
q1cnXKMzMEO3Qryj5aBwKLXWcpfF1TDq4Z2g4sWy0218xxBXfw5gBZu4kYgmzbaL
Y3vlIvd4GfTdnLbc08bfRcd+sgoa7rI82LuIcgYOVm/HsvKYbn5rvEymLU1yVCKG
Ocs4WtvBfLjw/m2dF3qf7J+QnE96GqtBDAJhzZPWAEmH0IMCs+5CfpTjUT3TbtmF
Wtm5fH0Xo9E5r4jLFVm90qBuwYIf7wCUTFs/ecxxGPexYlZiy6SYUS8Cm4hevW3l
ot4kcx2grSrhe6yjiYG55X8i3+XepDPoBME+4X9cjlpsFBiNIZ9cLGoLLwsyqeAC
z3bgMTDxV4JtZB8Mq9XaKLP64csWM0Zmykh1mW7BowIALp5BRxhUdLriQP+LN1hy
9UVfLd5nq2fUtUrHbgurzf6Dmf/jfwtOIbCitj8tpUeLqc1OMlNOZNmSnnzmnb0/
HRy7pm9uHGN1wAiWgAzOxtlgKTW924dihEo2BQP1WBqK35kUxPdVnGt0DfFXjdWR
CmCayKrltCazZcPKZ7IwdoQigmV6+6frqZDVvkidvpUjRey4Iu/gRqZKjjFpa+xH
z6AnZ7tbcTWdfICU8wY8tV2wla5qDfY7es+nVqAx7/aKRHmmz5X7hNRd1SeCzoz3
twRx32NeB/oLjYuPa/D3IDoBkTNXSA3tlsB+33p1jST+c2tlH19VqeQ3ZV0nh7Dm
Z9XpJQwmxi0PQYLW5kO7KmEjKabkvEd1hcLrS2xqCYhtrMnpApf4Ibb+V4yEw/TK
bN4Sw8qLJOOHzNKCymnG5qlUgtNdL2P4KV+Yy/pD4KoGqWeoKJDPx5zhYhc78Pah
yRjscLqOqZUU4IyqUoGDUP8dANt28aXMvp8ik/lOQbcE2gtYrzUcg2lYtvfGKBOe
4L0/c6lVTj2idiKdkK/D4Ljgt89Xk6/Z8hhCGfxi9dIoVzF2E8CQ9IBv5kYKmwie
aQCAYSYXZJTGrdHb8lJIoQOm/3C5zjLPq5AW5Lw9jH9W2aJXAdZ/H+fj4H95BAkz
Dlh1ek14L/pROm6ibLUuvifvGPl4VgvUVDBKPG47Rw8sQjInn6raeq1xZYNKECF4
N0ViCxT2CjHXBX/g/QpmOr+0rkGnStA1fFXPnY/wc/cngfbC+quLXygo+hKUFsqs
5wVxyjN314mYXI5+iv92jsKsqags1g2juGkwe86bIMbQHMKMAtYWgIHyBNmJQdld
5IYXCETMpOTcJT3Xc8IttvoEF7+FVoetoMsh3gLxFl9m30K5eJrkOrbYRVy1Wv3s
ccuvIHltUTuwwDr9XM2mEj7qJMjCPDE4qyGF7sjqG2XR5DwueIb3ova6hgrgMcvL
qlh3cVZcsryQ2wf5I9LW2krKVQqjZTNGef5HyxE+djrSm+X/DY548s9EBK8owHdB
8gIAYyxqQ7ISGEmxbzbvMtAm5A7N0pt1zBUIJxkxyk4FVvAjX+LMfRZzeknBLdsa
xwcNYvl6OoAxBJMlHdpdjajrV9cxbR0daxPh6OwN5y0WXA+PdNnLCGC8RUM4ET0S
AHzCqGCcTzrj0h1BsfD6h54e4dfMZ3FJANYZnpNtxEPBFdv3eUPvGhCLqnWU92cT
Gf62+cEnW/xoXNccgro5ST/Sv1fPAkBRrTTeS0MeHyLvfAd7o19wtbg4Sm79WEsa
DlK8HuldN8fL4bpB7NnKJCZNA/s32IoqVogA9izeLSgqTmghlk/+Ic7sE8DZxIbN
hXuWzWpn6bgJ0vV4trbx6mjILbXxaeAebsfghZAOI0wcZXwnJksRxNe0bnftNqck
BiQOVOEl8uCfLsIysViLQwqJPdDiYFg61/qIW36xgRCxFg54rvlwfnpBbzGgys1r
aqqWl7+98rWrIK4E81Rith7oipEgqv7z+rQ8x0iAdyRN5A46SX1vaOw5k1li7AGN
7bIoaeVvrp64qByaEMgKcRWtJuXZuoAXVi7a5mxmUW1K7gcZme7B+mFlUUJSQrQ1
2Tu8fIZIwgRdiWje5uT6IplwPZsGItDJA2O55TiQucUSkf0Y7GFo1nkO4eNveKvB
OuDA4AVlgCi/4o+riPPjy31Q1eW3NMUKnHSdcJUlXr7m3fiG1e/+SHKmyN5l60Lo
64fCBiYQvDBUVn37zdcAV3E1gAbTkwzWmXDPApyx44ueRGrGmdeT2af3/StuPUE5
velrI3EmRAW9mEQGTraa+cxwWgEeZdttA3wLZHYQ5ftT0EfBETC6k0DhZCKpU5pp
ziI9zgF40BhHRWkhNCO/6Keo8e19+Ik5tM2NUvcAI81XxXR2nSgcqGsNuC4K+fip
HLHi9iTBai2ojCi8ni8ORtd042h1c6Y7+bvqGcQYKroIMAZ+RTXtTCyv4wucZGkD
6B3LMY413MD2ey3/EAzt/HesmEVLCZXCbAclZ70WGsl8lX/1MvGC36NjnziLBNyp
jj10l4sVK/0ErRs9GjXlJType/0q4qxYeW7tBT+iY4laumxpDTtXEgwVsQIKz2TF
xfRZG9B3UZZ2ZrZWB+tSG3JpEdhVgNMLqjxulAE+5qixBo8U84R6uolb1/3AXL1j
opVnBAgh0po68gGHqIq0lE3pXVRJObFRqc0TqOvecxyLBi2sjNQjkr33pqqWiA6P
LDyvtTlwzQrmZALcmulxc2vtcq4aXXj+ToSPYjoJxzXstZQAJLj3EUQCypL8VL50
89/OM7UQW/7FUv9oiizoE5G9vZpJKw55MHMYEezrOz2AGF7n99BwwtkJYyqTzLA4
fgxOYYaT9AMlCAPjVfXZSe6QvUnHhdR2TSFPJv2OwTrhogjAub2y1iqh5EmCNJYJ
eC3eK2F1IkR0XWqfZFx8JoBBfiupJlzkiMBOmwuiVjkFI0lFIhNbKikGz2zFKz2Z
soCW5OTDAaaZwo/Pv2G55BuuITevqGp92tQ9zRqwVDXsqtmMz4qya54fN5IvGhwK
EGcRWmJsw3YJjjUW4GNcyQ6GmKRBeihBqTht5fCOTlnFhG9OF6/Ak1ZT+Rjar5KF
nEoJzPAqnw2HnIcMB/N10MDji748+tdjTtpjsiZlHKfJlgrIVT09C0yGpc198Fq0
T3vEoWLIOlZsvdwYr9ubpiWVwVGG4kTpWKdOl6jMwtmm/DK4gb7FiReYzQ7USD9/
etGc81+moEhJsUhdkKIeeFxopq85ye5peozjz4gSSn4uIPudoBvbJOMoy2kQ7oyQ
FLySdDwWyeBRNE/HldIPO9R2c/v+62wR4w8BzwgKwavciuq9chjPUAYDUj0hIt4f
feIBNKWIGWnpSqhD2PSXlJrn1FHb1sGHSiAoOlkEgaGQG6YgYsZPHbEb/BAk2OI6
dK81o3OsU5WkedO2LJ3K4Smi4zT12EcnjdapVAl6mSSSN5cbaXTOBWQ8ewYFWb4L
c/dq77j1cxokZbS6oNIrTEsiP9AE2Mum++jrN8ahMxeuKVdmgWnx+HtaESd3fgdI
PT3xK08k1uKeQyZhigcULi5hQ1R1ItHkxD6Iay9MqGYMbGxeywysB5vSyisaCI6v
k5m0yiOnk0qhgpxwcrk5LMtmyvvoY+XvlFUN3EE7q7Ux0ygqeMhxgj03b+PN8PpQ
2fYK26eGYNf0/Ge5csOkBsNhjiVGuaO9kneUxfRcoI1Ocj+6KCgc6IC+jJ1zMFhO
uo/ZXBccZ7G0PzBJ0uy7OvV135kek0s4HdwlhDrC1qjSfYMRFm19QZh3sO1WG1Ix
kiqAkASDCi9UaK/aX+8VKQeN3s2wdg6u7BvuTwYASd4oZaQYB40ZA7KdVdTww4DE
nMsGmdMdXiZwTp8lkP5aLUjjPamof2GIegWv9KVUeSCbwdZr39xRWi0djoMa1fRe
IwFT0uDbErQC3HEekTXh3Guk8XhF35Yxn5sr9FSuNJf1PONjRmIcAC3VwZlgHldc
VC1ZdWHpFnDvrk0nhP5yfK2n+3nJaqTqn+QtlsJ+A/By9gzTbUH/+NfXuzBNVOUo
Le9iPqhMY/82JurE4JIEko/IXLsmJjwIN3CIM4vxsdu1m2gQAaNIKZqenJQnDDPo
mWFm/9I692z0Th9UdF7nKQWwPCOpfDDQAi/PyUym69sSvRWIqyCLXy9PdMEGA1V1
GVj4g+GR2NTj1Wpqn1ro3QTxIrVJ9l6SpVqE0X+bB3eKag+ZULTYo7j0OjlGvYVT
8NizToCMvT9ZSBQHjVHDXI4zMlxwkCQKPEJV1+f3HVu7LL98UY6lUa9XeZyt8+Eu
vzVEsDDHiuABue9SGolANwK/czfmI/eXzHd6pSs1JfuAVefMjuu52Su1ZRygIBaL
QIv4hmDYEGvfRxC5Tzw5mEqjxQR4nZV4Owl4RaLQJvXy4EfPK99Da9SYH3G301CK
f2l2p4Z9V8B19y7NHBYEbLCa637iTsmO0vwY8C8igTfqTs38aWYV2EAn22Anhcz2
6X1SXQq88S5pQY5zX9HFDsT5DBEossyHfPqmxopOgjXvnubG1Kd8GyHnHuDzV3mL
NqV1PExacNtUgH3IgiTg/n0jMHhwopjkUkEAshMwlwBwcMIpMUio1yD0PjzwCxeE
zp0FuiuqREVmo5yhsSHvd66QVKLaZG9To+sxS+R/iAsqB0QF1Q12NTzzhyksamZt
Fuu/H33Q1s+4WGYBekdFaYRVG241CLxqV8mtYoUWT3QAX3pD0/8YFkRH6AmhAxl+
mBtIOrMspffkIjZaN5HXyywE4MaCLTfj2nlK5SQM/03S+sE2ph9QOvU+c2uZ0WdU
d6cncNhGa5B5OR6NVWsTazIienrUuXgko7w0/pMgPhZQtuDfEKhYpOUkwRpAiB3G
w3STgNI0eIeZYWQvpncGAaDn/qUN8OkX/0QSfCzeF4CiFOADXI9JaAG4k7cbY3Hx
KiYNpss8IvChfiGeve2bGv1EcrZgY1r+kWC01OGhL8nppDO786gj1qyNOjrwiWFi
xUZykSn58BzXAefoHv7WoCWXNWc1xd2+zo4Ih4hUhYM6ixBc5awlEGt4Iv6FgS+F
sGVJ0VzQO46E9tGPo7vyRUHmnElPkx+dl5U0QiC9IjGR7ct8d9gVWn1xluC3c9qV
daSC+nr7FEVyH3e0a/66xnT4+JdVPz2a2HYi8VDdcbI09eaVBilKup46XL4/XYPO
5w5S3VGYKZI6wkRsWl+o9JNUiZIGflCUUAks1AMm/rY5c/u5OtJJkyX7dvVB1wZS
45MahbaCFw2L6UhPlCTVitFQlOsofKlP8bw1yvwzBOVEMhzbZLWeySQXps6+zhDj
1KgGUD4TVsGtio1xyi/pNTGT7MFsaUJ+0tWNgfPVaR1vQpBnznLXvDDu01VDa6KZ
8ercZTGyHKDsRmrHfyoka2S/01EeS3CxY/I0Lx+YhJ4b1uJH9eLTHk+NUc9CoUAR
aXg94YjfpaV7Cv09HPGYkLjgd4PzegKtZHVZ57mvmZJhnnCwnAe7up7MdHd43h4G
qOqrcNay9FFOEM3ek7ZERlKAPoeau5zyCKJqLCK1iidZ7jqgbd4JbXJpimlwuiIo
AzqgwAAW7AAwbmAZ3Vspf20wmHlq0E+fBYbAJsFSmN80matp4XAi+fSFtXJWhe4a
o+3/SgYHD+cHLdNSSmqeroNcqcMBCdgv36L20+fHjfs003NNp9FZR2mUQBDuXPls
xrtH1i9OBatGVFT9z5YkiZLfc2yT9pZka1jkSuk7rzJnIVb4HSqvEIKnUOn3PGcj
NDLKFbmdNx4yCnJoK+Hav8Aam6m3tVWEKHQtij8siHYPMA4ukEhtqZY/w4YvE7+1
5xSeWVIxn6oEHXf4vKQr7CxwpatS0GreQ71O78N6eKzR1bk87sjLRw6UAfH36SWr
TlhGpRJY6rclKBV9TuNrMDp77tKRklJpxENuY/6GvImc4fLqs+aMN2DpmMU7HYkE
3CGHNggG0rJWJF9/VJVpSfTozQ68fBBsBddkANxWwgUiCYvt9VKJZEEAdrj5nGM6
DTuKgvTGE64ITV2fj7A3R0Cx4fgiHk//YZXjbJHMfZabptMilJyBZClQmihD5sPl
ssACStUXCveeinNvRzBqfOyksKwr8E1lxkBpaJS5HDUWDXDqYA4TR1651gNb7/jW
7SW15oPybFxrMZ14wSQEVJwYvxbnXgdfadAg1Nwgx74v+rnUxFki+C2ZrbZS0Z45
s8/bO/huViEy9RVJriMAloind64TzVFiqP5Ggk5YZVTjx2qU1X3wYpk693EY64yP
2x/s3cu5izyNLt7+koA6r6ErEpdTV3/WFkBSic05cEc+bFA50AhE6LSdEbWTUE2O
YWnlTN8nYTwDNWJVMni0+EsCx7JyVLwn4HK+ue5NPELLIY3PGJWu3g0m493rpawr
k0q/B5Yy03w1Bxg1nDgLae0DqQMXvCXi1jysmNEe81SrkBplZeGW6sAXXecwELUf
5VfuxXZGlpiVdjLaeFBSwPEwjF5FFELE5VNH3mJow/LD1BTrqlMmPORyYndqBE3+
EBcOH740yUmhD4ylFFxMOnm7fnY21V+X4NlvYjtiZyzYMCzpn6WnAZT9qyFzlSdz
HJ7ctEIxm41dee9ZB/xQNDQwgYaRo2BqSOacpmHlySx+ktr08LCZy8ozq/DgiBOp
zJDRPVJSGaeDC1yEdGWesHb//lArF4714KekXhIkU6UXxZFwcoeuvw40/J6ZZInI
H/NtR/M3uS0qwlhmFF6VndaRWKebJgKt5LardazQyS1216WuqboduLqBdiPtKqz5
I+P1nI15trkKwqHcClakwHsg7aGZedXou3+I3jZZenTgiL+O1wy+88+ma+hAfnKE
JKi/c/W12ByMSgzTz4NrLGO+8EPXeODBS4UP5fkFeOI/lDL9gVAizr0CUIgFXhnL
zw5OEEZrlVy3Hzor59tUjc6F9WCJSQjBOtPYjbi3nd+JrnmW191VIbvHSxuxfZxf
kxV360dGw7ITjkg+/hei5R7b4A9/f6jJBrPjkCWZcoHMAC//Md6HUSP9w7Uzv/2n
zi14+6phz+2c8k/hOQl46Zvx3+tUhQv0xVnH0djoe7xOdTt8d7ClU8LsIU3VNBLL
WPSRBOf6XY10a9/YU2dxSUsI9vGqufH0L/hBpdZhYQeKtqdBpxf5NKO7AHCbul4Y
oo5cok1JEKR0GmXfPk/PZ2jtWYLIwItrGumYb9wCtYklc05jls+mysOjzAj3+TkL
LcU5IPeU/KlKKJw3BCwnBVIancmRUezyKezNTIjIeBomLyQQAnqo8xp4nkIagjAA
skYUgR9158VW2XCz2ZeAyuf36OCjDtmb49+1neopAw6l4bdU0ags4jsmT9khNO39
Nb272oz9afcXUWr/sLo6XGni1DIXOS9WNbng61+4LPbJibgn3KyoTpg78B1c3pfr
GHj1JXKmRq8SjP5MN74oH1ncwCW+Zc3GYDooDhbfVIMYLJKRpLCXoTqIuwoEt/D7
I4ivxjFKcNfppYE+tHUs5MebG2QWd/PM9fwY4vg7yaBcY0ogSr0VexVr/Hp5sSIp
5PvqYtJLujYbk6L5pE1kJbpji7qM1HBQpt9tbfzbXxpJHp+0CApNlDyY0AEMLnvz
lzg5YvfoMA5jBdEuUXqFCMXCOLtC8sJ6mBt0P9l/2HpiyP2YdbPEk8bdXE57UMqC
cb6HEGfxdERMoGc88sdttXoDg0sszBLdK9btDVcKs0rRHJifwAdp7gkmY34waq7s
tFMEvaQwPD5tqisfX31dRS8GplnuDRTRybCUgKsLpgAAwEns952B18ZqrymD9u2B
vXN+S6R2mTF9QheIcPHLDzVizEWXoISccs7TARzH2YqS/xgUpsvtbifLGT1KfA1p
MQavFxILC2vx2b6NOrw7UMmUUo/fWZpsBrk3e1RIxeRW1vIqyKbSjLs+m70ZcyF0
TLmmTEbmmcl4vGXSSZCvnMDJj+PCgXFmvqRdJf2R2syjj9VXQzlS7flBE+XTM8Qb
jy+5yVH7KCwhZ54bIYb2sFNDncm1aSvRYYIpqKX7vJrIKYMOOF5PCievJSPCpE3R
GgXw/0/P3jQQLKomRVgvtEDk50iKfLBAtkHY/Ipfa4NwgmdlMgn8lYPCL8v7Dh0v
sAmQKBMZ+0wRA4vK3+n3ctQONn+OTLqSkTsRedQ7q87GkOF3P5UgUzBMWeds+IeV
OoWKOO7vZUEAqmQE4JyTp8Ygj57cyqjllCUQj6ZVOZPqtI2y5omgyEmaON1IyBC+
fWvtGC/lPgxX6mfo1qFAljHDwVUaeIMd8srXkZL5HQRJntyzqaZSAwymFkhEWvf3
BHz76O6Y3QFpkNPr1hJhP9XUIKBvn4s2I85ZAi5QFi3yMDKqW0svWzJuOK3DD1zv
3JT5eCk1fVHJd4vqMd8ebV+nYPodaZ+oag9276FiP80CXOXaxttva2MmtL1TDdnX
LAV4V7r/oCo5+eHeUTDqfPqhXhK+94AoK8GBKe64zY0sWGbDbYRCV7i/hlvbiPNl
0esQ8weYQiqoIZt5KeeI4y9ognleorjaBP1Bgvi8Qkk+XbVRo+iH2DkE4xboND7B
H2lEq83RriixZulUCbhjFWF2Uns5ylwx4WasyGSOfLFcFHz5oEOnNe+pUeZK/OPp
tLHq94dfvTuvMEgva1I4mb8yALiCjtCVGcJHwYDXCyQJ6RKX46sMupUv47vwLQhc
uOk4yst8QG/Fj105UetfrgzCUPG+06eZjqMrYTMiYmgP+0ACEgyhJkMKsf+2Z+5x
EuFEW1J/PAzOSCfNw1DWT0oMUQcBT73lA5nf98yQ7UHcevLXO/57Zi22biybGryA
QTQ1OFA6xHdI8Ohd+fQcpzNhzrOP8ED8dB9MDQIv3tB0Nug/PG753hPGHKIuPXDM
iFvqXiN0qChGJkQxTRy6XLpwQF4EVksqF7Hbr3XhaSRDCOJlQ3tOFy5MWv9qHGMS
ExOMvSgbO8niluB8mc6Qdo2UcvD0w+q2ArmUNSb1z9JtSMoJtLEhLWB6Abs3fZ9w
lPhwkyB82lq2YFgqAlLLcqx3vD5hVeFlsBtKT75rtiA/titAYkmtOmjLWsRU9yAi
OE9wRhBqUmfBmFJneiXlFEMUX/1pjgDa9nFTJ2itrNA5CMODGCy6tXHwauZAJ2oV
cOl2eaU3VBy0IDIKG322Hai6hRAZKZT3/ppEU5H1tMOSfE9mHHnIGTA+9X5/g7Xc
HQ63Tmv+tcKG7gOJtgB/D6CxsqJ9Ufirwmyk9Z2Nx+v+WBCpn+SxA24WRJ3LNANf
rCextP/O8i0HQos5/1lCwUUEtie44bSZcLk2yrAmvID0p+/qOnqXEvNOgXtfP0mz
IeOBdaxyDDPZLzzZnFMaDvaovrm1xbFkqI1hc1fmyKxsVKgvSkNRdrSWihfvgrei
zn9foMdajN4ZTsQCFK54u7IWNzPyDXHuDnO575ezdwUacg5hQyvJIdHLVw6D9MFq
CItisvxk6z9qARKzeR/m+Dr1uKOwtwfKQw4f2sztQ1QFxV+NjnCHEqndg58WLebF
10ssI1TkdwoTzlUIYmjbC229oVz7o+lRomGUsn+fXWkiIzGHiLPq+MsDpEp0zxd+
8ySTIyNMX564PCNMh51yIkAE2anCLF/LvT9HlAHKZMhhOSCUwwyBEc++YVLCmfR9
PNj6s/YrJvL8OCl7wgxFQulXDuYqpIvByah3koD4phdnMpetmcxthgFp8u+oZN6U
XRpvjJUYVefwUU/VLDveyyd0r1oQfenrlBPsK1IZ4Fdg4dAQf3v4xhbCqZsaK4WW
rMggD6uA7sALUjV6DbU0H6nhhud1pm7wT6XLEBRG1VeFVpLLysifFK3PwVQXxR9b
ywKK1Ns5VXoh42BjhmYO5ocGgHvWlVeohkwW5/anFIy/deYrSCIb1tMAyNEFQt+w
puh5uYcas3NDRMchjmti5DD3ef2N/ZEZ4Hd8Fibs0bfBodRqX2iUQujjUxOXQx3P
ENag+p9ZVwJO1Th2fGCCxZF3+TZtFIVRSl1wpZ16wuMHgE7crwV2iNQTlm1b8Z8Q
OpI+jNTcwXZ3b+GVOoR3ikqWpkFGmk10bdni9nYNPddhuJG5T3OLy1nWGQnC9B9w
4ELXrOnGvoTeecNqr1sJ1GKPwZShTrxYpGkHbAXX8hX/Hj/sFRyQPL1Ne13INu9V
o9c/AbEqbTV2bZe3MmyQnpdbQjzzlzAOOdFdH8mGmQ3QJ30xCCIYUpxxn8y9qxy9
C0ZpgzC0/WSM01jxRdqPGyQw9heqdD2QtSOjmXeFcOqyqsaZ6DlWzjuwmshjLi6l
gk+9r6wY3VnqcdkiSYUGXycr65ZRBaZ9oPbKuGP4BHfjkxSiAFqiI1T3SbWb0AHY
8TpyePpDMEjFBbu0TntGrEepEp8VtVbKCnQKRUd5HStenN5qsOqba2gCyJE3D4Ca
fJ+8KzNeZVkZkBPrgbx+8sozW3QMRh1CRrb10Df1GfTAtOpSG3VD5WcAOE9CWS7M
ToT+vobdDKn6gvVjkCfb6UP70S75ORmgbm8K1uiJjFUfSOEV3eF7cQKBWPbtOOo+
YcdRxFI1/+0afrS6h57bbXiYdSN4hMTFtHTDgChnfqVP4W1tx+cXC0iHS8XB98+h
mJhJE1GeW5Y08rmhkMw8youvtbcYepk9ZziJKuQvJqqO6Q5AHWRa3UCYNCiziVf7
vSh/C6NxEQoupmxLs1lPpIy550GLcDLsJbv8YQOLpCVrhphhOFzbiJmepDmAGGcT
wxJ55WMR8nRM2fwwinnGAjxpBXtliJyqfEPpzmDwoQBG4FvU7I2RqX7ATBfg+bH+
avV1vsWecuvh5XkQWVFNy1SZcZDWmF3HrzEXFRurx31I6sC/Iv/NyKXWPWL+1rQs
oUyKNRpkzp45wUhwtzcZxBbCLBBYKWYtOHTXqIXPIuKjoOH7Genyo4a4HdtpuVhg
UmHc9TcmWzFpmRAIiPQi6s55h2wkBZTjXSrVIy7sG43rKta7M7KIWOcBK33PcEj3
GJk1nc4UJ3AQVwygrNDimLw29YdszWLNVpJkZC8ok2Ma0+7uo8qyOXrfPg9L9rUN
sxob6uDGbnoK+cQPGKGNEVamBIcFrCLBD8bxp78QK6/fgeUnIrinVuoqzvBwSjam
c07NGkSPq9ZvMCcVfbuW2V5npjhuVNRjkNgQ8Oq49pbMK4ClS+9qykXf7kRWTh+R
EgF9VWH3DJREF8e0aeEfhltQEKRXgL6etWEIZmV0bXOnqCSS9gvmpg6jeLepc4PZ
fMxLBxvUZq62Zx4LFLIUYSRdZIyePtYFaSFByVwZB756esCQSt300HdWZhsFUSFF
IARO1UgVzuRkKn/OsmLsdPrzMEhBYWfGGXwqKK34sdLea0dPLwomsmHoSiQc1mBm
TjaWH5J0wgDIXOFgSEnmoJRyAQIsYSEsotvChMvP6L2j4Y6qXLUSQ6erxoHldzQj
oCjlzJHirA62DN9t9zpeS2vrxAYhlMdvenzsqev/N9SY6tLRVoJQcLJfCZjvwcFb
TPEWJp/HfGvoG9tBCSM9SaNp8gUtHHh8A6t9cLjIHDLAhvAfB/VnRXEVc+B0jmgV
cE2qa6NGkZbSxX6EhIESfTlWZMZB/kNdfXejQrqLFYIXX4aGhul33yAgH9KB9hf9
RxHHFijNa7IupbypQQjt9l9Kem/aUx7ZThCVqDGTCvR18CNmP2cp6ZvFQ71uPVBj
9LjViYAnbtqLASPSIwVuNVS7EGalOYUxxkcQSX2BMM6cEn1rxyy9VTJMd4QFl9FY
BRcGL7zPKYtaTVC8u1lKnwBpXdae8rDAkQotd3mWHNWHP8PkrHrXKHPFX0R8U5FO
K9aAm3+J4VHHZ/rxrO+SWFM3hLdPaBA0bbY1StTALiE4S1+mqfFnpj7PKGrjaASd
vIR7HXINeZyhwHqRQtE6mzChaiOswtWIkQ3hQj/2ZiCk8ksT2wi2yS56Hp4F4L63
XCbPD7OQR2TzQoLAJPwAGWV0bEYhGpVTQpv5GrrNqyP0mkNCrrPdXyTHi2HJSprE
CBcKUay7CW9FLQ/KvrIbKzMSCca0ExHlDEsWY1FoMaMvZFENFYCGJFH1XEsZJv3h
udhY0GODsdPumI4ZKWnMdkrkKwGd8NTxlqXh8RduPSjiMvBIA0mEU4JznoaUgrKC
/mjnwK2XrvbVIvY8l0/1obKTtCdM6ZyuTPFkn/MemcE275gPLMwvi4wItaJxhpCJ
Z1ld46/7T344wkkm8KYKlnaff+/H6DHaok+8R6gNTv0Q/aZ21QU9KWwJOnH9EoRb
71tunkxHblQmpwkgKNNMGIqtABquQ9z1wJAD61se8wZ9c2iyp4inFRvaxqyNzE2R
7ULvLwggp67vh5hpmCLUrE4pDQqvG7P0zcJknGUSB9VIXWtQfxUrTeqAJgSkjoYt
0Ir7SWmuYyiTTQmQQlQ54O3/JoXhVV2aiZLU3CNBAl013LIQ7qoi+iomU7cnwuFZ
bX3akzWDk2E6gJsMajOl1kQuqSeXxWVgmMZmdJgNfIDLV2qogZ/OKPMYKHIyt+EX
D7pV7R1g5n0dykDX4w8K3PR3MpmoJ8QNlnXcX36U+nG7HGcj9+OuTp77qVRst55c
I+bUUZmcay1k9jLuFzaKqg8XTtOGUm+Nz5c42l1MRGulD2vW8PMzK7kGjmhEl8Mi
qzo0B1dw91RUhG9Hx7wuhlHA5MDkVb9bo1Z8J1R3ed8qzSlZLPAildbByo+3hcgV
zsiRlUdJxM8vzAheOf7uRfIb8NcIy+G1jGNTfbYUgz50uJ9SM7pxK2eoeWedj5RD
scMT0VmdwntZzPOOYhvSL4Np7g9xHtm+BCcpX1rmdKjbxRdoG+QDCK1xKpeYVI4a
GBDT+Dr5fBTFldeqcob1A703C1pha8OBN4pHC3f0tE9DrDue3bKeUU7kgaeS0NWB
MPciJvtbaWZoFTbPY6PabUUlErjDIZC9F9JRxcDtMplixgoQXQUkH8ml80jtoDOR
9BcTHv2VwLPVkIUlJ8ymOM2p2IYO71Xa41DY2KpMKSga2wGoyt9tQW+Lr0f7SHbi
sLDtqhqzrKvghOeutMpuuoVPb43En5sTcbaJnNqf3jyqOyBkQzQ7Q9kHwcje+iHU
OAj8zNFVST+RTNySusVw/yfrNB3KO7DPjp4O/64ruvTMvsDzjfoXpvRQZDLbJLdh
TqfaoDKuXah6KG54WpYJvzmSTUBPBVijfwoLmUtIhDB9rEjupzs+WfqogjLYIVWs
lt51jHedW3YhqRY1F9P2anQuUWlkLPUZf8lFbBavKDANxUqF+LO61jv1mjU0HJpW
FogxgbqSSsb5kze+TovNfm6BkNiDRMnE+SK1hXf8Cyyoq+sQmvji+CCkOfbc2BWb
KKFqhdymAyr5o8McoPjaDHfjoYd526PdLqoc6ujrteIKNZp/N3GP6ingYnXyQ2zV
0n783FfFfeI/VZpHnmzMVOl+0AqhqNTDV6qgM8R0ygQ5/boh21dI7+vOTXm4FHl7
hARO8YNqherUYdyD/mUReDhT65WR1to/obOz4H+V/RTQKO1CCBrAzrwJunG+LCo1
k7zbf0sOfr/n06tLqMPIe5k7PcSaJ5KIL10rGO2E/I+to8R7xKVOIsgGvh8n1YoO
f6gV2XdoPhLZwJc4BkWeKMH8agrcRJZKGjYzdQTgvOvNfJMrffghqnX0Gb3689eg
nhw9LjoqW/bLHRKPU+jPpzwCU4LWQGbBfNjk4oitirHH0pTMYT09BmcZn52DDJPA
nbBy4Ze2zLvNIptYBGgpn24QjiAodzHmaCR7VeWS5qaV3T6VBJhxbcgLwhmuD+tv
vGedsOa705iLelM0XWfyZH8b2xeG0ldpsRXzBBNDmEqUmo6aOFHEP4dkNNvTB4dx
4+BTDA1Y4Tnmm0e3jYT15tyNShSKQhFiGHs86ERbbiz9DAU0oddVxtnQyLnznPa1
MfxYQ3NuTi6O17WZmWPaef/sExDDeC19te/LOLjncH+47bhjkxVTL5pvHAizsl4X
xNN01IGplRbsQRluxHbgX9GfSHj0gfYDtvyyKMTpYM0sN61KayaKOjEOyAJr6kja
W+Mv2diHXHYWv/Aw+Ob8XsAM/FpbhE3NFyUY/yy1AROrMfCcniyXijUE5r1Lbmp+
cnCFRTbEShp+mzD05Z73I6vUgK3FUM+FwqIKQD/ODcYZ94Dct7jtxhK/Ii04Ge+X
Y08QO9g0gCC4pPLP8xw5EtbgHZcPjVAHrBG5e5+II5n1JucJ65BsQDQyuFS/4bwQ
d2NuobC8WAQR3dJrPghs6u5AzqOx4jVbmolXzDD7aOcvwL5+B2MGDCkKty30bUIY
RzXiOK7iRKrPuUgeA2DAUkVjfe8qGtqbMypAh4JGEYIx3guZy0LO3H3SBkZJEm3j
b5/u6ho5iehofUQGkD8qQ4o1tVxrrer/8ZiqOkwfgsfL3agF3P67Pe/vmKwxsu8F
CrmqYCOU7fLG1EVT6QEOXc1AtDjx2OJJ3bOunQv02BD4wc9g7/h7g48mmZWkCffk
mQPQeVfFlyUg2SjtPoPwkle/CLXhXuSXiCGHIFKlQLS8g+YhWswG9k30Cn/g/S1m
M1lB6UFpj+qytaLUdoTjG/I0H84y6JSf7OBcbm9NhiaRAXTK+R9tRWq3Nq3rnkRU
XcRQowEMqraiA5+siKcRvpei3aHuLP/vlJQeUkHT2D+SPSn5AihNVBtqTIlcDkJ+
uwR8tI7zu/Ewz/D66lUeC2w0MwO3+8BcbVt8j4LBm1XfmOoX3vXU2dVayB/Qv2gJ
j5ZtZHsFBds2Mb/ipv8xYBupW6wFp8jm6MlgHhtkzID5Mw0zj8IjfuzGVcLSq0mv
FcYYhH5UhPHVASgaZU24FTlYtt0MhPpM+DZio/aE8hg102LaK0QbEuRleXcpoiZq
djIkTonFw37xrgEvY1YpaO/GbGQA+VOlNYyADojnqQW4AYmM3nZ72YnCjLw+3UUH
o5+7fIchPX+byfUMVW0WEkJYisqcpkixOTAJuy5sIrXW4XGououorKqe3LX+pQFA
5cYIEPJRtfvqWNlt5HVdUbpBltnIoYdWG7soIUvNPZENRm70EMjVx7xIjJNtJm6e
uuDtuq+LOveL4NmVIrQyaeruaAls6T2TD2+NXck/gtLXpFig9V+a2lZaouEYHvMl
0CZgwK0VORBP/Tk8MkEXwJL8aFslQr9zgleoyS4hCa3FGbbjzkyIoPrm0CAw1F1b
bhbcYSNiyVyaXiGm7oPhlKid81kdJlaTWkZcl/rk///2Ck0skfKYFPNGCkOAKFy5
9oRluZe0pezc1bTdTrHblM4W32CyHua2rZwRQUPxOzmMXjSCmlPq+K17xfAZXiPS
vzkTKbksyU3z0H6I+wUPYsmMUtdxhoK3laOEWNIZnRvE/0Pw2QglZE1mpSAPv+Y4
MoNdy4YWy75Rl/x6nTzCcUoyqQVwVYI69NXhjSN58/aN/7qTpbfUUdvu0Ym0W7So
UVfw+hypZWU1TcCZPNx0espv2QaZDZZCHJo93wk1+lDGw5hnPFlFEJXqfTAlG5b6
aOc+RAcGiJzb2IoONQuf0KGUZC0gQ5SGaC21D8g4xSkQq1fLgCzgrupLWMSfZ9MQ
mj9M/8v4l7ZOpCYKC9HnaJR2UBGus78rzZBWzm0EeIbWhPOeCSanpVxj3DdlxyH1
zOuTXmvfAI1pETS6w9OYjM+S6s/6BBSZkwnkirpzxV1TXyn0TfCxhA9lUn9m1Uug
+k81thQBaYnh7FT9SwRisPD2RJqIZaF23u9kLdVrpPF7KmHgXFDTbTSFDCpy6WpU
LH2WQBdZipXcIBFWpxfnbpS1hElPATIrZ772WGWMBrfNMuSgqIkGXbfP0zO/ZJee
5dTXzw5RvEHtTy3WbhhQNcsLLkKk6ndqc9JytFlSIxFdwMwPsjYwPlyXBiLeIrUX
s6J3xX7NnFF7piY4hV9XXvXYgC06lrUlNfhkyKF33ImsCrKmlyvuZrdCzB9Gyc5S
tpjn+aMqZjAy3XOrLkSB/5ooEejv8Ek/Rr/0yfzLcVmEkVfnABfby+DdUSgArSDb
fiD4AoW5o0gJhy1PcoShYlfd6hTjPpDdFQO1Rzc4GV+zxQKeUjhL2d3tuknPXuk6
SPJZ8eabI38BHb5N3JuFDSqSv261ahypE8kcWDSHy0zLxwtULxzovSWNlbXWTa8B
HYON/S2XDvxhd3qczNFvYzXPyG/uOgEITH1JSsgk8YzH7uloWToIN0UodPo3ttpN
h0+4TSxTcS39t5g7uIXqUj00Z1cxU3MuweDgCcmHB8cZZYlxwUeV2ynIJL6VIABe
DsETtfm0WDZI3VanW6BB3kyNm5PDzYE3bGgKtJk4gxj5bxWgc6Wx1XZ6FrK1IaA4
BdYZbCc8jz+Vb5lN1hFbO6TbgJB1E0VR621hw/pZu2UWkXy1fHkmWlYzDEmFSI0K
U2EWbKzcsVxEzKKkgmujyvscEZqPm2T1sGw/4pyBheo4bfV1fD5Ysw2peEHsVNef
Yd1IQkmnN9Gk3u64qRFII6TjoX6tamEwf4AXUKeh29MfTCvdcCgZ0aqpZCLqOHl4
pzbGhz/q81CyflY1ti1x8XCk2Xy05+ckOzPEF9wM5int0V6imcyzfUBkZSObUEYv
v5iTPIR2nza3qVZlOBkiMnI4Ycc+HgM5i4Kz6xCO319gp+aldh5LxgNGS3I/ie9C
TZeGW4CQHZ7h8/tRnHdK+CYePS27qu94kSowYP8mqFi5y/+I5U7IvtJztJyKkNsy
ERejh6b/bkhh8ZAzIwwN891LWRgqiRCHmobOFPSHkE5Wb10TzPyZz9s5rjJL1UtI
fQ4tO4eR5Vm7/6NmxgIOPBNW8x/8wn2JOnZkYyOMmm0stN+nLvwnr2v5pZ9JToBr
OnwbppVXvf0UaP+F2U4S1GUQkfoDWvMmdk2XwZtRQcb4+rS0Sqzk7rOttNQ6kV2H
fOVacvXpspEjcGRarsBVJ1yWQbbWLjG3c5B9oc8AdJW/UAEujGV0xZV5MxZP2gS6
vLRVLfCtz9TZrZmPaiVZ1+rqebzi8z8Fo6+o2M/p4FDA1xFZdJT554Zzi2ftaRh1
aZc9s46tkru6P68wxeFXXytE7mOxAHoLbY/pZfHFyX4eWzy3hsjWzw0WqUcEAVNZ
ZiHx5fOsm8x00Vz6sEgMuEpMTVd0p5GCU68QoOiGdOLU4ACuVneUyIC+PGmrRli0
pMswUTw0hGBmG1CngK3A/WAVM0muffsQU+RYDQzNu7ivgubivzw6n+oCnSfTRnoI
7wcjOIZGwETfcsfrp1Er6yYk+5wImy/M6SQjiEFin2DT0BhNXuOx0Fspv89Cy8Fd
XZIQKchVv+Sz4VNP1K6gsjs9TFd1Y8bEWLXo0DUvD41fUKPQLXDbmUPrPfaX9SJL
SwwGmHJFkE3IMLsTxR73db0D5jJNp4Nm7NI2HlSWCwrtP7cgDXAWTvq2s+5P1MXE
mqlWjtt8NPp2WfC2sIofBDe2zF5Kst8jw8teUy8lWiMJ7M4gj4d5Qn3HW3Y819T6
rOdNU5XbqR4EEvaB6SytcIPgZeQSEXF3SgJtw90rUj5Y/3jw+F7L2XuRhWJop2nm
6tJ9BI5DfqCOouNPrmT5aC3IpaehiXXFK76a/ffqJJ6YIRgdxnj+nkWrmU7WC//3
oZmhtCr2q36MakmPDxN+fw9Kr5InZIUJHPUAlR2BGt2IEQRylDdn5oX0tCDhiILw
7AEzizS1nPCPHrfOOlu01T/Zv5P8DDzh0j3FefGZE2RforTontJcyO7Uw5uHL5QT
L0mb4qagh8XEcyzxLDft9dFHP5iGqjz3K6Hwg4A/iYFcxZDhc7SvrXCERqEJRkWF
XJqc+7KaVnOFJLQE7KMztf2R4fzGtkrkRkbX+oqn8WMav0jYwuhu2J6ppefAiyoh
AK9spHgiCvH+o5yD91sbQu0hHusoFd/3ktfuvNN6MMiGs2L5omEHKY0sD5Nhpk+F
/iU1a/Hz49RF6BTwP1NXvlSmUPHh6IuBDoe318DG2juOHulaLrlKrJH0rDPc0JU+
ecCs5EwQ5uVL5mP6aUbwjAcVRxPA6M8rcfNCa7aKdadQO2olniaI4HfLYF2i3KSD
37UladJ2yQU7i7TLM+eFKFdiRawfCWhntGBI+VW84DYquokTh7UefJroOPIaXgcH
CjTVD6eiZsCcLyjK1P9s3hP9iuJMYKl/eBVx6vxOGbnfI/TFeQsVQDyvOnvvK90A
TCB8n2GvpS/TV10suwM8/YmuaP6ubuKxIFYkBJlk7VRbAU/t8c2tnuiTe1bMaoTm
8ZkJ6tNjFaTjunLtnNsrU/+dwgVNRziw6phAd5N1uK1VpZ0GUFw2IzaZZUOzfTK3
oMAWfpu3BjX+JpJHZBkxp+ad8a8KPym/SWxRu8YMXUP+1F5iATGofgjJrDpgdtpO
ScAx/iTxcfJnSHt/EIwSyhSh3/u6UX9rSZ6j+NpnZTr9DO+QLtrNgAuxCLcRchMK
gP3ObIhQmWpg8W2aAirgGULUlxWGju5wwnFYFyEXoCnvgje57GY7iA7Q52oM08uP
Vjq09+qDx/VJ35fBZsen0Wr9ijTIagpLavHoK+IqLEKZdhyo9E0jydeg51h/Gwi8
/0Fqo/Cxul8CWB2sz5opcf8FnbJdARXDDZj36e/C1HjfZc2XIIOzWZz+Ujeldf20
Z7xTtNXEL3mhtI3fMVjBrCpM4ER5fLFo2IvaoBivJ39AdsILYEfwJZK/8o/hBPnt
XZCv4J1yfaWy6Ie5Cf9psCM7AKVhAo3OAPeF2BtZ71d35T2noQow/BIu7h3bB4yz
arLaZzfjshDKthQlPY/dV6werdwqcIi2aG26tlkN79s6phBPwQIKd9fgoe8KOLAF
ocMejXIkYB3nB5aQ64Qh/4F3ma+NWUrLqFG3QjMu39RUzKCeiknn6Vgp3248fnD/
8wKsySzu1JooDKyFRTMUSVI+OhcOSw9zuhqRs9sxgjbYS7FsPiV9eFNCO5NOwpO5
Q6gK7ZTyc8pe8jt0nn5sIssML0JV1ockOcOVDCPHrxzEIRk/8Rmf1n+q9Ms4Rrgi
E4FWEsP6CFskMULapScLP9r261PSNnM9SawZTKacHeuAv6lTnTsxwq+rDqYXmAZF
lqhZYmu0lHbx0n5gAlJf67o6O/APLtnBe9G4+NqQ3PyZ58DZjZzOmLBh34WzKDWX
ZJWU3KcqcjMTsu/tz+yko2vOD8BAF93gqfLsE7Gyoklt/O25imH0uaBnzF/wjABt
jY0Pbx/Q0HwBVQQ3fADNFK4q+wjeSPOCG6tb7D4IDoF1InUKKXYPqYguqfwAZb9G
TZlUU1PU3SdJTG9c3OVBkMkIAdQJcKtfsC03LGgMoIRTXgPGRICLSDY7aJAl+jj9
50a6YOlzAjm6MvS9xZOHRR5JbiTSJQQot8VV8KP+Wyr3+iSFm/WF7sZTG8uzau70
aK3it+Xf8gs16zDz6PbPdvoNovk2zA6bgY8TWYRYR6FR00QJC9xiWmFkM2odVN0c
VMzagOhhfpoBK6a4W2X8BgxKKGdMLbibki5cfvQlhKelYqLWwqNFgnzxG0qqWQct
8qc6HfrOiz9FUDS8KPgsOS6uMY40I1+69SZWwwTeyDkBCJORASZ0Hx8wSFT/KnG+
1Tfm1l19cNibpFH3Rs6qsYL6Vr2sJEB86WXwi/EizWL3TxGkIRZTCqjae41TKeMd
WZoVUi/kyLiVK7+cKzaxQ4JNLMaQfD9BI3CS7Nd8SAwQm01iexb6KlJWidCvcfPg
C4LTJzRdEWTDDzLpEcsdsxYjZskEJomTs8eGz9KwEv93TDvP397Ex9/zYtpU5PNk
fSyL7e6MUG17Qy+2JZGERZbYWQsxyuiX/rvVe1ezKY43IenKFtZRoh5i762r3lcn
6wzqZZ8hIf+F9EhU/ei3qzdVON78MaxaJgFVUNaYx5YgJMFO9EUKM6eDnKtpetMF
ojl0954CeDRriGg/2B8l4YZt4f/zVvQ1xMng5BoJnksOSVIyRzxS+EJgQ7xPxuvj
rICB10Rcrezun4dsH2SuJAtftX5pW/TOziffY4ukd2+LkC9aw+Y+6i3eZlemnoqF
JW/CKWvDwjU2+J+KvGJAU8RbJTa57xn2jxGGULGF29EAuWvRfiHzapH3Npz1S16C
GbQ3EcvKHo1/mKuNlCbqLim83vJdNnkzMK6VVUnCpvCmEMLs14zPiF0Xt84TBbvK
GCl0W1OKWnH+a/7X2KOD4Tow5Z2hbax2o5dNwAomJdxUqpeZ0QG2aQfwFCtf7nX+
F+paXFBX+QWBS6kBrSz7Rb+GbGq/TXGRuKfl3CgnSxcrRYiDXVBLrUfs5QLECHKG
ctdsgNLm3Imr+udiSmJ4xm3+TH1/VlH8N7MruwiBZiYob0VUB/mcjpNCPmO3zgE9
V9v9dk70g7Y6hI30QutRCH2MJWkh862qosOlPZJBfaKJA01Z7bZgHYV4PjzuY1SY
AmwG1zgu2tT4z6YnJmAPJ+B/lGOKbDWkPHkrHfNHWXcIoIM5cdJKNwBHhAvZBbm0
dXBmq+F+LQkuVEp7S851V0osIkwzMsH6i4/qadUR/GrLSXZcd69ZiuQneDXueWBl
8t/aFgNWFZU9QcTCcGINez8yfrJRAPAtYuLV9exqxI+2ENFgpQXCIGUBixNo59TZ
WbgYyMPAwelcBATnAmBbTKGcbosVr7TG2ycUD19FS+YIIiD7Z9Vw/0+Q6a5aXVgQ
YD23SczZF4nLs/9I9PIDPGcGFiwgfNz/yJL9lPnvsThD0u17yeqV8I7HgLlNZwGi
NL2nvAaRzAtJNx/XlfGBmiBSWdcjJN6iXMDDvq1hgyrHc30zUU3x7Rkb+WimUa29
6CifJOOd1s5kzM/gXpSCeZbXSCiY2twBYz0mdEZhezDpG3TEQ+S3m0Af9UzTrvbF
y/2QzV5CyE8TDXlaiTny9N9627K9sxhdtDCWRkB4Aq2AWZ5agc5kYNGCtBhg9m/a
240WS+ABO3QnN4fB7baFd1CApXBzQVrs2GkLb5I6t0aBIOuZUiyxWbVk3sKZ8lpi
NAHHdS85eivO7tMh2biNHrAExUy3lKK2Wm+CrRMKbpy3vqkvSgjybISZza1AJXbx
ycCAoSVKDZNOkKHsiIdGUMpuqattuN3HotP5n5iKsahZ56VlvGGuDJ6LIMP3kwgr
2BO459OtJBIv8J9T+3f6mFH211qLqX2tHQWsJ5nIfeJbyH4CLGPWa74qzsDbR3Bu
8GmEgYdAHjw4pySOTOl3LXpOXsEidCTcIP07vn9GcaaGJdMPN/2Y71YDEfN/FkBa
qSN1LWx7cqp3tVNO7UUUo4fDpmaWBeBMh7Hv/RrgmTlPsxltuJ5vEdvtKg0DBmTy
fkw2igr9vMYqjKn56/hqejR/gGrXONG6PQKLSas1Lr1VfpujZfj5dxrkCHq5HT8I
UrKz1xHlvvO2xbSnUOCrV0nq9pr5hKnTOJwF+mvltqynmhiaFczKD9a1LzcTJR0+
HJxJfvkDfx0Kk7X2Aq50sWenzkJ3K+KvjPSPaBVUdYx2E44ZdaD15c2cospkAx/m
fYlz987wBEyU+hJaH8FEhB8d3UQvN0AuAr4rAMqU2bwws9VgSvG+fSdoLx3SrpyZ
k5L7QXSDyfRjE/xgmJZgBkjw5jYx9/RwtGgn2nmE3H+LxEE+ZD+3xjLTfD9yMOFk
FzNUBhdnysAP3Am2b9ygVHWWyfixlfjN2tw36du2dnwwCLO0EZoCurhNK8MtrXny
7Y+mVCBAlQ3Yuo0VU5YKMe0v1qi/Hs3S1AXVDqg+jECTZKkBWKL+UMt4JYhJ7OdJ
e5bwvwRgJoqs9XvNDcMLTW4SKEi+MHU0a4cr/LiUAIGZu7DCtgJFTAY5EchIjb40
m/1YLgtkGzV59G33D0GA45jhjkGYXXPM1vKJtS/U2UjaOzth4bibUS+RvR7jNdnm
fyKB+iTaDjcUo/hi6n38+GmhdPqEidilH6en3T1DEkYO+2zyQOJjRe+ANd+8FTWj
N1U7EPx1aL3rh7RfUqZfZb+L+Z8+MsLuLBPHg1x6qLo4A5eJpQJMTTccNAhWm9vA
Z3IASsBPyYq4gwQLHPawM1+viirPmeObAYahKt2yl4JqmFr7QbbGAXs+1uHYVpMW
5kxP1GT64DrsYX1ACD6BPdsgCi4p4hnt/QpwdeGDVP3au1Zqi76OGMCqiDq9HA2H
TLtet0g3ikg2hdEc9O1rX6ig1/ng4TAHVVPltG7zjnnZKqJPWwphdPtFEZZt1qfC
FecYRJpFz4613lb+cyzec9pPuQeZNX3AUg6VHkCpJMBwSW2r3FJQcVs4T8n+PajP
UsKFHgadxa9iznx7lKH5Ri/H4h9k1jK8XtGYjzLBhfoVPAwYjSG9V96jRqlpwqJj
agzYJejh3LVFZ7Mf37nKN8/Ckov0Ig3glHURFVOs1P+vbdr0X/Z1ryPrNZxQ8SlK
CER/WDwQt3LUGCTwnVsCfebUUKUHsFdeGseDBr9sn6ekgjB1nSVV7EgsVPbESeDX
+cUq52AliRMtX1M1m5Ph4KsYyuLr6sX/Pl7QjUe5YKjvIT5LHdOUr8RbUTLj1jnm
YUW3geuHkdi0Clyf6JSy71+PfaxRb88BuasGICh+Q6d14vpPvMOYdxh8aXyVuSgI
uVSAAHrAQuUh2RxGbRxn+Yo0dry3529Maz5QQroTqcLTi2I9tq/fiMT8JhT2LRx4
t2K9dQQJzhORUGdCU08Os3SwMJHeTkj1d78XW+sKwdCTx2gaXPmQG4uV2KUdA4N/
9QUge15wtwSNlj6SJLyyPpACFxT4XMCVuUWAOOCHNdin1Sg0fBI3SEVyGpn8ik0u
h6L5IDhTFQBTkohovIUSzkLKRwffcftoarWPCkgvUth/VHsmjEYzMLPSBF8oeoBZ
crVIz5X+TydV4JArERxQG+vZGjcVvL/7xBd5ul+izM970ttMjhu3yTV/OjaVwF4O
WmsyXaWxocReFe0rpuoWq8ysBAtazkcb/hECiFAVvk+ZtkNOq2QM5Y5zfX+N5mXK
aYL2RzwviqQmmc72ImduFbu7MgB3o58+Z0e5F/BH4Ch9vKpgucOcZlLIQOx6slYQ
uHIaYckuevXYSiRJt287i/DL3asE7RR2shTzyR1bou89tFjPSteitIIQt8Ka0/uu
mdktQDG74bUPFKqpQFfChy/cLS/ou+EAZXeWFKVcdQT9kxxiQw202ESvAPOnSm5O
z1VMp+BygpYtXsajZTrOmZCj2oS1OsVr3vfG1mCc/QAsTt5AnhqzXO5wngEHYljy
caP/PIx0XaB+T0SXamOdGqDvHlpolJsUleIPxv52ioO8ul4Du+EorYCS3TyOoHFx
71MkDnWGzAzMyMKvR+b06mVBVoM2d7fDuyJUbL40TDfND2JqBY8JOrV87CJirVTK
jBQrNBTp2TqE2q5ZkAp3SGQcxlILyvwX+TqpNgrdqe9MovsCAimKsWngJZggqKYd
eZztMU6GMZYMlBZYrVq8wuvlGyUkQDcfDotgo+d1YMlwCq7GyaaHBN8ZCplqTYpR
kUkPDb+LlsP4go+lIi8/V0JU2kE54PPc/v+Tp7yk0YoklSFL0MQk7PtsBx0a2mnq
GaH31uN7TUB9/8J4I+TyOy8kueT0rVfTpkfTdFrZUaMqRdxHnE54TNUXmJqSdKG5
75ErXOu3WDun511dqRKOUmiA6YWLLijeulfCRm/V4tAq0ixzm4p6WrGkH1qbbki3
GjrO0iiSp49bhH2P9UC+nYm6h6Dr7/0PtyHDm3tDaDNPcu80fD39gey5uxTzYzbg
sNdaGhDvhY3t6zc7ZBhJ9rmHIJRIzdVCiM8umAZzwVe7+KSoBgVESRwtKdxMyAFE
idIT1EoEOR3TQ9notrcKKJFocWrRBi6mJywjmWucRTWpF4XZXitLz/OUbTrz4dSg
ejrUs/6DHe/iugkj4WXulo6/dWUkntcIfE/OZm5kF10mbCHBH8B+WRr4Iexu6E7j
lRVARHMxYpPlI+Z/1ncx0nVUIsbwO+OR/2PrNvMjoIOaYZnekKilkL1jpU6wbyZs
bOeTtFMrrhYaMKBBbXFJTmfPZMF2tFNXUzcORBIUn8vETkh5a+ilqCK9aQUcttWd
9FwjjMT5oQcwcgwAfNgOfgrdEiVaDqtTz3hxiNhVVTfr8+121VXydKDw9hQB4/d6
/3oUkPiFgMFvxgunzzxUwG02A9KfAAz06RwHUJMmZ4rszasKSPvCZ7XRFex44QVn
k+KaVHKkHwQgcAbq7cgNTEac4F7szdk+cZUPXYM8d0BZXF0q+6vaHFtG0kpRK51B
3GH9OriT8R8eP+42xtZgfYUehONHzS+Is+o7JoRO3iMfQ2ZK8uhyJFjRpOona/0c
EQcJqfnOZyJN49knXW693jJNewWJFa+eYYObpdArJLiZWT32NNsP7B5uILBEGrlN
fChx6eQo/QEihFPS6xjFuCYefHL+U1jF8WiYnxcxjJHtYBcEcl9unnwn4vSSdKNu
HY/wCwYKXm2RU73TUoNQEaxVG0/PmHcoO78Y7N6uyWxdY1u+JXSsE+giWG9/K/Cf
Tj6PUjvCN2gL3/SCvxeX383EqY8/jjW7gfySYbI5Jw1T3129IEFxa8OHgGQJOQ6O
GtkeLqCx3od5u11i05docbu/Eam5BP3CWOK+R9vHZ+ap5gvJi2OS8oNOJoTVxfeJ
6s5HTjidab0Qa/DUrRInX4lRC+RsnXEgb81pYgrQLe4unZbfrQiJE4krgkM8M/WE
7gPkNA3HxI1Jnk69eFgdyKz6CmkOJNFuM2gfT+VJpKqhsKMEVXNoleP987rA3MmE
5h87LQrcklg1HaK7IsF76rSKJju0UQ27GSNbb7ae4yul8+E1Y5ELus0kjbrUCjkS
znWJePCmc4TLhSxrnMubAvA47R0W8hbzfysMWj54PYfbdvw/6Zr/BpS7LbaLJ5d+
wyEAhxCZiV8B1r5zbC9TLHtsgTxuiAYV67uf7vbPRHO7tglnch/FaKQNcsanRToN
spAWomWQmvVKF2YWWkNUoxDgt8rWvTKlQJrsFZSgvGX7di9A5YvCymdGbEFFaeFS
IZDFnvmZubdFDzj9shsREZbm6dbzhlpFqVcLLfhEaZCX2pK66J+NWLdBheHrH94A
p3F+CDOjO+p4T79RT4bka84TSua0ctM1AtKXoXu7x1P9S3nqG21ccV0sr3r5h9go
QvXUdCagp7OXV0oIoN1Lu/0I15KXGmsrHoNrx9X3LEceEPkPi6Sou2c0jWT4Keuq
Ev/aoSoPFmW9HTA/28xF5keg7L6NgdQ9Cej01VZFaEaM4wTIPbxtiK1j3k5vfZF6
9ccQsKE9FFriZUYDaOslzli+t1O9rXy9OzawQMx2H0A3inVDXB21k8CaoO8Ed9Qz
8V1Z0HMVtFTQjd5arIveBkeFJzRyUsLecAVleZQcOWuEpD6yH+a79z8VAgMzyn/S
/k7cTJF/pezHXAPaOYryiodqqY61EWPxKZ4p6O7XauENyjtBd9STgwR0xsaZXTrI
AO/QetNxEcnNHr2RnPLgBwNRyn3T7O3GuaFNPtQVQ8m6Ggs5CwT9xozRLw66Rf6q
2Qg05wwgNCilwZu5nXOFt9HmihcTSi4RT+xMbXnTYBWBqJRgdtVdT+BqGIm6OQgH
bpPEmiu7lXdLJ5xuPaOuL/O6/GrVA6M5/l2i1C5bS+1iFwmqJMOcBzekkqMI7xiX
7VqHZ6BymBIKuF42bVdT+cKVq0ah1LhuONMDtnqRIA+F8TQAC/GwR0ftvfSyG3TD
AtLHxlNNNaxqw6Zf5OisGR5KegYQ7UN/ZPnFazv/mnuh9ajib4lHCrBgXPuyRp4D
bcrS3EvFLhRrpdsA/oACPt78mREC+Y3ukk4TK4HddbOqgRahpoH0c6ggdGx1PuGz
NY1tjQbqRBzEy5w0fECP8umrGwfbmrFwykLQaZ8/k3T/20opIXd9xjQFZhXezA85
6BRjlvSX4t/gv0rGqxCxQkFJoSYXhaxpvj5x2+dxbpkcVsarRSr7gnxtw4Lar5be
ZlUId+NI20ilLFaVtawWkbafzTuM4ZEKCrwyFEweK/9cOpRqgbNHBu2NpbwRX19f
6CXCJSexf6azd50e8LP8zS79HCzESUFF14V5lhPBK0gc0KGDOCpFNm36bAdLlQil
Z5ruUCP0JO8ujiAHiuL0h8yPgMso9HE5b+7mWl6LdRvw685JWGBDiTO6x1fK7Dc9
mQHKTQcOHH2VsVBzg3ourcMerH8nUohYlJdv3eFvEMaw/bCpmJfYxBgGMilcIQme
ha5Zf62XMVZRUZAPAm5JIYxkNaO1urHlpjNEZ+Yw09TKMzU7VtYIboS7hCYFVhUp
zu2y7bspjMFNiPcL8Lk/Ixyj8A6IBtb9sWSFEfJj3U+SlkfvyAXktfanypumrQM2
wDvxA5xl+/ayB3r14WzYl699Mf77GZeu6UCLnOUCM6ljYnAGtMF+/rVAd0aU3d3S
K14aIeOLWsikIrKSGKA3TKpxeXjNf6tPX0B68df9irK+xHOAHAdPdy2MautHgyug
Z8Nv8qFGhNBYebAqztX/wMSup3yNeaXcUq1ft199rNGcoqA9sNS1o9KMZDQNGCIk
vn0EKKeA8XL2u2oSeHKBD3lH6JOcJ+x1vCqbY8cX14w/7UGvTVPOZsNbzHNeD2xM
vCTRajKveClSpiFn+XRhlrqyqgAcM6BQnmo5q3sS7vy0ErwSdbqcOJ6VyNPZ1OEK
vH0HXMvw86NuZ4ihGeX3vvUPLoYFUZnEZF5beqHda1wJ9qFtICPo9azS089qlpDm
oBP6KtIX1W7kJWoA0lrB8ohIL8pMNvrplFc1PZvP30nC8fYRgXnju0+BbI+/vrai
0DmeprRtnvPx5Nd5R/6S9yAPeLmjfBpr0hm4AiCCfz0LWcht0jCxk+3zjRyxGwZc
+6KmEPxI2o+TslsIyYnEDmpDUzp4cGvaX74CfTRJRIeW7YH4wXotZz1Rv4Kd3WPZ
O8S9TyOMXtj2M9zG9nqb1hTeqUmpR+M8bwuoNDp6GJJYC32lOTPso7A257fGZNpt
Qr37t2sDZD9dnDpRqoXg5+iFbd93MDVLgiM2wGt1y6+BhKcAHOQVwb4knaOE5/K4
GawQVRpoD9WpZUxs3i1ptWsY4gl+/u5MiJgUKd3WkQB4JSa8fDZMADBpoEKJR6kX
j5n9ZIyI/SCvNkpBYSZbJszO3++m+ZQnOnrts541kCANDC+4LQ9y5cpHQybZjsa0
z3fUq71UdmFexBsEkeGO1vvddAAxPY7eg/RZGR89WzQRMhliVajF6G3mFxBG379n
grvcaopbd2gi9zJhRD+vDu+mPH6KDzESMkVTwmZ5sHhfGmT9XrU6Ltc2vJKTLz07
FcC+8r01PaXlQcdf4LNEkZvmtWBjEduzDImOj6TYc4OdorKRt0guDW5sHj5X0TDJ
hAFAMy4wgn4ZEAcJ8fA7RAXb0TPZQsQ7+m/tZXufy3XX+FCiRWhtJx9tBd9ILtW9
8tyNrVUFhHrxkWf0aSvr2xJ0A1PGW0ToOCOUCr+XFiUjc5OvpCygNCWtnmbEaNhM
JilyvbYxclYrT9X6t++xEvbcKnHXC+5IcX4oXBzTQxHRXh4nfHiOtNETAab5e29v
hWr72f3BjmU8xfBBJJRlb4kOeNAVkuqqCcLEFe1hDli+PXvEL3QgP2hgqProG/Jv
7ZTfHRKRwb1w9dhW0QCn+uUCcmaMe74qu+4BHN137RXh8WvgPR/MWJKvnr3Tzxas
YgXqYNasQqid6bhQeaWK5p85jJiA2Z4wRnnlDjLKGiXdvgC/hx2XFd7tdNl10zZv
6JiTiJbz6CXbkNHMLeGX6X/bjf1uYJjJ55EHXtAoYl/IBHqoU3e/Ol6d9XQMWkNx
ux3BhnL5XRf/RV4ZTcHC+jHWL02KnBEn8VgrE0PcB52OAiNqcEdhKVYW38NnsQjk
4k7YZQqC902IXsNfMc6qWBUTc5/RgDwqOxRFxwbT1MDKoLuFg/QiscoNqk4VG4WM
+Hx3agAmixAjk6I/ww897QVvVHJRZkGMyta3Ahnj5uMIKZ+/HdT1ZQWupMV8t8xm
8daEUzBMEtQaBy7WDKQCf27FNQUhTxXj7/1sA7iu349LzCOSlc68MuzZAPPRnsLF
VpWvzwpUOMXdtd+ayjLbr+b/SdXUMgdig2l2VzNVcg0n70GhsUKUE5gVCbBdNvLv
C/Gls5NUDU6SqREwRAyO4plt293TKz2oEyqJney/fKRJCUgWrzYRrzSSQYpZ0Ir9
8QdyMSrEP12a+9tR/haKKuBqTjY6iuMf2d1PygOQdwpmGGPzN5ZyMEF3D8KK6lkF
MedvM4BuOfLz5HhEfEFoAbGApNFcGQA9aiSwx484AfXeUs6Zo62Z5CrC5tlVCZjA
0CPtviI7emQfKzbztYrb0h1XTSGb68LML5GwA5ttSSq0VWgoTxyJ88SQowkU2OcE
AzAYqHjpx74DllYbo3D2RL6k1os6maRNZXsQkAazegC0jOw5Y/cVZUrotYy+XXYR
niwk8XHYa7znvV0maNULvMOxRA36oqV0N2WpBf860j9IucBegyq/2ulZq1ovk3b/
9aQrFMz5LfRdfFvf06ZUQP0epf4uURedzNjDhM9W7k4SKJoEKTKCyNdmWxEkdgNp
LQzxgvHKjaZSmcjLolmosIHgTWa36480NPm+jOtQK4yvw49z9lyLrIW5whsPcxq4
nvOkqR4N1wmral1qcK4ANwfzgz16rV8tidD3XU3QQKF08dyzr9rygsIF6P3WEsi6
w5z6/tjmL2ikierM+QLrrAxynZzS36pzK0W64wEsP+Ri76VjjNR5AA1X38Q0Nlr+
iyrdC18R0NukpWZps9H3WtxPp56bI9JxEyoyZEgBQ+DQCS9KAio/wnPAu+XNeCo3
fnpQl/ZHPgH/HzqpCprqQP3nzU1j8CadPDFB0IUQ4Mht4/CK8+nE29XKK28TrTPu
ELSTJX6HfJKm62xW8KHAFZSBZYZQQY7D5cMQArV/Hb86Q9UFjf/RGHSuXy/bp6eA
VzCPlJGljF6bCqRg3GEpjNSt/Oh9zK5njvJL0spbcV2IvI3vwjA4AW+P1QfW+uZf
x/oo8BrHau9qEtI2aoHmu51CO1ILk/1FdnZ904lbzA7Y3hIz/axKictlSHLVQFRS
volgAlJYYBnjoKZSTK1V3WggUDa0Kkjb0Gki+hKzWWdRFAjWv8DR2vvhyyYk3Kpl
SUuvTUeQbmtrq0aGBQmNh6uEvlWfkuIBPCWZC/yNkU5YTb7TweALiEAjG2wp8y1N
K2vqL3maTnVeUU1CtvUOZjf89re2e+hVlyUhn9khsos6XwRyORuEZnEGkWQhcYFr
ntvuvQuQtWLMk9snWyr1ti8AlcHLI2HsUfSndg3Q4vW4urM3z70kpNEDEkYGo8aB
rTbec2IM78gC11xb2rp+VvbkGEjgEZi6UpQCtmqWhkwuImNPMzjibqCP7dMpCNpg
cOWJhDDmrprCLer4iOmDoe2Ru0PjWI6+nP2SK7wYcNn5rrpdC3f6zGuVF3Ng8NAD
WFJHoi1VHjz3Wr2KSdlFKYV+JXMqMKSFhLPfZW8D8nZQRS2cDBZgOoYtyeT943QN
iOHfPl1fJtMwzNchcM4NEHa0xLP0QQd+k1xisGVm7HWuz181QDdk4rVKrGSHwT2k
W5TQWZCF/4/Fm5cvAEJ+z0LQnhwG8KCRBZeFWIJvK1r5Toc+rZo9EHimwaYYNuwG
2J6ENz70rAz8J4ervFUNRONr1m5KnfXMiuKpIXUvO73n0pxtRHNICWC7ENCHJCS/
1WkiM5EPzELC21Wb8bonCF92sQISHikwuoWUqhBMTi1EOSlRFjgbsCa6hxfPM1FY
ltUgZZtgvNH3CUMh3BFC36aafvuTgUGx6rTviIVAX8FqWOvxa3r/c6FpWSjKh5Pb
9DNc0R/tRxhSMiVEnzvAu3JY0aEbZUcHIMqjl0lLQp6Ibvx9hIf0eDyPcf9Gn82B
1MGIQWrkE6H25i9W6t40r79Li9eINqPGWeN7Qby2X40XJVMfHl1rJ4aRjx/L9Hgr
7EP8RI77NXBzsSaG3uNyQOkos51pskJoqeIlAcfpfAvYgOPTrGPgUo2KRiRw2HdO
jRclsGADmdJRA9xqlcbNLHbn/R7aACwEMtJJC4X320oRFxPC8G75uyrzU16eTzgZ
t6crgvOKg5MRZqsfg9eK4jlTTFDqfx8mpIgugb7V7tH8/nYNx49I2yV7KDr9yI8Z
ORtgxA8gfDoGhx5h29jm4NfbRj/0yceY4CgO79Uehv/TKnYGgyL+uZdP0G9+hcFz
aI8cTVV5m5mvtxSxcBZRu/u1Fc7wupK1anYSJmOhb/kg6J8DAIZsevUMfuwaquEP
Z+WZaHLek8c7YICA+Wq0tnyApRGiR61+2pE/hMvKP2Y2endgNOthllbRvZJGQfQH
Ee8wJ3uXG9qW+twUXFL98SHzVWn+Kn5fv+5mttW3WqUsEr4WBGAyIBY2DY9WlC/P
0WfCj0XxwWIxtMbd5qmkFDkiw3Re0ZvYRduXlelcPezacEdLX2q+LwOE1zjWgNoK
m6VITEfP7JxZVofYxAPrCnWECvPLCzsit3tnUdkmeGBDoJZfZDrD8a64Azg22bI2
XHeBJadjkzz5A1+lteCNeu4dF4UiJMaonsm/7AHwRd5VHU1ebPZe2AxbNY5PJ+mm
2q5R5tHdvALeuUtubVOZOOaj2i2AiI5k+cxpfq0GT/tT6uyLTsIdjVghPjEWVhrz
1ddY+q2oNBAvemAv20XbrUvo8h1SnRREjNKzpyxxZKElR5rb8DTQfHoQYne1zim1
SVMR02veb9meGeAuY9DdJKGGqv0jSVKt7Mp5DKbHKoDXCPjUde/DQJ24Biu9pytg
WtMeZPrdh/fQ0XjD/ZGbb0trms6vc53JM0G1tK1IsciQWLWTQ/ewtO82tzxGEuo+
Mu+LwduVx3IMkwFI8lye8+RPWbZWzIqCPoDJbJwt28MUzD+Ui29OHIotxk/C9fs/
U5oGYN6EZibrbtd65fGwlj4EHclTGRuwDO9CqanjowQYStA7pqlFJGEWff3B1wtf
XmFRv5El53PrWd0TOC9bh6yj354T6w9e1xW3wByMDIMQMbCbeYdlbgDiQg5iyRMe
Ibj1zIE9CWfKOblOoe/cdeiUfyeOUCR5r5pIBou0tkWldS7Zjzq1QFZ6TcYhHrrR
H3tW0VdVkddzAew5S6BWZNB+jd32SbfrmhpOUCFMxC22x1kndRF0H4dVS5uQVsCg
8PahZ2NO19ypxvDXzSxYRTw4KIrHJPv1XxBT93xCNdxuH8iQIt1OLQFGs4KK3dlA
5uKXM9FCid34Pte+lFeR2VerFolRzJFA1M7ddUnSEix/KQ+Nsjd9ZFTh+us+ww46
CXencDiNXdhOUCFv4kBI7w/aN0f9P1YAsfowkFEoz5ce92cZsaEgEnOAnOpiUu2U
86GtU6PCTniQRIpl0DZSCu73E1eOAGVrVgi3MCpjAhogCKPKaOjXs6tm+eVwXvxd
D3c08H5KuXLcvDg6FNlaPamQcyoFnKSOhJ4jE86vVWIhX8usV77rcqjZ5kM085Tx
rEZrEqB4MiFHPXCq7CveB47lZ1L+zihRvfBpjAh+e3ybNvkWHpDhoLeXF4LJMhUG
5zAphtlpwsUKPZ5xBtXIxbsir9wpMM400UsI7tky0vtbVKQqTBH2y+0EYc7vheJ5
5kVXQrUltkTqW2UG0/8FSAkFKtyqeAyqjbVwPKLu2JNuPBHFb8cw3Egud8ebQTHB
UAPKYA85iuC7rL5gbUjFMRR3Awgq0s9w5L1spvtEB5lD0CcoIkYZ77kaYdb9WgEr
wYAnAjLi2B7fdf8GEeQzbs4ImzCjHoS7x8ofH1+S5qIgyBI7T/D+DzIG6MZNjf0B
rlT35OaPrgOSaRYi2qY9cnOwoEsLGjt5v09SxVlcIwxhqfCxVP230c4CqoHHJ8ll
jgI7DNwKyW8PK0lVZLWUDjmF1XDgsDOrJ994KM8v0LeEcMGFV4d8bNzKg79u4wrs
XTEMZJoqcnpiTZ2Cd+bGfwFPM6M9NIxixifJ226IJSQDCU7uE4uyCo7AXwfSn9lB
BTMiV4mCwanMRky3ph6+qQvTm86Xz+HnDCljJ8T4tfEzvu0Gt12awKV/bw4pzCiC
h/tDv4VpIqAvmg2BFOaobn3BiYNNgfeFsKrVBrpqpKyua5sTPPj8IFSSMcCGSQSd
wHuDn3/H6tY7OEqv/vwnk4N51WjEhUJ6w++k12kQxUtNYoDPopt0jlKjQ0kNPNGu
B6MIoUjxln4GoYaYQGw26h65j2bJdg6uYMpwIjSvBSb2tjK92jhHHVOXwXxpm5PB
Px1C+s3kUX3P0w099gFF4xbZD5EtHP9+oSZjPHYXL389I0lrNiK6K1QWWskriy+x
0JH0MNzaIo/XUK6uph/TfWXF80VtKlT61d5e6PKJHNdLdwnutr+anmMj11sKCn2i
pjKlKcP8uYKdZVH6uoMIKVMwaQLIhUEUu+PQ9pWVmaY/nvJ3tXJUT5V7mhQckzqA
Nvp/g4dE8MMDrsw0mzNt6vU/MPGnA2sHwVG2A3S59h682CtT+dvY4VzV90USP1jz
lPwtBLPsDJzd2lkHHCJzXGDDinr3KQtmefx+7Gi3gvacr2/Q3Uo4Tc3VwboR7Fl+
dWBn/yKVteTuXRlVxAXh53eO/2VqpkHsCIsAQDa6uZfyOWvGL/OA7m82D/SEgzEi
8yWHVwSWh+fLTVuB/0YT2NXro5sDpLaZxpbugIsE5pzWvCR9z1fdh0rQeFDydXWb
lrd/iFroFC1riWZdds0g3tLI3wvD/zlyxWzvXWEMMY9qClaRUghpBTMD68kQ77PN
AL5t4JRTq9M7rEXxZsgpocLP4LmiwaV58972xCO113+04aymgo5TbdxOw4mtDhGJ
NLPgJ2BoFDPCZeAP6NmqJwozalmm+CHGGHJsmizRaRX23+PMGI4hoWM61+sx3aU2
vPXHS1F0qhTVYlRAqS/fIrDgA604UaEFNvjY3/QC7M0ubsUX3sIiHiKNozMFt9ye
GqwtStKvJK5yZg8iQw9CIw4a8UaMkhozgyK3QKEWsXMt8YKJzn6uiR11wtvJ9wnf
4aL41xR1ecKvZNyx7cU6fDKV4M4SY6W/hELX+MG5iSlE5pOAxuFW4mK13+DVuTZg
y7PCWXk+lVpUXgeoz1GwdhN/VJlKjPcXdJNc+xifZ1jWFZO11J89bippU+9b2xt8
t+C6ngCDp1zEM2ASUXAZ/bpZgaXGb2zMbq2VYeCl9Rfn8/rHTiPx9q9vKvdZyU8b
+/l3ZzD45WM1ZqaVmMgkOZH/Xdu68O28dl+ha5i3Gwyv7XKoCGLyvIb9PXFc0VUv
2T/Mn5TQyLvrRP2m7YzHSKJoNXDZdPjg7mSI4oEYPEZvkNG15Ggtax71lje5WJad
S5fxmd233xAnfgOh4BUE6/QngrCnRJ3EuXHni7bASPnBYM6t1JbRihx2xfABz31/
AXIplymR0vlxTlxozEm6cLHjfYD/qy9mfMrAS4z/hCofPuPPm9HRQ0DmPvWS59ZV
qnajo60aXI7Kwqyn2ytVtUMxts1KZxTT1zkvRK3k8tsd7/8kLyhrsbUNCbtFZKcf
U7e7j87XWF5vXc0vulqOXXBhjihBpBeMFHxEcuuAV2iSII35GuHEtu0zKf5pavmL
csKztTzb7ydYpuMP8IK6Ty6NNO0pLEijXUntQDdmmObdp6KX1ZJxLUzszN3gyBI/
UAsk2jR0/BBzujAO8Ka7AmKVNXtCxCPz19ng4d7ujvON3vWhc6ne+3HZQj7BvWUf
cklItJwBp5Kkgi3GB5W9jDoLNVOzgWCTMH5HOMs8WfYCyLaOpPiBLe2Ro3G0NP5O
eoqLbD/eq+fsW5B7S7rGg2+pJsZkOFT71YfjPFn8RnFcWYdw2D5u4NWLTC7NzQCP
cwcv1Z5vk4RpfXJEzEgJN1W8knQVNURD5jEW3rik19i38fHbcg+RyRF2xhGe03C8
CWrHNedQWx36iLvbgTIICIyRTHG1AcX+ZkJOrPqJ+oNcyJ8RC/DfdbLa2LH3x+P6
3uSz763cJ1H94adi8Sv2Cyy8EH+/cap78ExqCNDi2IIMst1Rh9oYFWpCmbSKK3bh
dxFolWpz3PotAzJsN1JfWJnqhxX+udN1DmVI2OLbmsbYxLTieANyGRYB9E0wZxQk
oUro4sGlimdc9fKtmiIVmQFBX6Stxcq0zyfSM6EUx8R+7FNP3V7NPJZp9pvjNd8Z
3JoDJ5Hz9li+LkiPhp3n4kGC5FaSn3RDvw9MOcJRFBz+E/bggB/7T53/mw0lhccw
p1RGMPRbMpRbm92xihMxmnlv8AuE8FJDe77NiawnPowwHSqxpTJxk/IzHc+VeNGb
mffEixZGXdYNEujQl0Q7ONE/lrOD4FWltO6s8KQach8h8HHVkd55wJNy43z5LasR
5mzybZrw/Wd19FZXznq8TWA4j7BHLG37TTBYrDQc6dLx251DM8gPbMwoNl7ukPsR
FTcZejZ1a6UMbPAztY78L5MhJRgnBaBuC7L9+3DBbF67EjwwIg8cUsOXelDWnJ7O
S7jTzpZYKcieds5u89GJpTQFzbrC7BkDqsndo2JzoECHJS3W3S5Z4EQZuwOZfb73
55ml1rRK0yZjtZybFd+SHEGnv3ip/RusYXzBb3Wi76dghD7/nxKF2EKQLPz4iI2d
WDJZ8Ay1IrLu5lIYEdgsjjcUsq4maoN3ffVdSssJl13gt1CnZV6A0yvc6Sx0s68u
PsEdavQbxmeJl4xtRlfqHbkBleEG4Ml+SU2jlioKz10AATjk0Zgpm/wqX65CRSAS
/ZeOiiqK2o9vmNng2aFGTVBLCSXsrqI5o0OHlIebA+aG6sfFmcfNleu1ZuJFTgGu
CF4KnKcmPE8VIw5SiKazjbcZmib37gyrPbQkMBHIZHQfGVsV5L3TDsUEMFXicLO8
vpHHotiEBGXMOqWoJ1uosyH0orDPYXhHBfn+aJBmhnoZjTqVHl8+mWRvjIf6Rszk
hj5ByW5J1emoPD3BUZqjYgwgUSdwY6JUcEPi0T1L0UonqqIaGmDTUf50V6z8mp3U
QoIj7AZwd6ffNzpmOxSK55mH8YxDYeoL5gMCbCoV8x8A7u8+kXz/ZirZqAtjMuCj
XMvMsml6OfW+2iF5/PyaGjwffK0k376M7pXD4x0NnceltA/tX9T74quC4LwuN8X+
HRhQppkumW/7dMTdrChpcjfJjMz+iqrMQbaXGQGpyz8QQ5am5Qleea0pkVBy2syU
+bSr1/2Ulu5QBDw2h3Tq4BlGXR0so9iMh4iCBizEdMeGjjdXXRZgCUsHJYhN5ca7
SIabi66QYI4hBs19t4a4XaalUx/k2qjspD0AA1JIi7tTqRMxByvwLxlu+d1uudgq
phCTjFpUI/EITWBkQm7vlouogRGFcSSLmKEz+gzDzgy+F4qEXS6CIohQAvPCONan
r99YIQEUN+qLgh8Mu+Fz2nzde0VTgqMkAdu1opEUdymLJKTARqa2SkrJjsjTb4tE
haGQRATOY3lnVNhz4mnffu0dxZ4UiQ8Q9F6ZlXA+vOGIa6DSE67TQC009oJ9gySE
Uh4OS57w+Wld3pOrVRn4znsukVHzI/To0//1ewhfN+QrXe2+jCffwOoyRyr7lt1p
f9RsT1xmYlSTJQqR6/7kmqLDZh/82jN8RvAsNIx2aoLT245iNqHXKUVd4fnu6DR2
1m7hgC2a0O/xpXbS7FmD3MrSVmon+1Y6SnyoFwBUTZCy0QjfcQSaWjTFwGBwvcMb
H3ZeQWrmRqAljhdfUKGSwq5e25YiU/K8PutI3O2t9ru14YX14u1Q2fe56lPaEUEi
F4rl5ATVAwWwWvk4kuSEV/YCxgE/7dvf+qMKCg40UF9Pjvsp7/TQImBy6aTS/R0a
JcCjRzS0RqSeTJMoVsNOpIKEByZjX3Vt5zsz6XYPKQ9onYuSftNJKfRZTtsXJoay
gWaNtElEaou1uBpKFKyJ7XwDoziRy3OEA/lzb6OH6Bf/O685dMSzzeULZukUsE8M
BJHdyjWdRI3G/KoRI48jFv7qnSHvrYfVDQfCti3ETqV1ogBpFFBZ8TAP07hrXdDj
T5WVPd/ovBSg9sghK+ngRE8FAlTU0Dh3JRz5da0yip1GTGo1wkXpf2rFTSQDoK7S
fHGwF8g4k2EqmtEsNmy086FIjcEPkTXqw+NBK1xBNrbS8QfoADowci7aIjCOldtS
JiZ+jEKF+C7c4OEH0otpDXgMH7CUMo3sTdrLuXrH7pjBLynYy/B9c2QgaTPBBOzL
jqlqkUC6Q19acIQSg8r3wYfZnlh+1jmWqvgdFJAnuOEH7r1saZMmloUwlAobtBQB
r5EOKk5H99cDwFiCy1sKb6vmZz/tTw8gAxEBCfbTia5RuAPCo+Y5Nnj3VV1VVU4g
UGOqzSwhgZI1M/p0ssICSFqvQKJ5uIgYp6IlmMHR9TWTJU8gMN5V1zkdpjOcqIYh
50rp8/n01V2qq2tmafuPeDurAVy0MfktTxDPe2cXtY/3nctTpL5fpK2NOt7uk3Gh
Vbir6WazbF4muApPP64j15m7P83yPs+LrDZ9osJFwZ9YzzuSltjktt0ggIhDDv4e
bZ9HKJLu6Zby1lAon14gdc5Xhow23Y0Dzgv2B25vF4wmP1zo2Uh6MqbRVv9coE4F
Oy0GAr1IYka6Dm0XG1tCmyalf0zzRFz2LX1cvEqmkWK4pTu+Ab1+hKMZNqRW4J5L
IX92ZX9yBTKOP7HUoH0VJU78FtWzh0rve9KW9pOtAdhdRz0HnelWTIDpqemQz970
Epfk0F6HiHzc1NmLI+frCn8tcYDnsXlVkUx7AIkIeXJbpqqoWX6Wx4rssk4x1JO9
4ImVj532BoxsJgRlPeYf4T8WnuJ/HLCzGz/HKItoRfIozC29HtoL1rZ0ifgKv1nl
PTc/9jCrG4dylMfyxVvWUGQC7MJxwPt0zHBXO636WLcRRAMG2f0ToublCHQmkUJF
Sfla01ocxkEOBt8B0wOrSkqBIloTfAYS+D8hGDibhYd1my6LdJRwEaXcebwUOUXP
mvU8OnfPMuHvobNdA1X8El0muC66AmijSQMfCZ+X20zN6T28oHqUr9nPXBWcJmir
p+SPuvLn5O3qIW75qCM8Ci/2otjP85/da6nEQVXlsgD00AouADKZ7bKUdICpwMNv
xwzTTolWwd5Ks9DtIIobINQSO6T0AavFhr1ySeqhFUCRMlBw/WGYS30cG60iwNm/
1TbM2WzDQGbqnL/McMGjz39ArIZRer/Vwsehbe1d508hld6iGrG5dsbuLoKfz89B
zvqYPe78mZ+X0DLeJPwxUs/E/mrvd/o6cEV5RO3U5lFSo56+5QpkZHdM7wkjr3oC
bSkrx403TWMlT/9rJ+DLH9mXCAEXt4t0myOljVB2nQBcAwJECZA+SlVV77QBRnF9
WQDQS9Gmfx7aozjwdd5SUY0Kbxv8nUCO6t4ZqTmJK6ImTNPYtgs+ntLdtrXiA8n9
CVOaPp0ImfDyVGt0qHk6vLWdBgnCZdRPQw58nQp2v7HuFow4GRJSNjDeWL7iQ6YY
Si5Nq3OnZvXe2ACPTNev8cSNECRvRfyp/4ppo8Tv+5TzfEe+IzReFvq3zpUt5NYB
`protect END_PROTECTED
