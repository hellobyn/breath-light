`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xG1RlwbbLQHXp/kk5fLxIQLYkl+A9BW8SsFpzgQB2q1sm5iCc9zSSPhwqa2JkgkS
JCsrTg+rqLfB5JolRTxMyaKu/mncosEApnHKxK89/uEAzlV6PcFGzOMpPQTOosCA
edToOu1pq18t3wq5SF0dKVIkFTsrNpblxIcek/a/G7ziv2DHdl6doXWTNiSwgxzp
Q6VTZQAEQVdm3MXudTkpE4a8KaqbsDwxNJmu7aQZqCz4Lp1XKyavl9x7cjFUlh0r
SHWpTBJC0nS2AwY7Dfim3g5n915dZQJzjEwpLr9sjmxUEBsPZJwBvz/FhHSyInd6
A+KmvXfEbS1DnVMsZv/kdy4/xvKSQwNt9KbohFRzt6spnlwsbKHGtwRt+GQusD+z
l9nMN7SRnttdN24LYWhLW4gHnT6t/uroXSBWOWAEVWguqV3dpJkJ3R+J5PZ65wDi
mAHDTF2QBPf0aVBMr+f4mJwuwPesrKcAcpTCsxOsbrRH+/3dJpC0YuzzPwPzBXhv
OnOH+0zDJOp4NZHs34KYyVJVmXjukBycmX5wMNnE8E+gPx0T2dZqFSWxIEmWOl1l
+M5iPmUspKvPfAF35mU48n41VChvL4iU0/o+K8Fi3ThP8jybC2LKnR70Qz9a9mbN
1idi/r+FotBw/bvG/lLIALBCN56rjJJ6UOJFFDs0O+obGxoB9dn0GXuwO4nhFLDa
RmSe8QypZIp+zAO6fNoQE04IqfnI5BbMZEyAnjRkztJSHnz+u1ytmp6leUC6t3cr
UAc1Xbh4AjX8aXjVw18RpAN6o+rBByjtMsOWhyUp3ocX65ZthcFQn0HaE8FsGQtp
u5NEzWogUrCCrine+Man/jK1vL/PU58yOMpdaijd7/V3CCcfuYS0TSIJHG1ow/2u
RaQNY4hFcvsBSzKeyYXuJTFpRQGGV/GePOIcFD0u+WwmB0tGUprW7UoavmwBfDsJ
jPIrp4dCTX+cvtP3v7kCd/PCGK4Q+D+Y35jKFMdoZzZRRPJ8YXlrejsXbA3X4owq
moOu4tlAfuF5AJxKBcW9hWSFoRV0Nkg9cv/6YaE1VEQ6RCcpo+6GQXKs3Kzb7QVG
l0MR9hwpxFA9OjfbtsuZrIJ9bdzrOM8nHuzVZXUe6mtWEJJDwZZV+9oxy+2ElncD
iSFnGT9HNar9J90qBKN67Bim3adHpXCp4oTVyuGHY1sCF+jXJ3/GufydMc4yICvI
Byl50JJtxxR6ScGYRHYp3WYln3yRKB2QFihcZOdyhuttNf7KD1jmrxYyswMbnH64
UDP8POPnNEXbH7iIV6v9xvKEf7At1DTwn92pdP+t8ITl70TpJPZFXGbqlftco8CB
U6yo7dVWu6mnX0NuaYPMosLs6VOvFGBWs6BkHTRlO64zJrtbwqv2zfwf6XMRpYbM
Ut68wJeb5ciK3AkwOccsVNcGEmOOtKQgZo9pO2mAZBxiG/MKxF+j9U9Fomo40IKk
IHPGB0geb343IrCr+McNdXWM9NZjGIwgiiZnlf7BQAz7CspIHzfxv5Z2znX2XDEK
jIT7aUEuAcwIpU2FNtFmNScdMLKc+Obs8zoMkTnlHfg5SfiahWniMc2OcRMQYVZ4
ST6O1IUnOta0DcD1OlxgxfBIUg3wQ8XyVAieyyUHu3LMAuHWT+HnnH+y6889S9ef
Nggq0OrgadFgFbupnf626Jz4CVHKK9j1ErcJIzlO8bYhUCpT0pnrwBZW1nur22rp
Yqr83t39eovwhL54TwGSfH4fPttoHQCJ9EXzAXg709Kxb9DHu1hc0AdkrMP22vnI
wsbWCHHZXV9ABKGtQ9YA9RMhL41LlMsqLf2Jrgc/0QoB0etvCUO/1dxmk2bBJ3L2
ro0liyI7gsCoK9+Z4/eJxTKC9kQTjQAkE4QlQzeUlTOW56/s4lHae9LqXuWjfTHV
EncEqTeBPlFwSbJhVYtro5tkUhVcXVZJDzIM2GIo3XwbCphPlOFgfnuVn7w8ulE0
hnxl2FEO/uzN68WO/0781zHvYoXQF3HAIHm/9hTgHmZzbfwT7mmeH52jC+Q1Vrn1
VbuvVEATsCJ+cyqfpSXgNVwe/leOLQuD/HP7Jb441RQwpQyI0UrI5bZ0Z8y9eeJR
Dq2AG3mFdZDsFVk9Dk1waPK+Cn2b2oEVVDQXTWQkYytoV6mRzFEEBhvkffXziMaD
ea9d2Y4cW5jW3NeqqpZTn5CWn/I7BqvkBRkj3NRDSBKdKbjscQxJkZmHmCnsKAdz
rQcGDNxDJ2dN0NFx6HPHA4WyVmm/odkRGWbDcdrfHQI7JAZS5zSCxCfQ5o2EiOmf
+8Xk7I9kT2ui0Js2lFYTUiFZRCcbOAJzqU58qwF0ZaUnQqPxG5UYjRwEm//Q+/n2
47nFVM2lGFpviqk+5GNsr1LDt/d6cw7ylz2CmI7fUZATXm7aYz7f4qYA9VtsooRo
tJod/8lNs6g2iExyJB4zVdi5LXflMuPmgJcBh19jlnu3Vj8sVetSo5xawzcBxs39
K8aOiYApU6wJDceyTdE0RaNkMXBMYHe9jemkcTsxWB4IUaayMdrWUoCvdMpl6ItA
ZtJ6XdCvOLGgwmV8sfYD1LMKI/wLxfDXg1Lkww9ZieWkk86APtGVfwYaJJ0KaoJO
mJz88fKyXXwtEWvxy1W2rMXLS71P4eiAxd0hcC7V1hNqoATZ6LCj5bcqWDRkpnRQ
OaJ1hiq1Ghx2Xdd1h06TUam+culz0UUw9C3NR1jF0aHiv0rXNrE6C2/KQk5SsSxt
t6Qyn9lIWJsgELfbaY+r2nvTTYWcOpEZSjIQ2AhNZETIvAWX6FJZ4jG4J4uB8EyO
vcOc59JQYAezTuRYrh79GE/euauEpcJ8g3uzZauaffEtW2pLhRX1VRCPpR22/If+
rz8BoQwENw9fbWpxW9mhyq4ZCbG04tvfUkGK9hHY7J2qLQUe6GzRDGJeaQvkYd3K
RcQwBCbKTHsQ49aZDLqZXyII3tVC7eaL0ilKkLcYjQ/MdvCp3yXRTtctoYXX6RfE
bwVuQC+oNR65v6pPhcgM65yMPyfZw/1Ek0RpiXydKC8ftou5g5FHT84mVTGh821P
9KQG6ecEn9YDOMbsnhzFjwca5w6OTTaTkmEKHdjQbeoiV7DV6kyKSM/LU2zX8fdw
oNDws5xicaV7o7Km3fZdncoRv2Kcu7R6Ky+LAR9ZJz6H5jcN/tgl8Nu8nqTFCvAR
UOJxN7/IX4fJl70IrpIbQviWy4/kLfRjELigYM2nmr1KH7hoSD+eN7bJd+4CLpDy
RHwAxrPglcyDZdmIlZWK7Z285jwvMSe+9EH145UCdYM=
`protect END_PROTECTED
