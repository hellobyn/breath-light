`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ls0cDs2vq3khl11OhTxza1z1IlbxL53rzhedK0puNwalLtA1gWYdR5w7pKy8hlV
IsMaEWeENxCMmg7nOUtGtjFUHQFLbSA1OG7dDg2Rjk6ExfCyogp26x1ar77dS5F7
lEtTIt2FIptMS5uTnFe6QFVzE9ZoNN+ZLZmgFcTqd76O1Bc2dqjNTv5+yKbDfXJ/
Np1DgjHuDTaHFsK0et4DYZy0iaqumNpULpI7IADQ5zgtKCWoCbG3S4pgFVHNUSBN
Js07OHioos8g64J73BPDM5+YJFEknxOYStcpcfDmi4U5Y2x3aSM456L1cfAQWsv1
pWCbSl2fyrAO5WPKEiEQ/BIKWOv6PWGAcV4R7r2h4A8jN3wTjIwvYOWr09y8p2+T
utG9jnX3WpLQkmljcm1MoztnSmEcuS1fK/2ESCqAHe45/qQmQe+VPr6Ayv1d5uj/
eHexMCVQNu2m/q3jrp3YGkfsRNIUtgL+/iHibnmNRpBjiVyCrS+VUAFjRBRsmvL/
piuVqkfBY8opPNN6MTj3pzFv1DuddV5PzzlPU9QHlsbG+2qx68BSJljKQJvZsGC4
7ptyPRS9yimfp/TJLWKcEbbG1+O4cnhJ9spQhg30OWVeSjjm4E8lAMsyycul0QhE
GgS2FHZPG6tY2aDu7CmNn8KrOlUzTRp1CE6IG38amTK+pXu+E0CPt3BpDDqVpna6
WlyVlPeqt1ytiS877ILp4FQujt7IIpfn1G8SM1WTEb2DbaG41OuHNWe4M6tXfowt
ManBGJ0xgYEcAaZoW+DKqu7YPPI/Jo6Xyw0MFTV0fE72K3GY1AQd6Xh5WOeXft/0
LXlCVLAi2qy/gGKnxYsRaLaknBtOySdFWkZDcEExyd6YVfkaUbszf0tw9QLN+omm
pYocqbYRc0end68ExnwIapQj+hwuiw6/9DNaL99FawNt6LH647LquEqTYIHY2rPo
XGIhZ36yDC040DcjjuLY63hCf+uxL6CpurmOi8lABcQQwpdNBrw/EsoRoIMkuKrn
Brll0sb/3nrDHjw3G9nb3uAmLIRJWPiLcVmaNU3MTEztpgpeHNZ1YzxNZhsFEznR
TCFLkaExYP4dgzT6nZ40GFkdvMsUYZKa2GwrADE2sBwWnEwyub6Zu3jOcdw0wH9P
CYJ9WAZMJEVjTsHXH/+RNJcqpX+PpAqEtHLrHeZdJY1g7S+cil3u+fbu1KW2uqv2
B1q2d0K2bOP48SfIMrN+xqeCh7e++ZV1sPu2mgGQnmnEguJT0YbHxiOyCne9kr+a
i7ETzgmBql2OPXXukzBoEQ==
`protect END_PROTECTED
