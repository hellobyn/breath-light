`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Msl9D0rOiN+bT474dXJBZCXaKIE/YxBDjvSKFHwtqsEEmD8t8d3Fb51cBsLPoV0B
rar4+MbjWbIatvqxb7eSFoUHwkzeFc9n1+69Hh4n2J7QwcuefQWSM+0As8GVOFwj
eqI0Or9gQnu4X66c23jqlaRWFIk5v17RC1ebl3MLVZWIj5/LNJzcNpPjmCMBKDJS
fEIw73amNoxiRr8pZeMpb46SfGv72Buy0XgyW52/IXbe817OovcJGEkh8/cH1cY8
dhcW81x37cx6AGvhDN4LIbuxxRtDakuPXyj+nfWyBT9PtVNkS2VNZ+PAzqJMS7mq
J3pwuEC2g+Kc/A2G2UDwn48/uUhUtOtbivFbzWGiKtMD0jU4s7XeKrowE3UgGFN5
3NGcMHdEo2JISjAkZpHAFRhAqrAeHrzgWPJoSAVx67HLHFnRU35P3fdjvQtghz9I
KfhwvNVNdyQsVprC6EqFEGvObHnyC2y/8+Oq6+U4kJrFXq/2kA2PqDLtO23Yf4Ie
VuGsZYOHMs1kYhHHGuusnm53JWtDw9EU7vxD72nr0+8baAAujWd1C5qM+ib+aOSq
xXLjCEVTGi8Z5EdEs7m48ZrdK89u59GSN9zMefFox1LRIngCN+WrWAyf6d74Cx3t
zUg8FB52HpddbmjiHaANoCNjrFqtMEqwbymiC1mg2U+QwJ7Zg6KWKUlmXdiinQ0T
`protect END_PROTECTED
