`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
373GMXgnSbnddObT384yqdeheH+4gCf2iwmTG6EeasvaMve68266KfvJj2sr0wGO
5jx+LSbxBZEk3EWO7l/3vSVdQYZfRL/wkHMRR/Iyc7ERQ8lUgcIO8un0T+qRzBub
+TyVhfFZfrKoWvcp72M+LW0LmK9j8BV4gOW1350O+XgmHy8LzUdntgTWzIe2B2DG
Zjqy5jK6V6NH9CYi+tX1pcFn+Z2WQnPETDys/XSJ8p9cGcebnaD5L3oiPYjA6BuG
cG1ntS95erVJOmwY3E6ARp48QNyBt83jSPBPoZGzMgBBiQq9yyLEE6ewTymGPOBJ
VhuCm/wjxH65JDo0bgQ6YFIvYp91BeS4i2PdtTZdes1Z7NBv/2wBtQD1LcfJvpC/
r8VFaQbA/vYkcZTBRwLwG0anz8s9btB7xCyTEy814deau1cLUOtwjVzlep5IlJoX
WW+dK7KMBb5Ei2319k337mfAMqQbePN3QzENT+G7EYZY6/Vzf0ddNTyepMfgySHm
vI7QBBx1onsD5VKUAUzEdVmBnwK0DqTNRFD+jIK9bpXP3/rhTM/rrabYJQFVn62u
DVzJMR/NQmcyHhBqv1iDVqDVz5bXiVCtvp5P2P0W5+NgUUq4yAAbEhhvKy3zBVzU
Ulire5SCykrRD4xvM7KdQZ4rCIaDHGwnD0bAw/qeX9SjP5nj16ykLdIpzWZw8Jc1
sMhopb3McgTMhKrJlfMuSVICC42DhcjAsIJJHbYwsiOWATxHxpsj2UzW8AzqrUWV
+FUilfbtpgI93yNg3Yl95UjUZeyXQ/8RjFJq229hkcUBj5WIjGsW8DXaC4R5XPeF
0Z534IbX5of4yiKoOe6G5DXcQK24T2G88FHsYc8bix8/d82SrOFssEccQTteFu52
azvZGTOchWQ37A2/ZbgXKhoXNGLjV3evoiHssuN0avLC2Brc8DsVyglVZMZxhber
`protect END_PROTECTED
