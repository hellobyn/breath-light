`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JPp2LmXOw/YS+jJRMmZVh5jxeKK/7jMo2oouct+BqDClQsZpR2LYpVdpk1wzigsO
r/QZZAeOTE0KRHefmxs/1Y4o5Vvka1LXGC4QfMGkGI2q6oydstmu4Qy7SCLsChz6
0GKvMNMadzwfpbPgRmNCQWy6WPhO6+YBoUtdauRg+2xyTaJlYJ3rxxvVRjoJPfQm
k5uCdV79eV9DoFDZY1EAnKwBAAO6I0FzcB5dYTS1eiDAZ0iHQUb9MdfWz+9oFn32
eZ6R8D0+Xm3wqf2Hc4EJ3hfA8WvvpVRftAFstjBeNvyI+TRW1NK0ddVUnBaj061a
GTYtrUulrxp46q8AwMQS8UDfyKDVqwAP4Trz5+H65iNsCCZEg+bgxO+UtdT0ebKp
tPHxG/MDYlyQKnwm9mpZb6iy8A4kZqyZiVZAHlMfeklHYX73+V83wWfu+CPxl/W4
qWVTfQxHm/6ILOJUSncVw2mRQevYfiQN2zpQBLN4xFa7kNjphvE79my+rT5vT0vC
ZZmU2EcRKbl6WhVNAoNI7LQvMgqMlnG4YIDuDAyNjJl4t4x2gYJHwtI7QwMeW3I7
t7pzRO2/IHojvU9nIccpQYXGxWICOTRWYTIPbAikwOtku+htQ6s+XHOnRY/Kkt6I
`protect END_PROTECTED
