`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XsOC5ddQTL5vY+/H+jCtlydHnp3VOdNder90vxXdz//yVv/BitDg0gpSokVn6tU+
nVTIJ+Qes8+R1F8tuAtj4uvN4aeXgM4/xlILUcc73ox7dk4VjuBKdi9CYLRVNDdN
w00IxeCELNj0/iaVBgNMsi2WKHKm9viBEDuGF6FiTtykYo6uS+ICfnoRGW7+r/on
Plo2W97ugQk4MLMq0xRaxo18kA88q7tWRS8illXBR88mTocHOIITrVD3/LtZxZBG
vB8zzCNg+cWDQKGopmOD+gNX4p+ozkLay7wqc7B++x5GsdUH95Q4HRjO3OjDUBQN
HrgYf82kiUR2VXtSHlwwGQ==
`protect END_PROTECTED
