`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18yA++uzgC6lZpMGUSGnPRSJdh2Kc8z4T1/7LJW1KPTP91OkVqUBGGYrho+AY4cF
PFogEADl0x6S82rOgl6TPDolZNi+2LZwZa/yf+PdJHbOjSZQ8NCRKBO64xFM/AAF
2BPVUz8CWXy+ud9eDbQ10948QSvU0ZuuUa2K8/JuvTAfQXJjUxe1EFlas3Il+BYX
lsB05fQDxN1q0quRm73KLdUJwWauf44YpbLLxrSP6F0GGF9Fx6MHff3EeYQaAvTM
moBzX0snaQjB+8kk4L0atwAFXzuKIiGlu8nR5jmHpEkCBYu7aoXf32914/pEkq5W
A9dBZ034HOK3bMESvKXqMT2A04YoTLFtt6w22TiSTk1ZAUu/1as6BwSAkOPgngZz
Ot7NdKILtIA7d/G6jDFSTJdLAcEkUjee2wKVMGssC2GopMlxR5RE7Vk1YDMzsDYz
pgSK4avJVa22BuJtSo0YBQDAyJEpMbSdS6K+QzjVWUNh7TAuPXHcKsfZwQWwdKuc
ScLSggKdXzvJdDW1C12mE4bdbDp/qSN8se3YNmla28IoqGSMJj9NKE+zSVkc2ICN
zz3YU9bxuPWL6DR8BxyJ/pxsyTTkUkqZp419PIDgYbjzzb5mVCPyfJgDnJnCgZ8f
YmdPzsOuoz2Ev2XBebL9iVLSqLoQ0W/EjY5hYv9+Ei/Wgcs2vW3ue4xcuCnYZeGO
h9UeJEMdpia2Gjjthjpihm17RwCeCX4RhKtphYCA7SbEZpjlcmVDmAgbpdzxQNUf
+pjVjVH7Ac6heQOzthVg4fxST7EnwtGElGNu9L1oapt1wrOf7KLfTfZIdUuKjQVQ
VX3+vh6qoIAmWvTs1uSq+xa8xmwAQEFNFaLa1GPv6nS2d+ZwREmV1MXGRs077W3q
wZdIn4TAqntwyPgrjKCDongAE3LIhs7Juq/gsEOPFLB2v8+ztmA6VbZaGR1BI3yz
5Axindys/UAhC21+Z18HYpYA2A+rSxcCKmMxZXAa541LJ98mSqbfRQhmEGPW1kcr
VSf8US7s+Rgh5hRX1RopI8dHGJ8Ag20CujDgn779yMjw3Ga1eoqB0awetvMQEDF4
xmfHwrlIPZHNXm3Nt1mAowPQCSIO6UQ0k7riv6EjxEWKkEixQVI0Ch2C1AmoyQi5
6gSCLLu442k8ZzjxdRM2SNFmoYjXSFbKoeUldQtEJVXK4hS/dJi6ZmJg1t9rIr6D
z5tyqmVzQRQwIQ3NRYaUtdXkRxL04ovDoTzTmB18dgPFRTTnwatRq526dRuNnadp
JOA3YEJC7/v0AQe/KTm0HHRAEqXUcKYSuyVDxX/hj/TnQAVkojPLI2sxLbodRaFF
YLmV1C6aFr6pwZa/aBVq6tFVEB1UdNnKqMdP9oRYu/1DJTpheBqVg5nJPb9kuVHF
BEFrOdUH7D7zt9D5MasXrRLdZo5NqGIpGkIAC6DmEPWggMNQb06P7GbiM0QmA9T6
Fn2a9AsTB+u1KCboWDb7Sy+t90ZqyCD/lTqUDWfJ3aw6E2ZiESFFccu118HAxsEy
UbscGpuoentNUEpSnaqBdYp46V8elLnR6hZWhJTeFoZKV2JgJT6po/zgRx5oE/Rz
QtmI953hfW2t/dacovNrbFS3BfOA7Heg5cBsd+cvhG47r+mD6pPujyMpo064m/Fw
jvodwlW2rvT5wJdc7HVYS/sfsttRDIGOm1svx3B4DKYJvNOfrujwnTL1UnBeox/L
ib5lurKK8OPUQ/a100gP/g==
`protect END_PROTECTED
