`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbnUu2Gjxmsq6FRvzZg0n5ku1Piaen65CGldffihW2bnf5jrP6QCkms3j4Qf8UBu
VDhpjFRJnbof7FlIlkUfJ+md+nqhBxw0g4Psl3ow96FOw/CYHHq+wyUgHFTk4/vM
TED3JjXqqOC6qzTnWMDJU7IrsIkDXRskzD4kTqqJq7Vmhi4Ij9LecWHjgx//ylyW
hqERnn5MLWpyhvYJGTomc9SfyOSTosEJ1+bBhWXbzUZoKFP0ULoBLCZMqTj24cg3
+HaBDn++V0SjWB9XtlV5NKmA7qYD/D+Hq6cFZb6k9G0PPuTY0nvUYawPlSc2PUyC
PkqYCGuOZ5mpV4POvJGQpSP6z3ZfqVR/qIPqyYkAkeCzJQPCKGy0MyEceH3aK/3+
jvvA7nSyMPuuRGHUUROk0iM+kcg9XYjAtxVDL/qJShSqbeQhaHB7q0aw68Zf+mj+
GvnfridiVBE04R3UMxQrmeDRmUhfzOZq1Z1VnBkPIkZd2jSDjkKI5i2MCh4Vh70P
tWFIoffkQkbO65lmjkw8yAADp+iC6owIrdIU3bQXi9MArK2gpjQlD//44asxBVNL
Jo7jumKQWBtie7+tZufLwQUg7FVTdoDKFgXVrvotUJvw29rzltEWrQJ5+MWMWoSn
07/uZsIGKVfIP5ucwaI7Mc67pD1y1DQcG1NsbymZQjZ4fINaQigaZtvqB6mThpL8
6d5FZ9bAZLjghRbNVEbzGvmeCwDq/iFlBUm4JYikNiB65ISdw+LJOCD+SaySN3xu
SchR3yRMOH8D818WGJwqPeAkpSge3DdIiOMCSzL0q+olpQCtthSQ2PzjLOGHAdTX
Xz35nNEICcjVuLzGagikLw+uFTr6+i4WGy9Wqe9VNBmtLfLe2LBxZxP8JepiThzU
+sJ48VTWSMHbpNR9rdij99MfP5YoWs9YlcXpuxIdqfDENoMTzsmDM3MlOPVuxe6f
aeS0bqS9Oi0uk3Zeww3irEIqT8fqkDq4tq0RQjjvp6pZ3fGtKVVj3VZpBbyUEZcZ
T2tlskYvOi4BgzUertGZsk/riDWhDvarYmmyKaca4rHt+/KfeJTZMR0ndGSjbdMp
gsD4v5Gw5L2S7k1EY5GWRF0BlSYK3IYbLn2NeuN8worjmOzo5M2psoI8cFPAiK5V
pA2aSJFsls6hW9P2J9cmzPOzA81X+auZa9siiS02Y4pzkmSjAaFVFNAlMXQCQxyz
fLWISmeGgmgsUzlTSRRrpS/lJo2b3UA7ObxM59LVEAnt5dDLGyQFuqSgF79x0rYi
hHU6kG1miuuqX1r/+q7kRGOPxCrJSdFQJgp98KC01QLeicpaWsNUDuP6O691dkgT
IFa4IxtBy//At8gDXRTIkQnWDfzHPDRrp57CvPYFuOCIzdIs4Rikb8GnPVtoX2E2
VVjRmfnT7mBqBsXZmuZs4lecpfe9sM7PcE0XhE8KtiaUpSWN9NpF2wQ5I549nPeQ
ZfmUOz+oRUd6IHmSSMyOs9KxlYNnLsq3W55fAnASdW53lpWY/YluHOugM2/+4d8O
NGhGgyq9oR+jQHmiSV4I//jZwqFMYvzx25DgUKtl7ox8Bx3x3/wN+v6sNu8eTJ5a
66Jfj1qvbyicZtzCT+XZET5mm+CzY8h7XB6MzalSKmzYThCTryO6OIcBHeo1PaZg
lpLUcfNP9yM4sfnhmyWgSwXMjRXa69KQDr1qF6K/dRF5Xg7+TDbeyfC+qlJWcCXh
AYV9eYTAEkzBdbxJY5V9Kdyf7sGQPhnP9UXCI9W7pPRD/nHJbntL2uRLigOVa3ZM
Umx1Fw3y4Tl9fs7HhmtYd/foR0ycLrQw4VHVp8cP7QkGm9oZyulRFYqFYEENvLl9
bhSKuNQpFuWWWs8pS4je2LWkwCLbS3GgghbTMWkoURmMPgR1eN0r8eAHRvUwzzjL
VjFFJr7RmzOnCrFabAqiDhABtjkBzy9l4/v0twXwu7kRK1d0FkqbLzSYmyst/wsU
hm9MTYZDZR/vWKxxdDvI8cAnta2+BpqBQbv4BPtb4tVWfpaI+dB13juH27Otewz/
ObyraUi5ETs2GK7pRb1tq8oje/IvzmXj5z41eeV0TX4QfxjXgdip4ndG9CM8naZl
DlZXQxjmxBQhqQq43wk5d7GRMn+87xgGOo/V4pMm9+P4e907+MIASgB4ewLLRm4U
DjNDCPT1pUy9iz/l0/TgjJssKoZH5ptL9La5kNS6a+p2EH/jHa26aGhDyRrjT3yg
Vn4knhBUGWIkWhw428h6caTmh6PZyLfnP4pNoj6E+ALXI4QfImLiequCc/CRxgDe
Xcmn8Y9hv0TuKlmWp08BhlGjSHxpULb2TQOmys5DaZCHbNp6gnF8QK9ZmJsuMhfz
NTG+TtbPW2gMySv+6MWzWDNUXtKFEdq2cEiPNLPnIoTwod9DIx6bE7aq+BjhZ3M9
artSDjt+ZYY6zhfc8s+ledD+Nhk0+iLX3l/GIeoStgnTgre09zFV+WIokggl2W9M
gM9bcRyfG2LEtEcIluU/GCU/YzhkOsJkHUJCVADGQBXNBvmL5zuIcPWLOHnrfJiq
Jxq2kbRGZ8hT+74ZC4ItwFxnCv9y6tEGloZIL/Ax2umC1XFzvuLISPHHqGRUb6x3
8ltwCbOCplPnIJZ7kfQpzFF/PSnrsaF+bEQVOhhVAWIdWc64YIV8XR/vOYATTZtm
8w9f5xjpxhp5mKYQrZ00V3SRVmmbvuHjr739fhvCsg6WB60LIC2gRs74Tp12NUNA
NtcXZJxdMiTbqaurUOsdapxKyX3WkdQhMVOw+A/Mzq8pXjOLRbfyDm5PBRom9/4f
W5RXLXm8I2vUJB2gSYvqRdIpr5Ab1DaXlajUYsP3OFXMR0UMUWsL3V/P0bG7avVD
U4540GclSyTo18mv7Y6DxUwnFs8qDBOciEZlj/v2xZ9iN9QOPbpxQt8bGynn/ysm
uShTPVC8jnimLU96HaWG0DG2fQjJdRrrNrX/2vEutAUogWNKd2hAc92GDahRmoJO
oyeU4aodJFjgsr0liHaNK029LOD9guIqMEvu79HYIzzki0Qn+hCGgDtPl3INy7hr
wneMWxvRhAvAfs46np6/yB/GzvlK1jaaOt2wW8ied4KAYicoDzF6GyuK5Rw7Wqvq
FyDYR003tDr4pyO9edDM9SnI49/tGBOJbSv6pNAfRyOHUjoRWfswEbetnCYMJYpb
+TwmUtDOjL/MjbqAon0sWOmFmx15Ulf63Cu2+97YFg/cKQLa/uVumUqmBDKG13xy
riUeNp3Jbo38aAFdj7+TKtXWmlxIuWKmBzM65kWMAvZPI36/nxZve6Kq3EBQqlF6
bU2kLAV4DXO3NSF0qVzjqEvrqtKKOs7zjeRfoaKQlARH3RlkgDhe+4r+nrp+P5zZ
i7ru3WlvnntxnH2v+fu9C7QRapM33Jq1GC6rppTnQ4OKSAplxjt50l5WYNwQYbdq
PWeM7HkhcWIEN1qmwhqoWsBppFfPVXwr+pdChJBC0l4=
`protect END_PROTECTED
