`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vE1uTwhTia3kBt+MRpbsMKIlCMc5FXYP1M0eQ94hx/20zIQhK5Brvxv4wY8j8PDA
aqn3B3YGrQNFIxAMH4Wl5q3CwkWEmgiWuPNBnC5xUDU95S2BFQgQLcbzaPOjt2Qf
KhplIIHFyVxlYXJ4PwzVHuOT85zOE4Sz1s8SIiUdzoRmP4clt6jSDNcqp/i3ol1J
MFWqUBdbn6jzksbIw+VOYNVwz4zeQA9QTCrbOjkg4kUb18tLmIeaaJfGIo3D0zxX
ot/IUlDAsAtHGxjKRAcYkM2Fy10IOJqUkbW1h3ylx6npR8PaEShxfvcWhGPO63ma
MkAhM2WSF15prF2L4i2aeEkMEojjgUB/UcBHja8PK8QCG6l0VPzeDrvM6ZTpv+kM
Scm929C91HC8Kf3zLnrfOB9qltaWDAaLpY/+sQe4Y7VCBoaJv4CESgehjbdG1MRS
dnJk1sDmLEc2gmiZawdk57znERF0SR6yr0wVle3kIztYqIaP2fWsB2IkO+Yy7H9E
1j+uXAuIXBFK+0rMlRFMRHYkPVbRUlpw1GjM80uByJTvbf7Fc5cfqtW2geNbt+O4
awkgsU1StqosbQ7snPfzzx6CwlFYYTwpOVL0WKnYC92f9zosRuGzS3SY1D23GFTd
OSB7MIGpNN28HohTvj9WtxwDMtjAl2oXudXKmo7+07MAxhM77rTZF8GA0qzjwuSl
IYiq8tgThiGr9A57LGo89DEl1nbBipiJxwK7jdOpwVmcvprPRqzFyps4k5RdiV3K
sjDz7z2yO03zsGvRScCgnGN5NDEcQwgFD90e2J9ANDpfQ3STUDqehYlkdks8MlLB
0a7Md5BdzBXObRq53oY1SkFtEg4H3K4nXaPIuZW+jntcjf1b1Y8NnFqBnzpOu5D8
zQ4uqf9ITjCqtyv0YnIVALPCVonyUGnpKdCGMeSYjtDG5naz3WR3/f5AGHv2JKq2
9LW9U2daTV/id8CE+fSJmwl43frVhQ9Ks9IiNQd2vhzJ8rMJHyvb4p0L8/lH2UGE
hCzEgg/8uMsU33lmjdJrjq991cuxdAbtaYE4GuehSObXreXHzPaMrvzWpjuv8m6k
9K6R6yVH7NXF14VDW26epzlO5BYqCUeZhqk4taSrX4Kt+rgY1w7jqbpVrhBPbiCK
/jxXICsPKq9GFbPEJCDqCBAjpBHv7WFOlzcJaEak9oIAj2qWftg7BiIs+xCBlMdo
Q2fMTZzye6HTQYd7oE57t1vI7JcLTKJf1RMCe4bZD0OLIRhjLmo245G4VcYA4Uwk
A0xezzpLK9qokoKBkhC3ClFDhiSRhc5Y9IoVLvbakQ4AsIydg9DaTJtl+62alN8p
+3L+z85fyWkPy3lh8ftF1WA5otmpjw/E/Nyrrrz+gUYy1oIlvzYnV5RfFy689dIq
CE1f+wK51QyuYPxIaklbqw7Jghy3UopBvlXWmG7EwG6oVE16QCCF3gdHB5/A11JD
5XxzEGKvPSvlIYezMcg9+jC+fTLqs+qe/ztd8I/I4xRomaCMKMzsNBxMAZuZvs1L
FQ9j/N+gD4aHbjc/maw9DMLUBNS5Fo/A+CJ/V4oF5rJgwwOLw0b4B4g0h9JQ/ZA3
7v/HLIxHtvngZaRYg3juqhnnog8Bro3ZNJwBfJTO1iRwoe+xNfdDI7VAzooviVU9
EsBzSCo8Z75S9lx80C5LXcpeLC0kBD7A6jiYA64BYyONdppACrg53H5YiKM0c5vF
Yn4ZUAJxnn4kPq0+A7UUWD97KhCtueDU494QIJQ7aV/fQJhwq2EmmLV2XucBRcN6
UgedwppOYXBANIi06gh0okt1WbEgOSsyxDfVW25TebAsgSmcgxeuQlybCsVQBZSr
XLAHu8vKhpyyF6wsBs87jx2WdKKjEpnc3XAYVrDcnqx2QYa98xd9c0LKo+4Am16I
xGwgW1HJaIC2C7unFSwRL+xFIuWzVnTJ5wIwkw984zvxGFbcJRXkDOdgSbdtRhvT
B+Gw6l3CpPIqKYHX+NpxYF9g9LxbN7WZQliydBCI4Fovbx/5c85zCubXezpJpYN7
DBtteUW1+8R3PeWWUcGPmd6GnN42FRBpkeVomLoUdVkjS1lySyqtF0eWFo9gghO6
u03D/Q/GKVyLxuUgnmbSyKgOtclqAt0YZuslxqz+KXs=
`protect END_PROTECTED
