`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbdpIqjFjb/0DGsb8OjejCVvX2kcud1W2wfOGbs/DCLDFEHQRvoHijpp5zHpjduC
bSwHcSrLEGMajbnseExfzjkbND5AhtHNZbVJEv1cdJnMOYFom5NzYq8J14SCo0xn
sRu2EC4HGwwTeWswLbzsOEahsPDIKFCnhyXIrNYNNVcboWW343+rCDTC+mMNLeHx
xiaqsklC7tEttPQDxJKVHL7Dn3UlmIy42Kks2ITB+1JDSkVvaur9KgU+TlKt51p+
e+i/tJh3MEjrwsDjwuLR+lDHdS5tdJLZqzU+tDhPtdR7uTySTeftmcq2g5oYbvd0
nR9/Xm24lYLfKSsQP8xNZpO9V28YqC5NQ/nuqbgquUVay0Ez/DjfHiV17SawhMdC
y2PvdHynJfP8Mi6vZ3OkFCOV/77ec7jPa3iSoL4TAOmEFgz2wFk6PQ1XVdj5YI8f
jyz5GtS9y/eELNU3meo9Y42fwum8OpXXS9MYL+e3QtQzbJtxGrPT6pmmZtTNdRoh
8NZpFvfFeihD5MPzOrzHRm4w+el01Nbrz0ep9df6WHzt6A1glkQAb9psJkS7c2IM
U/vDKBscty7U9pSceoFLaMLTCcjbH/wWSp8tL7Y7GNiqdXbAs05tVP1/X7pDy5nv
foRg6TKmSsOarto5SeJwgGMA76m9hedFlc55upYXgz6ynp94nlc2Sxk2rBDTGfDb
hPZXif9LO4FB5BY4una5SraEup44eSW0l9/qUTWw/iwdGC6WbtxzA8aBwcuMjzc2
a3uoK937jIDvZC+qXyT1FTP5O2iSB1Jjj8kn8a/ZdAzp3i9DTviolxTLm+9uQmvq
F6b8tPDiMCIGr6H8+AfOALJWIUj042oTslWo5UXLa0M5D6/sUZ07JbzA/KwY/lY4
44XgqX/aPCm8VQRVkRPlH8dY2PKLPzf1GrGrzLyF5yX/ZAzfn+wYR6yo/lQq2My0
cXAgh4Yt8/P+JrubZ/ewBAT76oHeMPRPdV23idmxzoaL3IBndUfRpyYOM1SKikND
iCs1DRemOiJi0c3fSPZzVP2DmzeImSOylf4mx1/v26knPT8AcN0f6d1HeZKaeZJv
+GjsCW9l3EOSyFXR6qhscA==
`protect END_PROTECTED
