`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxuMi6mLOoYOamhB/3r1XYu5V8pmW74mPKNalNNu23hngG/rGRB3G0OecMuaVdlR
kvoSjLNR1OZH0Q72MJbBm0CgJtrOELE4RVsLYJKX/yVOJyUj40/bf+PuksyCgtPe
6gb4oSH94oVwp/JXCb7r8CJZGdlfu1XT4lCfY8J05Lg1P2v2gAokS1yfwTUwfV5A
LjN0d1wrfQhGx+ZiZbGSKd/IIe1yOQcxSZmlT01CNrqb7Pn/3csHhXVYPZocyoE3
+cQ/2+wUbzc0CQRivX67AjM1QSV1hj04hZKT95C5oCH7dkdYV/JBhaIOsqeNQVIK
WCSdaovdZyeWn6YsVXxNSiQqeCzyTuESGOZ2Y8vWMh92W0xfV8RiOsOgS5ZD6sP8
7MbyTE3Pxem9LfCcoXcNMNdwLnsfgHIGiBLczilR0GDFJQup0Nz3MFPlLNSYXEmz
9lyMEygJzv4MjZwKjUK9ED/QlqwWHR0Gqy9v9PEGw1bPH8U5d24rmE6clqB6NQMF
j9C4ZNCfJ70Li7Pf8IUb4sUgcBtJbmxED5zg4ET49ia2+QNtKG/wZEpw6xSXny65
PqpitdRclTuvuHPOvYJSJ6YBynZ6GBTOQO44caQ0HT317ZSREvEv8LJJ9Du1s22B
lJ20oiI7YTRZbIMk7Ndih90BawW6WRdhVHIj33UdniV6XSqiGEib7cST+UZ9MksC
PhNlcW6i8UKywNH0hN1YnsJKvWBjEfFxAPnkEFQQ7RzmIOUH6u3ih/irZjLl78k3
QPtMIscraXuKma0LwNEZkmx9dJzev+hPTbVIj1KXtiQFYVd/4ezkD2SEFFkxXQg+
rRr/MjZTiXMl/UW27N7RaWUbVCYImWk9O50liJVPh2Jjns9hVZEvfEI7VW/zstrR
gSFp0RdhLqyLtxXBiCxqs6nXZ7OWMIbleJFBu4CDjAz7yW637QysdaI+iqF4An4W
V+68EYQv5ZT0ZHY5Fjjmdos4Gmw5Jyer8qbuFZqRynz6chsbAoqp6+dGKhWjTIZT
llMZGwPei7+tODFpnfbp2qkILvaVzjPxzFl1cP0rgSuZUZnRMCHAnlC78M0y/oYv
mLnWh+7UP3CBm3sftsDW7Ln71hNjzQ+vNur3sSQQAd4=
`protect END_PROTECTED
