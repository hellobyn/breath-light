`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aRtcjC1EkYKYniYGLt8frsFlh/4K+zwLhrar3Kh9Pq3jUGJw5kjJ7MRyqrdkKWpV
spp00nh06ajqosXmigSCpqJgYr2hQKIuQxvQGv/ZT4uwjjQ0qqI4Nz+Lh3BfvhGo
tKfoJOFImqb+qt1PZU3maxNQRol+QbESv/i/UPrfch5IDMGVu0zew1UH8cwaGlsH
tBmFYGlzg9dhI7G7oKCLWPVxZwgWZVcipgA6cuF+M8byTdS0J484rkpEsI9ftjg1
yV1b7k2i0SoG1t6V8pN8CdrtIo8GRCZXkPA9W5bdYH3UNLWlUbjqKp7mzq4PZmv8
kTDKjsp+lCcRaIJFRdvrys57TAQN1HpZBuJXb9SWLY4Bvzg0i/zqmQ8jdzoZzNLN
n/hXursMDa+Z49yjuSxwo5XoRU2bRExEX7f83ry219t9OL/LlIWOq3sCJon5Danv
04Jrb1lDg19MwN4cgGyRvebaa7sVtYdJZ26sioYJ0RtmRSXnHDjc7qGJarYA+ilX
poCgtjtqTkobqzwgj4z9RCwi+t9dBl/9HqhLA+blmirFszP2ZfY5FPU+lUdrAjj3
+zvTYpPB1GrNjIofODxOgqmpzbCv4U0shGVeEAG79/grKDFyNKkVMOsHpXYWfgDC
ul5u2hn2Qz8ptqLiptd4dtOqwzqc5MiL6dMxX4/wr9nSfKwdzw//nTRyUOydWIyk
0zHRQW16cE+0AQCYad5maQ2bJtbPzz2wfccToHhH5XEwrY072k509VofwPkM9lVt
C1T3pQENcQuhRolbMCdWftRZdpweeLwDGysaXms2nqmQTWqBX+lT/dVn8YKjG7ml
dUp9YCjueBXPiBgEnqSms8PZ+UrmC+U6a/vFbsc/0Gkz3RYNOjYRnbH8NqiNNFnw
dB8CVo3iwHrx8K78lB+AlcIsxF/3WXJWi/VMa/tpQ/o=
`protect END_PROTECTED
