`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UV+t7+T2+5M3o1fXpbJSNv6BlMrSif3+t+M9TxrExBe1GK4jCRahwuk/R/Q1txyz
U1QvGuTfZVftKiWIbq+low4I4xnbZQFDf/Yo1D2V52OWe4cwKfmlEvYcBg5QIwmu
3s/mmAMFnyifAsg1A9x8Ozqh8q23ZbwdHpQhJD4HyTM5IjabMEMH+uzCFvDk89VS
oPBoKjJYK9wIt8GEBDdku1G4WXF/wcrRSEwQFY6j5OsoLA1osXo09Pn2BYE4yFRo
wXGrFx+IrEvg8wr37S7Up4VBFcFMMPBAqJZ6+sBhSDieiCh5b/o3Qe5E+FVdwGH+
5CFZ9QE/UwCMJwU4F5OU9fQoW2xCDshwlKJGlbqhVdsDRTNRepkUDoPEoLxf83Pb
QxqU+emkysZSCFL+tKsuKlTmYICP4YCHrpWH5UYirfD4MaSLZy7icCayW5oA7mXS
9wR5NE01yRoIUHnUpOLVc3PsrNWPjpBzNJF0CrAqxsghCEDAiKYiIVRSrk5QtxuS
oaRpIl4UR72thglW8mOOb11J9UHJ0VOEErh/0RbPww0w3FvFcvQUFWWs1uavZrFW
3K2ApkXJVDuqCGyU33ed1xoQL4ioe5rctpoxdkJ40jlVJCC2aG4/MTAIel4nEgoX
CaxsEm/ys7XXgPvQDMcQZakzd22Utmp4mURf8WRko1L0qWXKYtb0LSrMy8qgTucv
+6tQuEbaz/O+LbxAmSnW5FTpLaH8LxX4zMmKVpekOWcIwiqVZACTnPJVENs/KVO5
2V8nAXTqSg+9/j8SsrK0N9siEU+Ree/nrlzWZEh8g3hdCM5ni5fpgLd+SRyBBt+A
BRPd8ZKCxbm/kqYgq0sU4VDaIexlA1UxoZeWL8E4SZW4esJ4P3/WtDTgHxxFSyjm
Ds5z9h5K+v21az4DamqE2JTgb85kWYU4ixqiWdU5AjHI5Lwl58PKCo5lkfX4yb7h
6GTlSL16ciu/+HWrehXF+K46TQNuiJhoXLX1znQPj0k=
`protect END_PROTECTED
