`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkAOtkEZLMYvA9ui5zwhIaWiRNVAJMz8hgLo00Mmcob7K2FqAobbBxUf8n6+5b1v
Tz4sBiYF34V6TSfnX3/ZDiKrUhk34wANgYul6SZGGHLa/hNivgKgU7baToTKt6PF
GekKjRzL0ovIsggxfrNEbZQZ6aSPVhSSeLg+fgONZReT7d19ca79C82ynWqcDq+M
WQTcyxH13KOz2its4cIvYdoX5ID4IScblPKJN8o+q/QwOh4tgyRixsjXy4J1nvoR
+WrI2BTwZs5TSuockr6X8+8LReGd+zIH4hLFEo8i4CeJAMOBSwSMTN7gIp3dibVa
7r7FFLM+K+PKkG1OxA4qde9EXoxyMARp/Bf0JNtZ7FY4mLN3i4JFP/5fb2jblQHl
0iktbOqpqRQgYnGcErYGH4bx+j4kTN7jQpOdXwa+S1i20abw8wc1lEsFqgzBXWDj
EoL/6JBKA0BsvxdJQRcoPvtR3Vc/LfvWTfkBOQZcTImFEbAoXMDFjPW77cej0oBL
kskfqH0gGeqiImgWlg/Wnz11SQLwnbSwc3mAaIreEeRszigY/CbHswfcpfaF3vG+
/6rvmEKAbGdFVGVxU9wwYueu2HA4ea7Xkln2Rq6Bfsop/aQu/tHAR3LCqVMR/0fm
jn44p7law+utZe3+0mfVYuXHpl1Z5yPSaUc9zad2Zx58EcMa1/adbbkkKii+B/fc
xY18yvqAku5WI6APwQqUdCKCPj4eif8zfJr/T+XHGtUCnKrINHaWHgU35i43dT7u
954RXPwsoE/zmXMOjatMHndphUsBsN1d+iZsxvloINKAQfx4S5ju4elcTmV6EGxb
pvqMaN8g8Jctes9RzBuqACf1bKwGbfjmQuqb+U/aCBxQ0jQoqRUH0wOQ2/asFtZv
CRzlaDK2nNBEi5tOKdz81EmijDFoizyBBufneiXmPAQB6XeyqXFXhjls7uxyGfRk
KV86mHupwR4Jg0Oe/1R2SlZu41IFBar+AefmBMWQoWsaTBbgHOEdRKyLqTXNmcBX
k7ebdi37olD6JadYglSgA6kEtY5tkI0eGAxi7M/UXcSW/dnO+9Ylqs5mDnNs0qVR
fiuO8X3e4HWrF/YcMbmpJ5Lrmjkf5s/oWx20v52JED1eGqHUu9Pmkq/zfOLZBxGC
NjKevl2Jo+pvQt/tUuwRlE4SB1JV4z2EeYuOP1b0n84W6xDIicJdLWuG08GDIc7A
Jt+Z/mY3x7klKucMFmz1aQpoN9ighV8nQ4Wo+e4C9m8f9ZQQ+GVE2oyBeYvBS7A7
`protect END_PROTECTED
