`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtHlj2cpprh5Pzy+5vXs+XS9VrjkpPzBJcylBuqZppYHZT4QmJUBOMatk5Dji4OR
8+IO6syZSqu+r6KjAb7JuKjHEwDqfq8n1Wc+VHok8UuG0B8UfB2+weUYdmX9N97E
7/RwNmsrpXNF8g4jR98wmAnQRaVaOWks16SAuP2Vs2c9GTMjR51UuR59W+vkkLXi
UcW8lbzOBVfFFZCNGYAizricsmV/YktSLiDm55GpEY3aJv2tcphJ9XoHnm/FvAA1
JVrQ08ahMtLTJgWqH9BSzMOxf6FRBPHHMenp05uaPbGG+auvGgxqH9SCsYX4zPNe
VvDi2ygbHBXgdAjguLf2lojjdR/dLLwZgt8ZzuDdu3BZpCwkqKrfuR3Yzj8fPBqh
RvT7PD1YmAhjYKLecQ/pjjMqZCyDLZLjuVWLXiiw7wZYpYGLL/sZEmLhhkStD0Uq
UgREi3PWCdaxNZe2zggz3gxQxoSN2mA3ISx/Usnr4WgvDqIWzuIEXhuwNBtoOV22
1YiMZY6bdrya2RYB+sDclygX1Finj0QPJ6edzesxi19zk4XteOk9sYKUihotet7e
a4HmkOJbvsyuuelPIcSFDx++Beoxyhv62myfUOq8y/qBfNvY/OpxBn/7AE3uU3b2
YIWWGOU4fgqeEbUvkmd2P8rFqtaUgUBGkA5Bki/EXsGIvaYDqQRi3nQbChX8PH3E
IR4MpFElkcj4VIHVU6KYqF0+sjAN9qBW5ZzBZMebswWM6dhwrf9ArCo/3Y/6B2h8
vvPephPZGvAgA3I2M7bVZWyr/RExxYvFLooZWp6nnINbgvYbQ8z6Xi0YawAY79mH
JnmmGE9ufEHcr4tbrzi1FwpNdZYJSrokkFp3mPv+ObkqjUFabxh4CYFxj/aZSi5X
HJ3upecCDCN4hKgHRBk2VCRdQbbi3a2UyP8cf+Z79R8Jmw4TeHy69ywHn9N4+mmW
MX/UmA/INYrclRzlN+RQldbpo2xl7ddsnY1/szL7yhRLPy1rff0V8ER06Vc6UGQP
i+TpRUM9OU/mzbs4L7KDNQllHdy93pc9j76pgv5uPDb+FN4DQ5gr/kVESqnMlv4b
/BujHW0T38JcJtTIaCJIZdGMupkR7ZI7Z9hZWEr/53AYfwoYiFTlYztmeMke7a5r
REznA733oDW0jivMDG2hklVmmr9pFgD9Obui+ZECM5r/HeJjO9yASmfK44lR35rl
fYe6ihUqIrlCgUcoGHlDuqpBTZ5rzxsfLK4bqTdB0vwCffhZecBkwyKKOEQOEssm
R+ihtNglOqxpyQrIq+RTlS5GisSAkvDqxiKV6tR5jhi1IVv+AFJi1X6rQt9zngwr
47lfOhi5Yo+TC6wVENB98+01gUqC0JcReBDFq6ELifAVRwX1g8E2Byu3i56bdEze
frWl4e1Jku+pWJtFY+LaVnVIvSjK2ITgYUU/WCR6DVBhBm8DDHIKdy0Z5NfkNFoh
h3+BS/BUTBJmCsQvGeu3PPTSfLuWbLWm2yqj0Cip9aVgVKMWs5UJBUHtq1/Zl5Tw
RGvA4fWCTGxWNRijnW2QTB8xnT4F3ZSadnEv3Ip82cF2HX9zQGX6p3qX0NCJeFhK
a61FZpmRwx3E2Lo/LRx+pffyy/QIx4CjOKM7cruWTN8bckmXuS5CaVXAv1heRhhj
SXGbNIkQjv1WFRpxsVR6S0IJc8C4iPa2Ah3M1Y7HEIrwvxO4HhY1ojC8IpCBubgL
aSnF9RN033n9two1KoNo/l+862RKMFZg9++yhcUnXxQE4UsW/51M5eVIAz8LRW/s
6aYYlnvoKqy0OGOVnQcTzhTxGVRJ5KFp53DRltgTc5uuyVMHAL/s39Jhtc1reFP1
C2NUQjXXfdf8CR6n4Qm3lRwqN3GnKlP0bNIf54S3vcgYjFcXRvqqLsNeiInnTNqB
u61QiWDQN7V9HPWWxihOsUoEs+EuI1KCU36QTjh1ZaezWVFmSjgUs/XhL1PJ65qQ
gO+wXNi3V1aMowYiu/02WSUPjOXJbdwMd4/sZIqoU0Ntp39ghH9iMEmAAjDoQleF
xlx8yAbWVivK8SpKWlxHGROsunLlO+9FA7G20G8esULHKvDgvVffWBWFXINLYvXi
UZuk8YY13hzRd4RQx8VbLwv9iRSTSa+9vkInBK4iSOSrd5oclcl9aHRnY+rjwJ11
HCo4bFYAwfwtT0W6XsB+aZHwJVChDNkwrQW6jePcOD7kLJ3kOWAJU34bBzp4yDfp
hQ2ExGhLX6aGP06GqfOQIKcZ58t15O/bpVWBJra6agwnQlFLzdZ0gYNDLqlvE3N1
A6WtWBbuY0UYnisI76kg1B5mai0NvyGgeTNd1MB+qpVL7EqHvm8EUDThuaQJlx+Y
QQV+4erPvS8GAn7tOs21LiT9TvjczI367x+YhV/ggmqKc4OoG766T6ynQtj+TP2R
dPdTHI0Yzo8a7dIwyBLtfYSUA0rZjeb85/zWezKc/zZVr+ir0awWgmxwsj1eQR+a
9TFr+eruxlOCBRtW2gl7yATuxjcR0SyDDreG8wdrZIXd2YFTiUi3ZNiwWJrHToFS
iXmhHWSCRW85rtErZd+aENIKErbK63D7DSmBvIVJizE5CRyA0G7squrMlbhKtYJp
R9zVlY/Ty8hwc4NZAdh3JfYNFl9n4xO4f6ylHTQ3ZPtEkYq0TPZXAzotTT4r7ToI
A47toOERtzzybqmVLCtWFQYhoHPHheHF9r35to5O6kT9J+FmG/x0s6NfB0IlSa6g
Vrhh6QMxrxAYZyGCU9Vg/d1QD9KstsW8cUXTK5DTvPuu7RAOIEwAWmmhEZz2xShi
bnlXe9UJw9/dgLGFpL5axY6zvo9j7Mw1S0/fN7hwMEx9HKYiHDsLBlt2PPtyUTwl
IKaHwJj/ApfUVCHJ0AbyK+BGgMeZKy9ozT6pI/5Vmw4Ap+Qryq9G5xQEGdqMV6zZ
sFL3HKiX/dSpEds99Fw0PwiGHRVuTFFkyNFjdaPd8us95dFBKLznVrovrBlfWqSY
xube4xZbYQBHg+K72zGSbCBPVZDex6m9fVjexqaJGOhm8Z1lSmlLD71ADpgPLidV
PakODJa4yKF625ER2G8e6wCsk2UgEX9IS/c84dB/9AvVmdCw56AAE996lxL0rYVK
X3gLT/lV0PGzWYG32Ur/WpTVBMurKMGJzoEUaiHn9+fxfhOV+lE+wq9PdeOOy7Cl
veC9B4IgHkCuB9RECPlei7exyllKAI9A31ivK6QPzq4pPrcJbxrSy6vzXWMYULA5
pCsx1EYUtun3m/sZhF+7F/7Uz8EJa5AiG4/7U25DHrzavVLGp0m4QQ6UdNlSEM/a
C+F3hM75HQFX9zf9FPBdbcCrjvqDvuyR1fxrKbPbcefEdfW/hKuVM0i54yBd5/pq
ce9SVHnCnHHJCHUk7wSn0RqaWTBkcYXAqI9PX472z9iA+U6L5mRtmheri+v4d37x
P14y5AQioS1HgPuRAOMp4RJ2CSQC/Mh/24zpTrL9mlLBFQbmc5ghNO9EdD8NfqHl
SO/lmPiez8lVykiBKsJ6kwXut/RW16o7FnPmQvjWW47x3PrllBWbVbMhres48sa6
pC9L1CpiRiExgHInhS1YTVut8YMkRCwy/QVv9SVuQsoy/DHhipJPR2e4oPvkZp1z
/kdfrVQS6VvfljRVvRiKWLB7LpIzBT8AXugwsjO1/BNsg3ZtdCYiNDgKFJPVgrm4
J6l3rzohGmVr4+eeRA8y7KAn8dWxR8+GPazME1mHzgDWgShy7Mq8NC57NOJD7D2l
jLTsugjiL405tWedTMJZ+3tngjqhUYphYeqws5+mCMWttBV8OQDEgVLlMKTXJegq
6kRNPmc7hUIkXcKsGKPdS5NAXrcqF1+QPwVDOSPRtxnhtsVG54bhJ3IC+4+gvzjT
yHX3Lhu/S6brzVD0u86CwBk4Sa90g0t4m0f8re4YSwzLbHn24vvfty2vCQjO5+jv
0DZL65AECxz82k25uftYl4Nh2eimP4mPnxQ6txUtcrxTp+kngTUjO1LSqYuSJSLw
bdEtu7W8zEmEE5GZdLfh411OqPDxe2ibmUI109sRx7j9DJiNmwrnnKQmiCoM/DjG
9LPDoCW3gvlLKvWumn47KSQe1yP3kZK9EHlG4PXBPmtOhfRk+KK1GMz+XabAbdgA
S1PABoF1T3YrcmuIK1mUsj/qzVBhoW+ik2mddv53lno6zptRw5icPQTCRnkOFL+p
En8NzpoeFm4zNg1GKDJpFFptvWg8zjeT8yErvQrApHgHNNHNeORWjFwUqQZ+FcPg
gcr+3DxViCCh6lN2FiJDcqJJ6nukJkhgfbw1Bh0QHJpBwjGsFIHZxngCKKh8LwiY
0TIDjvx3CDb7Cm7k6S+DwARR6pS+QjiOsEVzU93juTEvxe/TQunW4di46q89KCwJ
l6DisDTmc516i+S12L7MfIqUyPEG7zjXOTbvVdw0s2dI4HP8Z3YsjTUm2ZBJjnFh
dxE1fJ881/q8htSGttjLdi9lTC/ps/bnrCAPhJSClO5p3ziVowJkqigK+ZjNYF83
SqB355HSq/4u5fMhkHCMC6D5vwVf9IDzn2wCnMj/R+yvlbM+ROWWkFJOpoBvjPRO
lpJwKmfQq3ns2yKEPXNndp+oHK8pMR0RWzw/cH28+A2TwCVPEkiBRKODf+VFbDk6
h3TNHKCXCT0P2QB84cX+Rt/E+JK3yECRALXi+/Pt/BuXoQSqQcmlMUKVAncnN+fb
NxqeRteBWmZXs6BLZlANZuu/qYYN8LKb4rZVTmU5Rg4wpnq82Drp+Gj3vuBlqcMr
NVFhx6SZlAolTOXNnuyg2LU5F4V/f1o+G+A2Bl55ygEcQJYA8+R/IEJtbtnG+1x5
C+8pSWxDXmNaDTw1GBC8OdS+wOSJcY18GLqg9ejMRZlBgSFNugqCtItrCm8YPljH
ThtfDG4BcH9mrCt5Jv+ezBVzBpd32iVJ1emSOYW6yjBy1s8rXALV9uPvAN2y5jVp
TneiX7GZ+0FCJgYP7BDO+8enJLhINYYko9Uov6ixbVvXUdK4/kwz5D5ujty6hZZ8
cTayNDmEroGryIKwYX1XowmFp5kWToCEv0nvcgDIzTKiXKIGMf9pm/P4T6bIeMxe
HaLsZV9ig6PGJQjY00rmT4dIy1u9bzecGG5XT43xO/F635mn8+02RloS8NpRgzqC
LzTs4DRCphWQp63Yfk/FNGPqGotqVoFntt9ZoIFAY/MpiJOmo2bv6ybU0+tKQvs0
/EwtRPiNnslj6RnOlnWSqxmubhHwy2+n6S/cT1F8KHoQ7vIrHuZWSR6IV4dOqT4/
R9lLjn8gMXpx20PrAuOxEPXmOT2q1mDyS4Sfilc5oYJsMpkVcTFnJMQilrkXpDrn
WbNg/FPRgK3/o49Yr2LM+kUH0IB8BVgUBPoCvum90bkBgcXuXUcBXNzCZoqmmiz2
IZHdFAQt4y6kuuxEeO32Vjhra3e42I7mNBCVQEuBzJQft1arQQ1j6+45Btjx+03c
Z+3GGMP2QWy/IHHr3fpvwJt5f1Ht78Igru/20UiU12f+C/fR05K4njoeKCj8GSrJ
HUQO/8PiILxfDaVwqY6HjHDIVs+Mj3HJQjv8XDqOmDMOXykdVYgYLjwWdBldvfIm
mtGz9Zu/+b7vHI3ixz5YdlNBCFML01yUnKiqrKg5D/g8TMlcx9WiEmRcn7h67Vha
w8TK+TLUxKocc13Fr0naO8IrtDzRJYisgo/KKEijWyxYmkwj2mDv0lyajwq8fDP3
IXyg9KQH9FmUBjV8qHekwZFAchbuH/zPi6i78IjTEG0soTUoscC7gRK4eyAui8qT
BPAMbeMR0Dntwesn2Zi/ODHb8wNkkOZCyOoum6gqLKEFuDJjKNiRFKLGrywNvYc9
yl5PxEeFba7ATCAijemO7ZNzVXH8yC3Y5MCCHKMvCG72tw6FrkjqZclkB/EB77ux
9eqi4RKag4u6aw9emrOIz5m7jue//2JlxWZu9ycuR+cwI818QqHhbwg/Bw0Iamoh
FSiaDNDRvVaizJT/tXU1YP8i72zrD8AkeFSpEeB+CtUiYtLqUEnPuwlEXai/iicd
F7e4bXUvV8kotQql4c1XCixeWCjntZy69ylqmT5vzpjyfvSbJlAiyzNVrABYPEo/
XDs2MLgC35Rr7Csx1RGq5vPPzt352dT9uGXz1nvpWsUj+FDOiBIRQYpVNUfEN4lo
X08cpJU4ySQp3Lff3lfh8PUZ2jmL/enPbh0CuL54bgQInvvkCJIpbOd9Ha/onu0j
oUJcxh1qF9VlKNqd5Ppvj6oNco4iuKDuUj2zOXXIU3BIIdK80I2M7bwcaqJpqEkI
EkW5UYXtJCVjglvEUl+MsIywjHHtWwCKgPjxdeTw2KV4WvMasgqLpUHL1FA4sRJl
xAxmCTsfld9CvzjLvGTLQgm00Fl4vq9zmmSVhBy5vpjvf6cYGBycTAF8szm7kylG
cS3/if8/KWY+obpJl1g8VNOFHR8vzSR4bLOh4tdmOfkJwAld8qQmOLWJ/T/boywU
UWWHPlm/iHa2vLkuXd+hqdTDBT7+0Q2pSJcXA5xjhjC5r42jPWbqDMxdhcUPvzm7
AwRXArNgBaP8OwmmCJgdgKJc5V1z/BE7h/Ld+s417Lvqu6M/K+6hkOIqyEzR05vE
ZMOvTtzM3+2FR8rqLEbAjVDxH2fabH+mzqw09TLMb5inq8/ctdtR878y+AXVgNKu
fMQFkKepJoNH0wWMcBIAeOpcB/b8455QyCP4OS61pqpuGB2+27WTzkM1r0eQyFT6
btxuPPsWBInAXM70OeQqiLSM/sBiEOf/AA0EM2IncpNtQbjS0yrt4q3sQzMETc8r
1UhLC1tyw3VFMijSzDYFvWaKg4P3iuwfUZA45Nfpc2wIiP/sp4yp41bRCIV0RMnJ
cYaTam1BSV/P15/op6Qd5NcnuK3Y5WgdCGBBOij3TUV4HWvRbOPC4MxrQVgQqjit
o/6YXBzlm9yjY6ulF2QQB9CT9S4wmC+p1NrOscB8LYTUDjBgyKHdYpBu8FLN+0P7
QZ5spybPRHsTOLLSlAYGLlSZYBQzSy26XBsytVvvaKdS2Lgkpbll+/Zf84k929t5
PE49SqaMf4PiUFSLajOE7wv/p3uNHR1R1H0Ny5o9r+tPZNXJWX3ckWX1IqxXs0pR
cLWzRhkkSyJbF53vSEwMlrTZ6W4QdPlxQXtxFC9KQoZVWz++8wwWuz7MeFaWe/6w
FMdkVd2pQGba9Atbf0CnggASX0MBgJTXQIMaMEWSPrMQXjGVrK2LFYDxhSNLAbso
WvhwYqf97FED8lRFSeP+CpqYek08padG6mE/R+h6J+cyK1Sr9ZWxO2r1wQWOZ9Z0
xrNEZWuBT0QljRasVEZld5g35fqrPn61/zcmKBYtd5IlWtPpe3jCm10toWo16WLO
ZYq3Rx30YINSrMpDDIWybueZpgomgTAqliGLLfVnBrs0J8tqOM3jUz5ZyuCVdjXU
q6CnkLIQG7JCg5gzOLI5NsrKgV++jbNZOiafNUSEL4jbYpkb6KInf9D1T3Bj/L04
LPi197yAzv/pd+LfDUO87/L1GZ27k5znWggMgLsbANZunFrZFi9ZNNDaqXrNnyHW
tKB11Ed3nAWZRD1LM6YyyQ7G/0awOyrYSd8uu/JfBGLyMuz35nd+5kTBXceM7VOr
XZUvvW2SmfQl4g/lSh6L01ceMomAvUn37/6SAE1NgAwoz/3FsXnZBVR52Q+Ab70E
PJ95hI07kZB1CMA2ooclmCHcIb3oZbUxdpnmEHHHhvkkF1iJU1gU+nH9ldFtp5aV
763ztbuuMAgJb8u5GQEo18CVvfTZCe7yoagX59rNDwFtkP6HOZYqQAyHiwXDO9lV
vvxCQTsxZQQeeqAQe3spZk8hKvgwkMBxJRJX/Frwu65HXxsOxcxMbef6LcJMsvW7
c7J+8AzGlijBWMi4/9H/f6muNXK7HBV3R9p/73pS1IRaOVKNdMP/V6f2RrgFWfE9
A2LjEQnxqNJsdavIEKXyoGHBKpGuwbcIWM6aFZqeFksLzKRPFj+Clci0R27Wvcim
VhfdLE6XISIGIOaJofcNRgV8AvcMuCtOVqR9ohiivfndUpYH796lLqI8amHH9ICB
JYbk/twBxOOCYfnsUkZbczeAV9La5ZPPy+u/EpqgFchETluwmz+rx78HK0FhTJCF
x8RYci3aZ8YOBEDYwE5YAeDmurrryZ4YHdOipa3d9nj4lSxvPv2DUsX6OriSsm2J
zr2qwtVV0dotveG9vV09sKuUiV5hGYqq358H6/K1ICpwDm996RIK8+zNDKFZxjk9
1VzBYqiUaTLcfC7X/zxXs2/+qvg5sGtA8NXC3UpTRuV/vW4Ybom6zM3lIWO8fUeh
rc1KPicKcfTBveM7keM75Ix3ZQFi6h/688LiprARPEy4B61OlLgSojR4jbjLi8wa
ITkr6DEF/aywu1myO/zqRPYWW6Zez694K321/NOGiAZt+qlwYYZypXVPb2xhA/sA
42TnQHHoHM5SqVcwXxbPZ2ojDzv+xMHUW7uz1ETy1nDRGkp9gtlQzMK61yI9RyfR
3VPnIb6U6KBEokOX4wxC05y7KCfm6g5OxruEFClNmRn3e6Hu0PkGJVchqBOQvSbU
e4b8Aq4oXwFXgV0NG+xevbuYxuwSYEMEQcbWSYa8Lj4J+Kq8mW/cb3esqDWmfnhJ
2kx9qkOOTsST2J4rihqZhzEucss3eSbKPscucCcpOEW3gBDKznxqD01hlh1NKVwn
cmaXdN4TwhRNK8qOIi/A0Xr/dy1jmVsek2tsCt0GJ0DiSm9GNw0+n47n7/lZhSHW
2hcsmuL+6xSY2ApEBf8DYWVJcxPJPxKmf6WxM9SaH+nLYI3hc6BF4Sj8p50vijFU
xeoiifZpHXwcMWUum0rc3JgBtdA6UUR2PGfySyt7lvccokE3zagSD8SGiuU6upvb
q2AMf8jfvudpXVGOqFdicM9ViO6JPskfS84KiqE0F+3nX6fAdG7LvVaWqXAMip9y
3UEHWSxt98S7qaajHyItDfjTPcqpWRDc9dMCHMmcr7AoVuqFuS8Unab7moIkKku+
6h7rq+avSlZ9ut3yywMmvVprilipnjl4UMP3K4AKEdCcksQETXBLC8whL0IH3Htr
BGWdlPgVWEuO7DAMVrmho3gzLJzRNvX+qoCVIfPOb+Lhv0d8QGf0FqjjweFe4Da2
CXLv7J/FXT8tmsQXCl6PkUzPK5HZbE+XYvC5RMSLvSjRVmsvmNW13sbZPazj89M4
XOa6RSuuBkUIK/5zj053C+83R+pKLKo0v46K5RKFHIcbXS0Mxpv7xh7j8KC1Pu+2
sKHwwiMliyZV3m7P4xQMOSPvbiWKnnaBVtVs5bJ/rRoCRya0pkU/JYINMMb3Ufmo
bvvWFqjU38hR8I145QIGT7ySC+Iq9r7FjS2cNABCDLvK6S9ZeKOkkJurExKMG0Vj
c5zIUpNXoKllGD8v2K5E/rla+ijqk5MA3uLGkZW4SbcwlDTv3KaA8xNnE7mlr97a
qLQAL8ZYPE79u+b5/X2ed++hzOlP25BNh3oeK8aZyhutybjZL66627tHEGhRQeop
EtlbGJk0I8pIWbloeSK/ZNVAAslCENiAo9QTi2d2LD7bl+dN5LkyWGpsBlSJ3IPx
MMcMn34mbJ4BVmC6k++IUHANVFV8nzmUxQ2XPyc7fad4R0XccdBJVPReY05uDh/T
U43mPqeA/SV59qg/I8HEKH2mWunzMvEFW336KdL+Yr6y2hIxOmSA9IbiLqMLNviz
PC7R3mBOYRl6MotjGs/EaVoLWYvnc6uj6UrYq0qRXCClsr9WY9GdPXRz0G2+e1WQ
d6S6ndW2Ry3beeOLGOFxh9/nGmm5Kj1OSG/Msz+wktzPhMbvXrb7k8wa9XGE52jD
iUJqtgqWbV1tKiLFtl6CeX8qqYDdptHKEydOZgaCt6kuaMbacAKR7afZ5wA2zLM5
aZHquwwU+eMZ27mXWuEHzA5egv5aE3xhs2oPJHUY4XChpWim4NEEzuf8MDZXfBxp
BCp8OWqi1BE3Z4m9Pilll7s5I8u01glHoqYgnj9wrtqxmPv0z5x7Wyo1+9RFxGu+
Fy4ixF9nyFZ5kdolQT6p5g411ky6CWDnm6+AkDV7smWApUnBUwA2wRXE4aB5qLyQ
QzLRRpjO7LL+E0/1tFFAzebKfDg9t+EEoh1Xqcwm3tGrna/qeYPD8xxuO2FyQK2V
jjFbkoHEUAfk7GGrLUEn83TeP/j+Oru9Qqo5eM2Ucz75M8jCBgqYWrowkeAoHM2p
cFu/DpEycp+OPCoImYhleE1jPCK8K2h/q/WN3n0z73B3TKcwbrsJ7NAneTQnRQ9h
Vcke/8fkgFk9R8i4GEjBAa5D48SVJpSw4NUNPHd8goN5YZ393DRYeInvkWw8Yn2V
XjQvbiVYwGpNTVLO/puCxo/Wgoc8QeL5pZ0gmNxvWfPq3nLM6cdgSTHXgbQhUWkM
OhGp7hearzSbYcUB2wz33H9jz+6SlAC/0Yx+SyGYxhrYtMcT9FbcGxQAVtY/x2VP
L8WpAogel4iGpes4vakZsJIIfSv6gsY+ntlLdeAuQYAZjB+8nPCjXneOp+Zc7OaQ
T0B4lPP2M1CvdRcsAvbEDCgWL4735RJYjlqFt63lgEcE4Ce4tuACre6NGLOpo0V/
RpVT40Z/8OaC+urClXzUnDMKPXvXNy5+D78i89M2hz6iYg3hoiFNUeh+4/6pmjgm
7TlmdHKo+13z5Nq75HsiBOcAES3qEGPpRX7/GpeU3PQe+k+5CcpQ0IUI5Wx7dRfI
0m/rgZUEe6exxeyl9EAAuHtsSkuyOgukpv/0FnPKvFCIvUHtHECs3vcKBHNOruUa
UbY7tfhowe2UwN+kndEpsWDko4omsRGsQUBaHk+vhy3vVtYCuonKRTjz0pHUyGVt
SNWE7lc5KosEZ/9NZycK+IBRCnTya8hiR01Ch/32ZELKC8AhcPDRMj3fRGiKVOut
IIOI0GfrfJzsQu7ZwpXATsUmFViMHQ1j1mwOIJ4RnA7eUntzChuCjDXjIuhdzLOn
uPmXQEZMwLF41i5oH9GA57PpOA//DO/WtxEDBRR7rkjrTPfIUGCIvXaxUmQn/bVs
1TNjRyR9rG8a5UrOliqLcnhr009l3jSXyZeVXZquZe6q6pBPvLUs60XGYTCDYIQw
H2JS2WH+GdZ8G5r7+HyQZXK7VJxT84I8crzA+99e3Rwlh4W9mBI//f/7JFq44Gar
gQ3Ho8GxtQi4XBhVvJSnH7Xs9eRGF2RgYJDE9oaSm2AbE6Rabaa+EQwEWU0hpkMY
501Jag6wDaPCYtnlyb4lqRXCzbGe8YZNGzS27Ia0V7Vnt/LC+RKabswVJw08lza3
4bx5R13+c5v0z0mA+/cnYpG3+BYdTsOsbmnYVPxMxtGnrs/UyuZaOsx81yUV76vk
ULzBtngMpSTFuV8Ml7FV0nAiUFsmTR4miNjd0vfMPzkfiUGzgccm7ABEF4QOLDwc
z3l1xzTiEKtiMwG2UzABneKWCLSJLf4hT7IdQwSadMN/8vu5w96FI7COsrB2ruBs
3Of19+KOw3bhJpoAgqnqs2NB1ZFubBXFiV74pZbnFOVOyQJJLRD49l3PmqCFZ1lF
pf/j6UvIfz7NhOXF+mH34JO3+moiTJqTBIrZppr6bthzqEbdDzqCXPDQTqqbWJ7w
/9TRaf1RdKFQvrAixrjQccaAHpAYm6KHTSL4AC7CqA4hd8b+IDvtil/MpXP1wZmB
iQejFdZHXfMr2zNuF04L5mB0mJ0U25Rb6ul9JQwbT17QTGu+0j6aSV5k8+Ys4GNA
wG85mn+Tw8gN3oKbh00suqomtBsjLsfsinViY99DS48bB8KuE8/dhs3TTbUYVxMd
TaxqbweuVfutmfL2YQ2l86OwWt6vSbBfOLV0/mZI40AbwP6gQI9mQArf1CCSFqUG
KtdVezN9kV7VNqcwMdUYAdRZbon0GLFQEXu79iyQbSkaR8D9dcV10K6eBGRa3Bz2
MOaahYCv0hg1KSw2ttazrU9lT3HDZD14eLOxi/uov7eufTus+eCcXv9+uFdO/gxJ
bVyDCe8xbDlCkBzZ7Prqgj4VTZetb42Dty2A5ZUj14Jin4/TXIQ6I7Vz/CP8HFWj
PwcjwY2oPbUeEAZoCAo3hR1LzZ/W4dOaoeiRZbxjRRJ1YPNgD5FdxL9FtRZo1pze
XBlKy51rFDHSGGSHhJCCMdaE7ZqONb37GSCSkwHGZmTfHOBVQ8cgkGUExZzxDhS0
sXXqIPvI9TQ86vmN01f55FjcaS87Yo8Wf/0KcbUV0NrQ2SUAtz4uqf2FMiALh8/1
t7McbNhlaQYzaW8nxg5G7rYoH5/DGr+XnxXETycwJyIGqlXXv/q0re7h051EGga4
/e4eX+1fnEBurMpjKMZtKoGT0A0prlnWhZYcTB8iJGzuOEdfbm1AQjEgJXA+80xt
CHL2Jwwx0cIuuRu35f7bGwtmOGBFVWBW7EmpCN/ewknrWHXq9OyWoRtgwcZvZNOl
t5LM014TE1NVfO6lsl9QDPlvDvkqY8w+SZE6EDtDNCTrLvBOA8X/lk0+sy0YWW3Z
QwINvVhRVItZLT4/D9mFOKJNlayaTi31c2Zzy0pCjkkHuyNhQ0pAWiQDe9NVOe2l
o0WiEMLsnRMyMaBtxL9i39CoPPFNsEhpvHv6rY8SyYuMCfFuRlb3Euui2C1hrSf6
lzfISWHami/hYpK4CAgfi3LMcC+/d/4aA3XmayNojLghquGUeEHxdRgqZzzbeUk2
WmCrqOlUutiVyuHxXQT/b2np2uUxNjs6c9k9Fm1r1iXqkr20Nh0MTwCbSaCY5jOa
xNEAFVNcQDyodwX7tD2HbI4AtkmKamO7kHoLxK9s9PQADkdZjzlJBL09pAuqBn+D
8F+a7RNKp3LyCxa0iXLIyOHNwieLBOKizRRaZYvPsqmh9FgGvC4zraDM4ObjglOE
m7Ns6aqRAyFZQLl5K93WPWBLmp8ZVp62PGo4NWC2dldhw6z5CdvWl0UeekMgIzwz
M3KnuWag+wFLLZWh0aTg/7AOJk22q+9txzZAWMo+EFfl2KaW+5UzHx9WUsog2xDa
ZRXUDgzdfv1LzcD5eMbx5mQ7MZQu17nssFCQpXAXa/4lwGBf4RzPM+SlHDlvLTbI
p7l3revauSFbOUtQyNnJmi5aX4cj+43KQsKUsjnIp+kwqEhivXIBat53CZetNdlE
978yvmmD92Kh4JjggO7FaGjA/Wps+GZqkvG45sD15BSaLcWEcuYgLSA3WD9tu8C7
`protect END_PROTECTED
