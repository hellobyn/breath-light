`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qLf7F9xKF5Pmyi0P+sFu6h620xlAeUc1NchojINmKdeH6widBAs3+uWf6gOw1obf
xBTcBmfDcrO8ewu8hTVRoWZGMzyV+9PmqOPSfBYWmv888p0yaNEYV80Jz94lIqqH
CHhLO+75/XOE805HGUT7I8QWpNmCwqTC8bEmTpc4C2VzC2DirW/5ymUPeIWZ0i1K
vE9oWfCrt2cUwJ9Ksidt90x0GVEltEetMlh78rj24PgznGQHZiCkhnUbRq8XMhCY
Ef0y9gzcVt1c8Jl+RRHlMrhOH3JI+SVDu1/GPMMsbxjf3YCG58gzpzVHKG5yY1aG
14xf0P5I5QnbciVR47VlDaOdrvkmgorqLbsblPFuCTSy45CPgpiJPNBaBAsDvPAI
dgV8DAhHf+u/6Ojso3AR47HrknJ066UXOi5pEUY3jtskP2alYbHc052aCNp7usjN
LXrIrucSAP95hnwaCwsR3kTHziRhV09OiQzgLzlBMeuqwUQL1W8VnMKYMI4ttAGK
+KKr0yOm3scJzd7Q+CRBTUUhEIwEqZ+y+dF4s5OvVKoYzWebsgWaT6l0pz5rgulz
Q8qNPvGe7Tak0RrWz+5i3EYVUT3nFwITl299QbDD9iCMgmdBa8TZrCn0CUfSICMx
MaK7b318qG2DHISFf9ztz/K+jPMWwyH559Bn2HFToqxHbZiFXVvpNp8lfgwAZMv8
XUnOZCAQ6MyVtWgldwIWFXFkuLkDYT8CvsH9+Eiv6MsxzFqn7DcqvRlyGK9fzrg5
wD1/EAqYOs+f+xiCb9rrcAA+lY7EXD7zKSb/863C9LiRmRGJ2hzV6N86NJEJ9rf0
1V87G0F2alNjuAwF6ErPqfwJpA5mjimsvrnhcvUsKpWLfNsDWtnuOTdAQQ86tMDL
0AbzQ/C/hRIbeLL9PydDA9N30rhBRHM+zSozRd4pPv8jjqZvRhBAa84+DSYWG9GL
0XesgPaNyYonqNW1whwNQOwA0iDdfALj42LbocHbfSr7jo+ABeHjZqhitpO/P2Mi
KgpkqybmHqsyHfYzPCQg7M1tFLPERTCRnC8+WaoVijTFk3V+EWpfCADiUQIqb+6k
dl6RTT8bH6jH+uW+YopCEA5jLxyuiSZoSX2OB00+s8an7RFP96Xum6ldbztKwztw
cuJuuV0NoXlOOqF0uXazI2OF1VGEEPEPTlxIima9qjVsjG94cFaBLChhW4jBw4yr
jI5CygOlHjo9lxZXl969JIHvUsjIJ8Nx8BNSls0a9fwE/WVQmTpip/0X96hvP96A
IRJ0qZeefGZcZgNyAbkxE87Wk8cPvWFnBn3xUVn8QB5pPYTGto2vZVu1hx33De8B
S8EV7YCSu8Nhze+sRPHVtaUy4ry3nk3fwrlLstDmHGU=
`protect END_PROTECTED
