`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93O/lkkup6DnnrgfW0vmTehDE84/4DwilggabJOwJtxJAviBTpbmM77x3An6R4wh
qo0B+U/rid2G+yz2sI1yG2uhB6o+r+NHUZ7fLHPOhj9FCCDC8MTqhEwMztuDkSaM
AdwdMdkyyQ3gJsWYaJanIN1qRE8tsW1aBuebyRQzvNBQAcVCBejhYMTZwXi69MiH
EAcW1hQxAnxEJZR31Hh0hlMi7zuChjHbMfk0EC86u1tM4bgtYGl00iZpklQQIu3d
sGCZiQ4HUaLLBYzKfx8g4WF9bM7LQZddh/yQvNvY5sTK7ibshW1pfbh6zixrmux6
omTCj8nxazsJY406d+tK7wbN+LLVxpyEZbWGN3T9EbUIOCe8RR/yY2L6qNIwzb6i
kNv8dLduVTvvHiHOEIXKxlIe+JrnfW31Gw4CMtnCSrg6PmM5b1z57I9FPEiFnst9
kAZFtaaS62UcrG8df6F9+OyjSDNgrMeqQrhZC0XegCkoFcc6jhEU3TS4MaO/4yc0
mDKraM0nR3gd3NF1AAiCjdbTMQ4nnX17bkA+IudIzwQiswtYSILswm5M9+cU8sSp
w1bS5ssO1G8HJ/QCqxLo6ezY5ibJebvVY41cnAcpYjmt07aJeMdEYkR1ppOztb/H
QatrKjVvt62koMTn1J+cUzwx4UHdaCiiLU4rH7CPDubWqCo0vgv2+Z/pJaORx7YH
QiHwX/DhUt2j00SUrm3BW0nEn9x5c85Zad+xUFjFltjMKouCYofnglhd5XoTJWir
DuGPzPPMSR5pK53iOsatlD+S6ge5nJGpnQ6S0tp7yC9qIbVzV665akmNC8tYxvml
nW84fm1odpUIrlhk9iKKiq4Pr8yBzCvRBRTnuhkLXC9E/aBz72TcszZm6cpgwcJL
6MMXZ7OAqahSqRRVSTwWyj3cCLQlsqdsoZ1P4n4G+KqbAovIIbMwwg7zLJLT6TSd
fI/y8D1XtHjRujoZEQg6X8ddALcd9KoZA5AbxJfJkr3jI95aSPq3fo8jQGr0UfWu
hsig95iiuXIRGlRF+Y+Ovbk8dIuMhGegOG62K7Tm29cuAk97HMxAryn5+mRpVf+b
Tu+REMXTs0IujlsSZhAcLhcrXb+rCnKYcmNGCSCQt7SSD+4ybpOAWqxHtkvUFjUd
hlCsFg4eyjA472cSbkjM4FhW6jg/JzOsSZke5tl4vf2WWcpsFTwOUT7CvpzmXbRo
hw3+fjN53oZZA1/jHTTGThe/ZIBaCTOSKj6+fDEHBJD6zMF/2QOqT+Vi2xYBWauG
eOlRphiKbiSYOmy2pYAAQmM7agC6suj5Wxsf3JyDH/gK2ySziDHr/b9qBg0Cy646
Vnhhk+aM/yXhqRFWtjLzZnsZmdLyR4BLDfk54YRsEnXhhv/SmsFHJZ1hLIstUrqq
ZA/nIR80BYp3VKSXBOygNjdK5klfkXR1Cuw9pv+cq1NSuD4dnRWjA+Su/f+8Lj1r
XKWImOFlHeGVOt2sCmvbwWbuvXiZIeD9mm1idfi2kf3MXvxFjfryRaIwkHb6OVgK
oMow9Y6ejzCGEloYcPwRwM6/L0E1dLyoEvuryvZfH36T55tDmtxs4D6DTCQE1EXw
6KLFvkiYXStpuhzignNi3rm9ui3XshUc6eiJqCQUGAv3AJC2tnle8GZk6L9g1j48
Hg2T+KDmvo0NiDsncTuxYvpT9asAcfaxmLVbeAwB8YYDuGoxNA2l5tg+DeOQs6oU
WZhlOOPDFkbHclgikXOg3+px7Bh8PaQYM7d/pvTkx4kECzVZiyx+DtPXsaBIyy9G
2Kb9j/zJX0cla9Sy4imcynuZkjP55G7ufdrP2GkuFcpK3TEvM1NOdeNWBskLnuE5
77Tz/2Zc2DBypyEEUmEwYCTQZOEWD96Qjn9ooQQ4iz3B+KcFkvdu/NfcLrBLlpgB
raOS/042HJe5U+9gYKz9GHVRtx9Fd1jeJTmZr2R/A1fcyvA5eN8UlPRLdWuLW8cL
hLZ6zubRz7p29YyHjR6Okzs6KbfPIBNb2TxRyxkU/b4BGOGEQUN7uJwU+MxZ5VWD
ywc8n3ZHAA1VewYmJD9BnxlcvkOohNCQ1foebLEdG5WymhtB6+f4cEZgYTUa9Ezw
RI6FLglWQaYrUysxSn+SY81nQUhcHAi3MyZzx+6MYkjOtnN3QgYiG/1LG0j8+CmR
zEwRT13066ZdWUzDyP8WtWCGevsPtvpjOb1ojR5rEVICzDIrfSl4IeWpclI1RM7y
EPaPges8rz7OP2T7bmFUt3xAEcgmhyiAxhchFQKCw+1gNrBZ94/uW0+g3WXFcECJ
A7NWFFMN1+/CKselsWiKppVq2vkbzBhzAxLjc5Tx0x6aO8WYzD5au8+S0tET/gnX
ro+cqrclEbAZ01yGT0YUpo7eyKHTYRikp+WgtdAiACzBlsxYJTpMJ6qwVzTHD11u
YXw0G8W6ZbWOQ6MYf2x68zkqn14ithU1aYdPBQLVW+eQN7SApuUmflGztHSAP1Wb
u2ZjgAPdL0N3kPlmPGxbcCBHg+BHhPmb3qqBzEhm/GO+9u6EX14AaWJdt9sGcTsY
udG0Zu9Q/i3cyI9NNmX8jJcVDVlU4iIyfuBEQa2nkxZ8/i6lbTj6ZZRJ6rekhi6I
4A6Uf0JZgtt/1m1t2J90zr8onARtKVM3TCpsEQSB+GkYs7lnTqFcvKTfCs8UFTNi
6V6klMBlLwesFTrReLdO8gekLA0avUvmjMiurQ/eVItuFicPtK1CYGJbhylUhivB
qKTpyTIbVHGB/xD0ZJsNjTLMUBkYpLgBdZUL7VRWmnKz86Si8bHIw1xeo1ruX/G+
qPVLbHdjgg2oX4TPI86g+9k+Sd7PnXYo9wy1acjImX+POnW5x/9/bPVwznmcvPAf
hynEITvxzQ0Twxvd91Xi98Vtmj5wcUmx2OD58y+YcX12oyG5XTexY7UcktaefYv6
7g+HOBO6Kk5ym9odDgjQzNTqMUraVbLpmb2+birDtehz1pt8Camsw8pDpOQKlaHF
PpY5RcHX95ntSmQjBQKvEFyCqwT8QJS7MckaGsTGlvaYjze1fPS8aw396NlBrsig
/gbojKlxTWxI0xLs+jPDp2ROsjKYGK8rAAK4KYvhdDFYS0zxx8erU5mEdWS5a0Y7
AwzL5T2T6iGB9j5XVMuX1SgQxz6PAZ/UPECeoL2P1jx6et94wf9wgAWQWE/F61EH
ENYC8B7ruudHByjrGqGq378mClhYgvJDHVNeB9ANoMWAs+hhqFggYFkZoD34K38P
Oj3EBci+lK4wZXRspeImbn0Fi5OvlGQlUbkqYwVocSfem5wA77bWtqvcxAYtZuO9
6Mg++OTA7QHxF1oH3j9mJugn60gs8Ha+1ztXFAWM5QNxq+XtvJaX0/DtQAOnLeCc
eyL4nFQZynEcp0fSvKxon9ppIe8f0nYWBv8cVXAdxo5Zum5sexTQn5raLNoEn3Lf
HaaZGNp7DoPx2uaIAYfoUnMSD8BFKXewttEnxiH/gbKVKXU+KdIofS0zg2UuQaEZ
cSBU6Z6YRmVHKBVUoHIsMtHWEdwwhFwTum9eSVHOk8dgsH/91TTVHo4h8OtzxETR
0U8Bxpy72ywZ2m5bWSKE/p8elrWhycq+oXPdiwUQRJ8r6n2t1UTm6lbZjYIan9RJ
Wkk817roAr6+t1YLCrkgLaKRiq89Oep3fFDZHc1XZ5dI7jw33MWy4ZUX82R4K57c
RFu+283llKOV0J2vz5yxdwTdxakts0AWX1SmvNsJz3UNkjioemutc3jipoVf6PUU
EdoEME0FsNLSlvN04OgkuG5w8aVmhbvf9zvSuwBmaYnUUAH3Xy9V8Wh+udJTuxKd
lVjo8HOew1TyAZfxv3uoEkBrPk4Dycv+CgchexJvqgokVy3az0NZtFgYnYGdYQkj
oHq+VH7n3vxK5y3j1LhL41gPsYnKakDKYZisU1RYQTorkomjXp+8NLjRnbrfAJHB
4VrYg/VguY59ULS1gww+lzLDY81u528hG+MVDHknofjEePyqRm97hgBjoBeGMHPJ
HtWlREhjRxYNY/S8qVgbQDNYW9HtG7O4r8TtRpXREFXhgyWMGTrkMknssrK3j0+j
+r70OJNlufMkfJ92t4rXMDlzI4hprPZItyYmQuwV5V02hKv8+pwsBai+oMYRYFMy
3gXFtpXdIxM2qN9/cyf2iGFwYZegegEhS5r3zY9UTLyFod0Uq3Dw/AVvszYBdCad
3g/mIjXzevfCYSx2weTkFIKONSimq/iWVP5kHL6vKk9VC1OdxSapB6npEkluMihY
lLWProj51FddAKMDN0E0FEPt6x6wwkqeQqb9urSB4gZ/uNKsEAcmmROC4slRdjAS
uiRtl0stusfyKlL7641QcMInmLrdyeQp6ytbAShxWWp7UhAA/NRVQKUxWvSnNM3q
jI0jd9sRJTGPBhhj6SKveUNrcka0UWOOQTh3OPLMbPeMexe25Lz5IDNfD65MjihI
NlzEqs0bzsESwG4FoDnlN66RhTpEmxYGO5hWHZWHFZZildgJgKLRG9aIF+9eaA6+
CnSsD7kq+TJplS5wxrnt1BBUN63O0KBWBctdBTAEd7ycxR1itpyMX5DuTuhWpwwC
HO36FJC2zcskjiVEih2dpisc9aoehmGrkwTdbs0ubNLJmrEx6yVtCJYNCnnbEMFK
YipuGpzhfdrWIvJ64gkkuHJvYJu0pKNrY6qBOM2GOM7jH1wcOqwpH+JF9Q8mK/cD
uO96r1i4ct52Q7fkHQqwFettolWr01INNL/8aRVOM53A0RtZ73WtQtdwbUaDO3e9
Fh6EJXEQ9au1z0MhLXmPhwsVXhdHlc9A1D+QCU4T/s3F0UHp38CNTEhnCmbSxP3H
tKisbMPnA5tjK/8YW6kNw7WT6w7P8pj3GzN6OZVrUqtn2Kobg01eiWzTarddeNkH
0lvrgRrT2bmzgEKr4109kr7KCNw9ny5w+YKR1V9x9vxq0PtgIHuGt0ImQ+Tdd0vk
y6nfQo/xmc12N6ggO9r915P6DmmFfj7iHIWkxFy3XglcCSnV2pSaSZo/SmfxnU5d
eYXjHS2i1+mIlIjSEl4uqOMBheyNavVlj2p8rLgDkCR1exGE7FSX8W70vXNkQ/kj
lchXJa75X6pOh3VPGY5SwLINlINFSJgIcDpkgYqp+EdqhUd0g7y081qDRbWU7yWf
Ql2qC9WqC9IcmzvVmomfbV6uSg1Gp9HlrxywH69EGg9sma0BBKRQYOI2DuxhqfOq
Oj+SUOZuWlONKjN9S4wBTcwjtccN4VpkwDMg576o1vP5E6kveyY211/WZOBkodWx
PVxTCcx0G0DOEmNiIuxc1E+uNtCdnswm4IuRh5JC2UqM2CRLMZ01juBCjNDuKj6Z
xScVVWGgZINeuXi0VSynxR0NgBhpfiBiDmcXIZ2hk0+efru2uf1Ny1igKAhaO1DA
lsiVOgODro1y9YmyLsXcGGwSW4Qsadf3ZvOKl232CxihkEWHXJ0PC0lf2YsqEZVq
iEoHuI4UyF6a/bARnNzF/TFNhOLvBKc8oCQh5223ZMYDVyOmHua7suNC7CfyQN86
yi/5PvKvPKRuoHD7jtvkt8gQHc4VV+5CEtIZpiQNV4F1fBgRfsBQuLEgrtwX1Y+S
uJcuTwJJ1vVvWfXOZ8AJFk7bUGmjtidxiFDzs1hQz1ecQkPCAFZr+ZtcE4JZ/c+Y
RlFxJBxwZo85WvKVysAsE/eyMOa8J9PSD05flueO/+YVdIpGVo+j4iqTtI0d435r
mGuqnnzUVa8hXgk7B+h7BzLuIElXs7fWUxE7PDuAIKGQ683w2hRIUtTLLo6+4tGO
Z9ryR9yJkDiQ9UZKf2kgJADpXBnp1/tV6M9b2FqXH4fRuGJV70Ld6me2f9CWkT1J
vvxS+43peeiuXExQNdyuhbB+RLxYbEQjxi9piCOK9l6Wdji6aEY0/ZeKQ8ebFzjm
miUxm00aibLngJPxPs5tBrfSwElwUq3MRL4+KEwHNvuWtMHez8CYUfeL6IUHSuKP
5tW6acccu+8Y7eKWUFf2rQsJnqtVrVKZ0llX+eTY2fbs75t4ZMXii2A/X1EVOCNd
qGKAtD+YUqs0XA0uTnFcEN88vPDyVfsRNPuxncWWKHDoX3cNWeJvjJfAAIfdBr9u
ZlLEbhhPOWA2IoFRqMp2L9LQiezyK6KMRptaZnhUx8GJZ5dJ/1nd/yfIpMG760sn
Skcl+Ck4H/MFVflg9XLbhCzWBgzQtghwg0QDT8cMdrDjbDXyVua58T/HOmVPPU6f
cscBMZAO3QzijZsm992GsiWl/G87uw6Ak4r8uQAc3oQM8fHPs5dZ89ykIpPmQW4k
s8IY9bNUEH4okMx7eRCLg8+MThqYYDkERLcANpG1mEwk0+v4sIZfEKcQPEhMXbBa
uY/Ho4CU0RkzwDdHtm4IeentQv0sVvZc8+u8AdaOVJDT4hGoJ8JXy+Y620PpyC/C
Afo19KFxEv2wr+VLCy7RU1NATlduLH7V/rCplwplMVWcwoylni6pHgbxTs/4Z4o2
/7i8saZ6fCOY+biGZWAAIp8zwiYKuHBgq7BcsB9vNIMEBLPPEsQ7S6Bq4RIDw9H/
vjQ99CJkYIpeIL/gMpX5x6ifWhFQ9J9r5FB+Rr6tZ+VNGrc68aNs2DwfhdPbsYyC
nlg5WdgQjn/OB5G7qr0dh9ofrX3H39Sp4m+ju7bWG3HOfp5u0dPIDjaN8GoL4WHC
TEwPO58a6+Ddwa6G/BQEVOpxnMVZ2MSEc7jgOMEZiPYO8kYtBbsIseVWKQneAdDE
HRh8oWG/6Jf/q8EsC3XIH+o5CfRh75REVP4C+0uf/h8rF3k14lB3mj6Uc9qp73EB
WVxKRI6n74VED2NQhp/eqje/oVU0xhiFP1g9b3I2y/d7qNScj7v4NnqXc/Czhjfw
WxhWzTFX2JWTbPo3HOempPnR3Jq7y09As7zV14wDXXOac4A182SVUWINiZfeWDWO
UJ4TLQuCuc6yRKCaETL+kttaBZj38TuAUEMaYuYuwVqJ7PhMZe4Xpeq5rO7zj7vy
AURpwBj3FcF5jWfmiLTUqxCsPkxlo2hw9RM4SCUctSsIvO+oOzzarJtHAvCuztlC
ctsYn0k8IWzgWfASMpAvfqqmq1ys5OCSzWd81noOsAzucCZGDL1qtFQbmDcwG2MD
tIgfeTRGiIxPBi5Etk6jcaIXRVSN7dZs93Zcatkte8XFMYKIHzXNUJ1WrcaKUk09
pEiqcVzEII2Y8X6BmilsL3YHmHbDdHbywgqzm0F2WAWRibcyZYDdEslhQCZttmK0
zDo8zS+IwZMtKBPPV3F/YMEyucwiEboZX1Tech8oZeiki16hvb5ZS51C7VXNY0pn
gUF2bSfpZpnO6EU9kPYnzp6SkAexIN3JHcpm8Y4k9WblHOL38T2Xmnv0gegCRRAh
Ff1D0W3gJFGcA5MVD9q2zZUpFAOkRi6pVL2Hk//bZixX0ut3xtXNnM72dCxc0zhu
r5gTiIv45wtU4Oo+HaB1cB07mU8a7e7BwJ20j0KDzQojqG53ACmX9Nkiu2EtCUIn
b5InYi7CHrFFD+6RqChZyU9Vopg6Bz9yZy8rfGB+PmUqg7ZKY16kfcWgx3iOTaZM
jwcWvg6nZvtAGxcl8iZvRvpo3On+mdNL++mjJbN910Fsk10OL9FU21XgU2jE2dc+
vvomVVXtNBl98WZLNvpTuUt+LmO6hJ44WoyidX+SHSutkrFcAC8BqFI/wSO7AroP
GlxluiiqwgSOk5ZIzktfkEAG8XFTtX9us/iu3pfAZ9HESm4RlDJYJZ4xMygx0NP6
kknPo86Brksr8VorADwiAIHZi8KUNHP04pvIAnYvpU4=
`protect END_PROTECTED
