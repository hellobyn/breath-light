`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpZARXt0FZmmsFlYYDHB7wQ51iaZdxNAwvJ2N390DL6V0cCd4BLh2U/ykpmkzGUU
mH7GwtfWzWr5osYOs1aKoonKixpVeVE6wW9LuChivWh1uuz8HrRVpaSifo6Wc4Fd
YRFbvl067iDbExUFsIbzjMgLxWd1ys18Ie6KKVieEorbMP2A+cNGusPx9BLF9VPE
oGuefr/AXaDynwUyTIOXWtzZrLupojzOLyAVqTecRsDkXWNAKyImgNF4yxf0j/9g
eZxg4y7I3WQUXmtWgG5Sw/WpOB2diUJuT9Cb2T82vErUA0MBfKzMk41A7rD2yp8H
8X0zAXBfPomBG+4+QEO8fi1ZxQDO0yfooKxJ6TJ6Qv+9CvMJGkkk+7l4W4KeYpiq
FMyJq9prG8XP/6PiVqG9S7mIB68Hl/JZUdcqOD3gUYPfDR5HWVgsUWl9MsQEeZYc
1vsdxubefyDo8X59CmtRLIyF24n4AFJPNjLmmgri4+hKKrWAKxrs4ftVItjAZBvM
n4TCn6b5eKq77RT9a2f5PFH0PIIj3sm6ghr9nliaNEt6Atae/9dM5dBnUrwyOtAp
qF9IxcKYmFcubE048C/z6w99kJSxKAx+lx4WxSkZRgby3NtYlc0vxiDa56NcTuKm
NXjjWAuUSCElZ+B4Fee/Gqa/Ngt7l0ewwpYQmveBqXZLFCJf/JB/tf11qgB5sZzy
uUonhXvLbqGAiw0ktho+mF94JIUbBwQMkriWZCPZp3bXX4AcEtYWzMb7bZXBDZ2q
Aiqe/pSoNaSjlQA/OVf0HPs1eeCDSgftNSZTXYnhN3HHWHvRRRQId1+VnpaNIR05
JD42KF2w+s3KKPg1PoVTuV9z1dHZXunmtpVRPrPfRLZJSi1nhYaqoxYk/8GK8y9l
`protect END_PROTECTED
