`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNSW7ucYFXiSpDLGYhzdeyljICZNV5AQ99HlISR9Zk6C5H5VnS/b/7KI8CJ6uQmn
33yegXAfdX1uUYwniYvYvK34481RT8xou5m36bB9/k1TmajpBG2YcU3kv2RsMixk
SS/3aCdiInwanIv3zFqE8x7Vj22SLHkuWCM3EPMLjWJWHxzhPjK61KkVXsFreE5c
7Iin3CYeBaRQbafl6s/4mFQpFsefx8i3FB3Sma+mw5fMr3nkipj8idylpZ7bATQ+
HY4iIX8v//s8w4rpRLIjxaxDTmF2/NMPIm5J0pfdcyjuqHgMAdPK9C764av5pNvH
3sdKO0H2BkZ+SyEBIeLMgXVde8+quUtKhVXYJ8BbCY8MvEi8g7IyGUR0FyR/u3XR
UXxbzW4iYSvM4csKS8Vw02q/LIteblsAkzqXq/zLWmcIEuZqBjbQvAswthXF0Er/
04AqqrRtv9EPx59QBqpeTv/c9A4b/OcE8iZnrT1qMg3Fr6Cz4uF7tP5vUwNJ5S8m
AJ3WlC8wQIMPgvpAh8tRGTBMsCIMJXmkXTt3hOdyV26KunbL1BOgj4jtmzoatSmT
3hmg3WoLzkT1bH2lDqTYDiaZK1f8QL5Y/aXM27k4G14gAnPM8CI9ekYDI5wSUrGQ
RrRVEv/Us5S2EpyXGZ5JL1htuCmSURk4wgQLzEpjZg5LMkDpCSuFUWJD2oT7GqhY
TVfA/QDJ7zxgUWRO+Iu+IIL4xWLD/VwFWeuN0eDS9TrJPctKkm3Vms9QJqpH5Uts
51AzQQopkGQami62w03eGPiZ5+ORzfMgKPa4Kbr8X4dWXbsDksAo+8LPOIAVHrEn
KD1GWRKptd2Enns0V9cb9EmiGd6qDmEklFu0Xpt0n25Dd86r3sLWSGDvGv+W5+8n
WS9RfULJBw5YlfoCljeiN4SRgJt2N8vIGq+7JgRKhtDfJV7q/yFtRMfk2djUIiMk
`protect END_PROTECTED
