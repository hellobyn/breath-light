`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORSI98eHPpvXdhfqLkIDcT9Uq96h7YmxlBrBz5D7qvh83FpYRqyw37WwS1NGgd/j
vwwxSpdI7W0wXhrq5hNUtZijnjBUvNy1cAw6Vkx5jpmjDMBb0vtrry5rqc3d3nfk
tYLrVpQVpsBJptPy9du0pv6Bg+yhN5VfqNhhg25tUIN3W8sOKd3kJGNoqvm+hOpP
/YpEigHQ/PLhCJZXmuiQAX7d1NQeq7rW/83IuoGDZiCCvt28yjCgSCXeqJrP/Zmv
hLF0v9VC47z0qt/RKyP8JJx3EqE2/sglqBsKr/Vvl7wQ4nvo/3W1a95EII7pKM8w
FRdjgwpbOWEpe83zCzYp0XQMBapJdCGmJfQsiO7pSh+g+LIrIodVomv5D44fgXm7
XLyQo5bW12HozUg2VFeElJ4A7FDDZApxH/L4Drmc/Iq5+NalVr/WpZGHjwIMIJmN
aNRqfWx4tQ5bhbJ/gK+Sw4j6VT2efIr6KS48O/UMlr5UZj3HbQ3d4WVibEryy95u
D9Svq8C1JoQ1ylsgrr+zRHRl/5KYvrdcyz1Y/v7NKV9Xk08Fsbx2n+psnBOrDrIK
aot+AojRdj4pFu5UimumOA==
`protect END_PROTECTED
