`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PAdRX+pazUNaZN1gcDhtIePpVNTrKqkzXy/U3SQA44GPWrrfhqDb/+FM4wKWPYKk
y15UchidMP2b6GaQvC7r/NCmq6O1KxwRVTyHOKR+0fu/PtkuDt6j5u4TNQRFAU6M
yBt1n320zmr+BZNq8+LF8UK53gLCC05/sVemVe8XLEplElwkQ2oJZAtfWUjWzAHH
lL4eYqoiIITawt6LmERt4hgE5bvw25rDpYJBuN4IwTmjMKQpgUZJyBJ9Py04auIj
VRqXSEzN0AgZ95A7SiEMEC78Kyt7WluJjxW44GDGK9vk3rbJPJyai5/zMMeuCkus
k5eudks5j80ZkJSLOb+cpMKbzGPCtdXgULnmQpPnE/RBss/WFEZ4X/kk01oIYyek
xe0lXfdGjyT6y9eGKlgPgL99uivIChR+6WZdw6bYSStXtk9JLklp/6eBqHEdi9z1
4Sd5Kp5TNW30Aryxx3bDG9Ia9OYhkKEtwIPHxyy8/B/vvH9umXQrFBmZyL1O4GqY
55kcR7QYe3AVeInFre1JCavecFYiK08F7g8KWQI31vbMmNcie7c/16KDH1vPxm9W
IjB6aM6Tg3Vx7qxYgNC3oXlaUOXBbqrge7Z3z1cOCllFP6Sb0qJ0lRjUPdhe9TTT
NniqHC2d1jj4fdnu3uGfXy5CfD3IYRutw9XGe4/MZW2Z7UIg5oTki9u+STmLYF4H
7uWJUob4ZzAXAmYH8GPi0GDIEnS0+FLMLk6qQ7hgtPCnQxrEEiZaXxjp0W1K3M/m
p5dnT0mtajBdmqnpFyboPccqiVe96xXEpgwSEs46mrM5I+Z66tsSya3OrWrvk6/5
b43kqxBisNLQcBpdqtkpyR8zMG5eKKHYH6V0HmW8aHUJMMuSPgsgMnFvZEnZS+Kj
YgLsCmObWp8pb2EBef2SD3jzl5AykjESDjnAm4Lrz6L7XUUaCq+7P9Xbc5dkJEhS
cZAz4nTBkfBGE+9L3fST3VKi+qhlO2ufSNft5mfBCGvQbRFSLC+GOIBdi20H/BFz
1XauyCCuI3h0xpIGZBC8bvPP82eMgdfcweFdnId7eTMl/uk2SK+q7kFZ2QK+m/hY
uOLCwWT3DDkmt1iwwppLsX1l7u2FPXu7Lp9efW0Ks8OG024DytYPPvOIl1ADi7Mj
xwdAuFuzXPbOTIzuPbPYSDRZfyKbKDwsdGo8rZDLqtorxHFRMGzCVwg4rDf7145x
4IwaTb7ZVlcfkaFYLSv69qZEN2r4dSWS4Wnr5VkmmBWnbKOfmMy4AK0lV6kwpINw
hgJ5UCvSZTaH3xzueEymRtA6Tmk1HE3B7VHO5lIUa4pZ65yjmFBHrZ0/GmA7Ui8G
vi3838Ztg3i6HQKS6Ul4C+kS4yw05FAwKngUPlG1msW1LpG9I8BHhbGdQhIIIjEL
6M803IEGtgMQ3+W+iby4SphMhS9fy4nBkPqJzTQfneDgTwk6KdI3QxIzutMz3Ld7
lN/wJXMmuctyrzqiOSKgiLdeDfFzf/FgjvjZvRFGik2apawSWidUjFUX1m8rgp5B
d0ZFN8owL8luPoT6yn+d0JeMK6QXVZZOmaYW22e5kNTZJFr3a+UEesDj3wKYl+jo
xcjDh2UHGinznv8E29MCjjTEivfhfkGPAb95rARe9DSowz8ICmV1luQhoXYBkJaZ
GfHCF0KOaWl4k1LJhL1TRoWZLvYGLQrqjHfotj8ITAE5g94PeaJYzxsbF1fL/2ih
u+M5EmD6WJ+VjsBq0RyGVfqEwA2cPXCsLcGCpvYAlpa00COb2IRxdw6KyUhv7SeQ
GP6/NKv5rFGUV8pl9QIvJfCawzEsts8KfMwivEDQGKprTwMZHKrg8shZQiYP8U7H
Bx184xDhc9HHlzVNYr//u+3IWenmQsYwRWg9+7N5SmQWbz03MgQjiD5Lwh4c+dJA
ubbe/7yyvrDWGB0aBS2XYHJO0Gjlv1a04ivGmTVEntodSs5T7d9nQ+CiFsGD3ddQ
gk+xQmbV4+SzBgcL4kfnWnA5zP3iNbfsc2Rp2pnUJSkSO594JfbAiKdRJWnJ8waK
T4vZUSOcreFILEGzET/zyu2rp9Vo+2HNq9gXHBixeyM//kINUVGa78c+dXHwleAP
Rcho8D21K4oslaXDm++X0WBxB9UouWw4OvMv0KsPHcUjOEdCzOdztkoBRw0vFWUi
Z8Nh5j0oHBNSPBQ/2MLK3ZmRyNJ+4uDzUdv1ImtxFsQTBRN2CsE69wT2lrh79WbU
F8fStFddC4IyYZwmNvRSfJkd7yznpsn8cxD3G9/NlbhAAN7q9N6QYT1QqtEcyfq2
3m0M7u68PHOw51TjpYdK3eHSPsaluv2VX0xMc7h6N3xtzdvn9UVm1gWUg43/xmkt
3FlTkyPUggGS5q2I867toxKtiuB7LFlVAnxWKx62n0MlznW3SNTjxMejXJA9UxjU
d1wgSBzrLO30/DwDfHcpseKXjjjMNIJ4GnGuGk0c6m4/s4fVKteqZ75mccQ1kAu/
MS2SEl958nLUbQM0v+Rcqd+BOZaaZI+spaDvniqsHFi+8Rqhj/9VfbZ3bk+TEdKK
dIPnXn6bvb3HFqNzwlkFCL/XlRNNgbYd4MmueCfZUG/VUAS1Jdkughk9I5sRTbx6
HW+TvuMNYsMjOLjuoep+x0wFdqsg4Ifl29ggxxNfmUQpiC+HugS6K8Q11gx4e/ix
srh4GUPhoiu7HUs4TcFjflx9KmRxCpqlflh99nDBU9Gln0cmSpS6gjK7i6ubmP0b
LfiPT8K6UoPsmtaNRswUIX7P/8n03dYoUjnsENYtKKrdexli5OEvqd+a13sSUZyz
RVR0odROEzOaqplR9B86c8bcgY9/633teNTH/fQQFvu7PR4KNkL5AhCftB1GAWn8
vSv85jEOv7Igc3Y4cTPfxZtYtRthRNLZA3ygYTNsiZhNCW1edYXa7m8eaAHvYoe/
u1QYaY1hCv3UBm0OsIBRjWBhqxOeFlgyyTRZRF6CpCP9tV0zo1vxc5AcQwcTwxdf
1V2xoKNp6e783W0MI3jZW/VjbndAs+//0UupCUwnKDvHok756iHNDyUc4HzN16kD
UhRCDoToJXKCF0ZyfaPG7gMPFz26CRtb1nAoqzvqrhLJD8qoqzmmtVZCm//7dT3H
zYC4G2QceMnqfNN7WV29MyHrkhvFZb0oEdf+dfKfVuU21BlIcBJ8IQG0dEnwedh4
SUZCGfZ58w1YT0N1T+vBHx/yj7mWLYB/ncBid8NZMwnZiLfkOikU7+Bs1qIFl/Dp
Bz5zwsQGeXWnQsw+fDYoyYFAFRGz0CwmsfHvXhtXtwBfVerFn87vkbMX+bImrqdP
jOZj4kGnQJZMkFTpZn3rNdG0vzaz0tNuI2OuKa5YpgAmjeTpJEaFen76QQkFHSg4
VPecALGQZEkT7JxSlojq36NI+Y5oTr1kmum+C/QlkLI=
`protect END_PROTECTED
