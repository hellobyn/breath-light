`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCyRQKJEJKUugn5LFDHsomt0lseq3fPLyLjpDFNYUlJdNZfubUUqZdMu7+J1HDhN
7LtEunVVYG1sfblDzqhNnmd0V2ics39U1NwFJgeLDLbrOcE121FYo8jdmB1X/6Z4
E8eiEaxqgZy0ApYOFm+319cyTcRUse1Zj/gfVz6Yusvhs0Da/hiCvoWAcNR7iYCM
JSTB7+B8FLPT1eZ23PRVdeBTA9G44SB16SAb/wdI8UkZ+A1gE1I7cVzShgGgFDRd
3XyKYiL1pHjQx/Ab5uhzWsu+RCcFpQsPF3E5rmtyTJNCiDSFA2aG4fJQDgRrrnyK
mEzsrVgMIwXQeetVCCPOIWiziZltGweSLQazLsuOLANo3ugp7Xolm+0FRKZoa/he
sQBduxkqT8JdiZHKt+INaGvE6I7FpLqib+oiT0CayTLDfeQcMg1tpQqqZEsvxugs
EYYoLvuDjVtMrTvSBSfvWnFmTh+mmYzLSxYtRYN+oJ9waytmE6ZW7XF1ICs9TZC+
16p3AWyuWncXNhqj+AqJ8kVSsIitsh5I5eSPUqzt7qLwvZOBkEsufDGSIjmjdxjf
I/ny/BBUPCkqtqhUZlExDiR4XKdbiafc165XVDibNPLFSXuint35kvPNjbATWMoD
4eQyYdveMX1p/nrxHSdUwKfBPeov6Q7KHb9p/KX2Ob5aiHUk781UwJ+LMyykJ33e
wLnyN48AoCjf1Ar5hqAEBu6X/qxdEWdwtqSUB9JUbpBniH9lvF7S0drEx/AqBoFz
371dEN4kHBR+N3JIDBYwGhQT0QdtPRoWbqZi0aX9Cg7HkYS29+qxqSOkgXC7/ymw
VjypIvzhMrggRSnFGuNDPS6Wykptvl/NX79HRGzuIqAQ2ckSuuHKpR9kRDUKIaXV
rlJc5SYn1UajfxFeKC27Tf+HVraiZDvy2kBsF4t0/d+Z/CXUv17aszCyJ3EH9M3S
R4jOKOcU5cOQIj2UVujTs9VR6m5cqqb+eNa1KCUK2IbpIqHsQlZRO0OFor+isqw6
XzLVdwxbgDxBXbGpKPpx5Pa/nOPTd55S8VPV539+Dm9j4VNIVDJw8mf+H+JVd3Xp
roWGsUMWzXqZ0jnrgU9DpOSUErBN5s0QDQ4GygLaDXLSiQlvi5eLVLrGxFnbbRn8
LrhwAZTLd+MMwgtdJacdyShBy3cqbsHyi/yWmf+lIFhTh+rr19/FgUojRaTQVt89
Px5OdkySyXZjnwwCPrxROFnLFzKMzF0505mYNDQJ0iybGrbxwWpE9rKw3kaiFh21
63Cft/ZRSFSl7ssdPla5CqVMnPIc5xLiGJrovUkxEmtUmpb29BHQY7f0/eno3Vp3
CDfXzuPaOfxImZ63uGmfj7ZnmDu1L2PK/Jpg2bp+jNwAi8tJqFCJKMxEf52qmHx/
eYqdFoRGFleb2LL5UbF3frM610ikTvmBXmD2Yoy5n+nERszbQIofoPjgPP/Uc1w/
hupxLCO7n8SkJIucA/AZ25TVFbxwex2Jb4+qCG5gp+XeitPFYDZotBFRyNdi1JDA
amk3RJ+XWYspg+42lXPHZToxHyinal0eqxbtKzSW5dmXZ3JBeJHFbLrCOb9l7BRI
81guu28S0cbCwAx93o1qFMdU3iRx4XMympHfSscAuW6MG92X7KbV2Jwliy/GO6Ks
8ndyR+0v2Fuga/2JGpqgXw/bW0dfj6aVlpUTwgeP/sk32HX90EqTJQAonXNfvojd
0ObpI4ZHnjZQGsr+/Tkgi6zMXzXNk9fYAHB7tqTlgtC4Vj5wJPqFogwr8y413ioo
AQlFJ9fHO3cQwjqKOSh7ee0DtdBEflIu5HGVwGvq16o4cjpsgHxjBS9Z3OyCW0o7
`protect END_PROTECTED
