`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIpkgIvqoFfOBNRhNojGDTjaklMVGAyievegHyp0Zx68zBB8M7g5sO3jLaAJ/z2h
PPjY/G0PPo4qf0N9OUL3/gmC+dTuJfo79mbOSeRqHJn6AxH6hmJOnfVD55hLICj5
E5yxF7gcpGClCBr1HFeheCO7sqlIUPoryM0j/rbXi9mIcPFLqESvCdO4Pp5rrMom
MfnZpoDAueCuWIJ3beD/LCHto+Tq7DCtdDAx+ZgPTRl9zwSLu6Oe0mGHlUULczju
To6AYVRgCmwVVtEvNzDo/PnMTdnCA6Zhj00BWZAo0jIjcAEhZWmGz9Hr+Ng5zGjk
YsdzDtMOwbAoEDbcWgHY5D11gXplhlgh3utnc5twcJMCPF8YYTnHbeVmjqAEDnS9
PlF4qMYLkEniq5zBXpfuaLzOWzsmDX9Y0JgyjWcadcmkZOdXThowEcvpE/Bz1GsO
RsDgf5ZqF2LoGBOPkrYZbhHz8BYOrKm1dUzTga7SVI4KjUnAz6Fy2zIFThkmFsRN
mybQZWwCvCzTrL45nx/iVwN00rIMuBLCzfm9mHC858PTJ/OAjrTw2t1eKhRtIUWm
/AF3CWPMUKZjij7UBJi8+Pto8iNHS8IeXwYqGSCVj2ED+qlrwXLxhcNGdI1zSosy
s0sTm/SVoxs4+9Z2XxRmuFCo8JBSKVAnqnt3JGUL+VyFD7J2WjuUpceZidVS1PBI
iT/Y185QPME7wUuTztbYCAasK5dVqOcCkAhxrj3AtfsHQzGIXhWS5fz61MWSu+ub
iL/Nxdcxrt1Uv6R2p8X2etfgU36uGWGZHcXG88aV39R0oXhWEmOIUmULFElSGtbt
5RAAwLVjU2XIBkHfusceLS4ELP24A+n3jyBBNa2N+HJ2YXpV5bcdTIw+uMkw1pRq
v9FTTmIRLvD9ukkuHB56/ma1/QCwV/nYycXFZ8enpuwB0zHAoqMsg02hqLPW4FOg
xUQ+pjdkeViZv7Ygo+wmv3oPkjHzvUXmw1C4qq87kv1qHox9UUpdYn9hRPAgJoBH
cyLD2mAmIyIzeGgKL/YEjppJTpTxJrkrJmJ7niLPhT4hEGnhPGreuk0ruPq8gBQI
FQFBXkDfMri4qFzY0WoV6ZO7mzEdXSGfElzvOCp4ZLxT7rk9BozS2aGNbZ8UBY1d
vtpMXeLSyHy9mPiAkUyHmVyPOn5tqWXFNAh0HeNJNO4ae+zBCDjLCJTaJoxj6uBz
3SpylDoB5KWlWkcbM5WzCSNL5jbftKA0aWLzON6qIv9KenBLZGZLKlsB/xguPTNr
CZdWo41JPhPHQaYefWdTHuRq+juWGpaMABlssJ2wFVKHu7x6KchCaVzuurt/TWFr
sYmGh17uKaB39kwQpS5wQf50DU+mEiZ+4YLAze6n7bwsuoMUXaX/qFU6MDaJgXQX
GCyaWisrhH6IqC2fslglfgTSW65kXQfOZB+wlYZCa4USMbe2N325hezkg/doALPx
PjWifS42hVQ8WMbdKCUvktXl2yw+dPB3vv05YalT8gfnrgsL3JG7b7XyJ7rkO+wx
AKzBjdQzzOZtoY38QOMYDFia+bDIHoF/E3zSAfa8wB5L86w0n4pnLhpHXuuDXLsx
eqlHAhf+LE3WIP7wNfiD4ZorM3qP9UUFsH8tYJsN+yYgt+Y1y5hpsh8byqEPdBT8
wx/lGA40IUFSqY4BYQeJmaOQJGTRzO+9qNRrMyRQodcZhJxkSch7BZp64PHM3BQz
j4E0z7z5Ei7B0wJYdRafKdvNgP5qajn9LkzTuHt1VJOOsMAU0tdlazacSXCxqFCg
pm/HAH3UTGzO4hXyEdBpC4ipVC05R2r8SCYU2GOZO1VEHX0TybAakuQJUmBvxbY8
dzQQI8DV3VHew0lAAN28aUCUMLp7sjZRZ2xfnkCnmIXBBUHbCFn9KiDrTq7ATjnP
0/uTZKSu2eDhVxvZANHIR6VGZerdeE+q67FTNVMZr2+bXvCULsvotu6liSd8GWsZ
uihGHBztfbiX1Yp1QqzIVbYP0sm84npVXFGNnJDIZGZcWKBPTmsDGGJTPMNu58ug
Od2FJHmqA7wTQUKQ3WXD8zNa4FjdJbXnA9DTgqsaxESouop5jQHwlMvn3GIeyHAz
3EP/NpoH6egyrimCItYUzkCjftyBAB60gNd2Qmi5CZuhip3SrONN49MGSwFx9HPN
6jOXvRhc1xBWJvk1ZDuFIx470Ol/QcMsxmg0f6ZxNBRPP3kVhKa/AQbbKITVsLue
VzB/W5uBV4QvrLwJA6OKlvzCyvBRPxtS6EvR3XkO72opvtS9dEu/wBdBDa+Un+Nc
dANZbkImyEq1/HGFr4BeixJ6HuxS1/YqLJleeMqUFYXXYEHY2tbgkXvBVOsknLQ7
eNwFGNkSHlOjXkk88ucTLY9FuAg62Eoh9mY67dygRO3yFgEyYH1m8EzmlpQmncJ+
LpeF9eay/SzOoqc0T802v4hbysf7MmHoyDJjtOnQ2fh0ZVGMujdc2n7jxwECmXKJ
Q/1ZG+8FBQG/c5Im/95o6W1GiTMEH1RFX6LAji4jxUJNOuqo6x8Of7Ej3PMMULqU
Cel/D3FfcBvQI0mI4GkcsEr5P5xTy3LF3cBi4sfW86jCN5a0MNRDtAa6J0pxQHBf
5AW1mcJV6r55BE2OL9kRH+LzGkV2D+yBhjedPvbyF5BT2VQFHJCw6owrAdxRWwKq
536qlD9op4+tqrocYgqMVS6LpdNKskks04pN1pG+3gRzRw2u4oGYFSgBlf3fQA9B
Q9eI0HiI625zrjtI0B7yhhf6M2oNjj2W2Ev7a1aWUouz0qytWNtv+gPXzCaLhrGw
WuUYtUhIbojyZkYAl1/5IWBrqhGQ7YYi2h4QdqciqlNjb9jdWoR2lMv2DuV/gQ2V
RCu4Crh+8dHwK1WuCVuCtY87WgD6Kg1SEZQKKT7zO7zfRKXXYkp3/hua5uG8/d/q
/z1IkuNrFkKWXX6Lg7Cc7vUrO72ynqg/F/HgrGkwxrGDzwcDFjRRWYm3xf97Dn6A
C7gBaGqQKzkMJge1BrpWmbxUkWOtZiGhU8HaC2ixfkB5zge9Cp8l08fTcsALjLnU
CRaJTrJp0x1NU9ev+nEnayuntgj9C9YuTpECK7PDbf3CFUQgwFggVY8iOEeP/2uN
XKQhsto/6Ave6iLRF30QL+stPOAcO7PN08rlggIcWcmaj54ln9J8g7E460j2Zghl
ZO4fZAbH+x9bIpdfpomBSjy02jaN8laioc61T/7zXEjpSraOY71O6FbH1pz/WRca
IAMqUIavJQ0F3/NNv96pB6Mfr5hYopW9rhhuQmJ0NsrJUuNtWYFhAUh085arnit0
FvHBOsaKbUkwy8VmdUI6/x4Cqjk9wENhqCHDmHRi/eZiYfEo/1BKwwKbdquQuj0M
KX4yNCmrC2TiIpWAdB2hSwfBYtm1h0Jze1oU77btFIc5fzUl2G/6GKH3cFGqBDoy
UeiuI26Lrz0z8+j1YsCY/D2WF3XGx3WjMG0h35mlbmk4dXBnoUHVZG4vKjnU2Rsj
iGz777LSc/dshlN/Digt/kowsCBrYOvo+P+6Ulvt0bAs1AHHYkqygR059dvGH+rs
mg4c+T/eIQm73W5C/EPm80PGZBFj1DokiJSpXPluzn5WZfKe9+lWgSbnAAK0uBrG
pW4TGUciecMYhfxJFcoIdfUWtDNmbF0Tx28h/iQoeHiFQc2vY0p6r/tue3ejxN9v
82W5q/LswxAZD8DljWqYiqScgPZPDwFGdGveuRnj3r3bBTlnJs4MHAL967+l1PAr
5AWNH0UlqqqLces5/39OTqc2uWAqPeQwzd+tVONq81WNIaCEbGR4iPWaU5MrkgtJ
p27Q0V4stE6odgN9bMtJklva8bj6YB+oB5QILc2QcfNJKVVDVuvVCkJ47cOZmDHT
/EtXAIAQJogD0hM+RBdFKYrb6zy9/6KtIk3IPU5eNmgwMajtVPQoxIWi93An3Ui1
sDJELIXhzJDccdp0WMH2rOsCV10Em3E+MQT6cs9VMXTX5fGFfVzGOH6+oYryN4La
pkW5AKVzrCN364Fiil7qfktVDqcvUsQWcniOzbd8QCzmeHdfegWUHm+iGBr+iOzL
Z3dQXO/k+xq2OGA4rKQfkIpmrn8GxuJAKZl52KYBkPVQ1VBpbRfJzwbwN4HK3zXM
Vf+WyHWbZf4Q31Gvlr50wutwSLo0bWw0QzBx+zkrBsRVf+TA0ku4ALQhuwa1ekCA
ZNqefdDj+hiMTSK/I2K8wMU1jBK3xQLRQdK7kvUG/zPQb4v6nxEzV6/Dt5Z2P8o/
IPHWsjdv11Kwniqr8TeOMGZlXyCdLfnQiJ7zqX4sxw164mZ46leWpn+S3H7PiwYg
VF0qgxvnFuRnfMTFgWMkYyR746GxBhtnTsUIYYE8QqJ4yiMJ8NAXKFfmvvldtwmU
XmwBl8zDkyXuLuhg/EkC7zLvaLAm7RfNqoOCmTqtVXX69BsnLCzvCbtrBE3k0G3S
3AmcRezP6exwce+XM5/hx4gYFDc0UYHfBFzPtOk274Vo/Mxkh8SL1PWt6v6Iv9Rn
cgCaHt99OCTPpgNEwaTvzaBMLlsAHYZLEzF1dcA4SVLhsf5RUEFK5T+Ne6+U4sAU
X9Yaji4SwKKJfG51qYOwKsYXp//hDX9qj6zbokRqj4JsZrHtE3rKZeYe0q5NHNJi
1nH4Tk/TzKyxKgqSEhob+b+WmzyQ51mFDVVEe58+Y+La0yLm+bbrKHRCzk+TEGiq
+ii7opaQJWPLouktwIr+kogvFKGwkB5+pa8ntU7SyKNi0RcBJzqmKQq0CQoZxNan
J3eZhZrjgcgEr56DUwYSdAZpN77JHdNd46elsAh/S1nyvcuuPVY0HS44T0J/RqKK
KdMtNHxd+ysBi60Oe8zBfX9Tezyj/OYZn1M99Xjhyz2YpoRtLoBqy+lZanRtiFmw
2ANo+PcTeUklLmJOYc/D+4jp9zfxG1yP+HnWOKPGCzUp5rllVFUfMUwJlw5tlxIl
SIMYDP345zXMUT7FGJzluimKfOyF1GiVqy/bKdsKJsKwMC7QEPq7YFHXMWWFRtiq
T6PEhtVrBa1dEuyXI20KbKNlKfEKuykrmTPtExn1ahQwBOdLsRg1KsTemwb0YPW6
VPj0F+ap6jt6pd5Qp1Zz+neeRdeP+upzO4YXFMJxiYBKN3dMA15hGaCnqp7epnKr
rDER+vwN3ho4EGVkkzV+izTPLOokmhwd3jaZqkN4haKCMsE9NZrHgvQ+1Mj8ubCa
KNwLSbGrdHKKcD+F84O8cZcPcZ2XsqRM/DwZXHPM3cl6A0ec3GzKLkgb9QjIdqVJ
fxWfl4B2n9hFqlejqhL04nD+FJdPf6LYMVDrn7tEr/Tz7krZfFSof0mZrjAObp78
E9C6pPGq3hxePUQdfAE83iVS6TBH6CqTo5Hw7uU+7Eh0Jzu8bsTwRGyPu2WJYxut
fK/+cHilMwBIkRI5dTOQ/JyLkznonS5/Cdd8N9sphQGqdGD3eOuGB8I2CcwDnpCe
fa5M6X2U9aIM87L4Zq11hQ75p2yQN7DjsEcEF27JXB6we3c8LM81XRhjKdube1QI
W4JIN+eCAiAGOl6dnf9lUBTXFwiCBUVifqi/b6yvIfed9YPvk/qcjsx4dgoe7i6x
nb/IXKdnsOUa8wkHabl5cl9RoE7K2KqbyKNEslsOY/7QB9Tz9whghRbJzCKj18oB
FFYwbSZF4ao50k6o82TZIcUOGEWXDVLJ4UJ8VdovSzOTS58cQ4BMTvpodMieZPK1
hNzzSmmuZY85M1zQL6rzcs4IFqI9SDavBDBkQoYCJpDgeQmHRE9ZumqbnWlbdEug
GLAm0qrqFiC2A8hufChcQc4FvMCdxoSD5hjdsUmPTT36eI3rgQHaT7jV9eZC9dIj
p2DTX8MFytA56O5SSkOnJvgLFzDM82etnZBPFAjt1HSaJhNhdKBWBg3pETInKzpA
4PP6n/jV+Ywa/sfVeUT847nsLYn5XipiPsIdP0TwXrSdjl4YXqVt8JGjUVJDxFYx
BrfHIFys6rgiTGLpdgCbzIphkf2hgG4Bfc6pwBwkkItkAePhgF/dDNdm8SN+4f7J
K2ZcK3Zu+rxULgyNUbkeSjIDn7W7x2NfxOXYordmIrOwLb81At4PFuwyOjR0MRh1
CHxDwY4aOi8GYx4guT8JQSMPwH897mK+CWazLevvx3QrBzXf8u8BYo4K4BXhzLOo
nQh5CqHSdyhU3QnWCErkc9eN2otrQPekK2RPm0XJ1L2aHPLOzhn+M3OuYOuRwoVY
VUDlT1/sOQiSpbLQODEc5KltYdW+hxLuX237zK+87J0PX6J7iJW5isWBtrfCcZ00
8T5OBR77dvFJ+gmkzD+xmx9ZwDqaEeVDIYgyXCALjSFH/yhexSc4WDuXtMJu36ky
dAPUx5r8B80sceeTEfAowBoRfjCSLSRYGCr+919rs6f+aTdHNW95qDhuCdQNcMQT
xP4jy7wgSRisVkB8yeG+n1nzuTrkwKDtdJJH0ogjuAYnCsUJFvT2DfHdBvOmhHZh
5HQwSPkFTH/J8AVN15S6MZwxMiYxCluYfzWrjtNgxNwPInGMYANBrydlmbCwzpfs
ZLv2Sfwh5iEIbTtYLRLeWYNJIbveSwA4gOO8KWQv719ryTNSxWsFs1HaDpF4sPtl
BfIbER3PWC2P1WRE770w7JA42RVA3wP0nlPpXX59VvIUi0VuxCKz9vClBzwk9O8h
oQ287KDrBfytgNOVF2GcbqulNVGAhoy1jq/sKCA9Uxe3lw9KU5Nf9WmAecEAhTP/
IZvytVEm1G/FswEwJU5KtE6s/qySWwzKeULuj+IOnkfnWpUQ/oNMhkSW9IClUEL9
iwUtbLGgySNBxEym0Kz3YpK5BWJRjx/5Zi3D5KFqJ09hSKHC0zZl0vTarBNlRQ9m
8ZElrUZUxU754nEJjQDX4kJsXDzUq6gUyUJ5Hfu9lZCsS9zszWMzEh4mzJe6h8tq
mxtj7kI5gFAAyYDsywZMwatznmQb5NicGx+cq9DVt+yqb7Dv/8MrYKcv5QJa4sqQ
XSWGmS3Dc+S8PqKs/e3mTQ/+p+pzr4iQp3Eqc3uNJoTzF6HS0WhJsuTxJ3sCKLU/
kLGdQZW4IKgCKubPrrZ9KHw48o3dLORmjHTE+GMCr7t2g+O6jxlrAiEeIocU7WaJ
MnZB5KAqsZUoUob6iCcPS2jkgV7zQOoEuHQCNAziSY4KR7Ir4bbCuWrCAxUY4+xE
d0aDC2/9Lx15YteW1y/0CDKve8H9b0Kg+3V/A27d85WPZWUtPWAZhDg8IkOj0QXu
89ViYTfjdqaNdxBepFKR88UETsqquasOtXxkii+htVGHGkdiloLhps/vJ3rGes4k
fNPp6PHwrkM/TMjhE1LgayELN0KJgCjs5XFN2BowDXTobsdGOytW4ITfdm+iBuvN
K470SiTZ5thYeo32MqXXyoov/20FnfQZZ4xj3SUe9QDXZA8prg/xnQH287b34ipK
JQzCeyPA1v5n+T6xIEHhEjJ1MxatFFYOig5wh1T3CVQOBPNnwtyGeE8Qor8XKg1k
aCZ/TkC39KE/ur02zUZOps4FxKaqxNwtCb1OGphOOPsThJwuRalei6W1LV3YyM/a
86cLvqLZVskql/8sDRYRZPPTbsKv35aCNJ6wP4f2YLlFYXMh0kW62Ce2Q0Yrx3r+
cS5RkP/3DdRE+gWQWpHG3sh/MueXZzcvyU2gzCt4hvVeHtKfBcG38OwZ/t5Uf/XK
LiyvuEFF8+gvXapzDvBjI4pnYgG7QP9g9cBz8Ah4LdLWjd2J9uTfoaRHNpitdvX+
eGv2xP3KL2CXdpKzEDL0aKn8sHzTZiS+1J0o/DiiA982ZdHWBVXgN0AqA41kKllb
uh7RRTIf3dHrU0wblShgiWUY/8qwZcfrRBqKlMha1t0Hmmh5paVxGC5cV2E/Kdd5
633JlRHE2XUGrUg/VaX4kmi5+V5X+3715ZmbvOIhCVqkIOg3bNEC594Lz2KNFT3e
MmL3HI43hfNTS4d9E0HxWqxJL7xLBBPkLcEjfkvHSylWExvhgrOHk6ImcsJqcZPd
Cq3rwMd/BErUB1RIqC4uPxfWMk8VRj7KfJWAKX+Uq27wr9i/Cn5NARVCKWrPzNor
nbPra6dGyJDAyZAbzMoZ0OkFCxvPXMHGvlqIoFqucDnhaQFMyt5SVQS6bogHTcA0
ZNym07B9snyAhUYEUGKMUg+vlBiuprvwqelflpIZgPtCotCFlspNBl7B3Ox/Ijxv
i09qKXG8IeBboAlNBpngAlIMzGslXIMzDX5+nxEih1B0KMkzEJp8v1EudQ4EIH0w
T0vhrGfyvXjOYK4Q1agikiXdc227kK3LkooBI1jevj/RWOtzDGk4lSjh/uX7qBeP
o+8Jdx5FP7pdMIbzW+efEWEZBBOu7JcRCNhi8Q8K0m+KDcLzFVD+vxmqIQ//qNjm
QQ+ThgqZGHR58XRsk8RxK3UZnmGSuWCWYdQ/QgTgFjTpgjChC5qLiYo/5AEvC7GP
By/XGAeU8tc4QJZnoG8kx8CB5zut8H76yHatT/+NxUII7sY2YeEN2g92KB8yCupW
R7P4C6vdG3jnx0zyI+za/JUAvnAb/oYIKKZN+rsN6eURLMAQdqyX+FJd1sqJAZWp
Osqnlctp1skCwR1z0uHu3tw4BqUVY7C0pAwULzUqU8k+oKjqIx0fM9ETZ0vH/gMX
QzMBmlK5ZuOSOZD6Ah3LZ9qB8jqktoECRsk50Ml8/ORPnUFeQ0H3asbUodKJpnB0
vKR4syMPx2xPtp+XsVwnQOJDJSGsCXmWzXZ3fOksr6mpgYfAqx1sZNHnNhoVyFdX
b2c/tDgYVmQ/soMpX7M+XAZdnK+3UtxOdeZge28N1OyQYPNMVfowNL5m19AVyd72
D1jXIE7JA8ipFxWitf/YULOb3en8ZLScfIP3bOMJ504SjKJlahKspVypiCkCkdU8
/k7i8YYZjGJ5cEiThQj1thE+Cvuf7yTesSlhORSKoYR1tcQMRBD4wZUM+Lmrk70P
7f+VUV4tjGqei3cmC9mfrgB4ph2Q3i3etmp0PIfWBZigLGqNTnPt5WAM4vGebaCw
0Tfs1bjGr64BHIYHVee8NjKCL1DxJ7CwBtNjg0NKeSKdYGDdvKaelhfNHT61WGo2
Zddc6o8TXoqHBJdzkQ4dIpjjPZpTfFfo7UCauG+wpA+sxQZ+uulLb4UPZdG/xESG
eP0xASsfZAr2gKGg002c12lPj7GUq7QSMC2Tdmrv4B55yRVKVJfBLeRslrxArluL
wO3LYxEjpGGPM3wZ2PS7Z/2qXlmN8aQRj26bJslflq4x99WgIJrNVd4OsfwJxl74
OxCm37PNJZY3Bjm+w1Cvyhx1STDr9gOfY8EzhqgKOxzzPgh7J1X5DNfaeGQ1R2MY
kr/yj/cua8yPU4MFyC8FV+ng7g7psm8uiS8DSK7kZEeJM0m3RyNeoe4kv7aRM6DK
wdjErr1ReB7tn9Yfuu4SCneI22c59o2IOg/6FnXCV8iDWW1bbJFBuIZRXaO9S3ts
yoN+dPdos/j8iZKwBAPLAej33h9mjIhHpNj77CJFa46JRTnj4odqWYiXdAYE7Ye/
K1OGnCKIciWteljhasvYIOZ9e3ZKKCbfbu4O0naxBN2k7+TZS0uRnK4MUcxn/g3G
VsyUNL4ycZPTxbIvoIJAUDzf0vNUM81xiJlKTZM9FmjatXBiV3ReUDe6QWvrUcej
gpCmUATQPQZtJAIbMed96EamambpmJc7dWcPV/fGdeu0vmEiRLvsm77wOaY9zK55
7klxzLBtfnz/gJn2d6xHyKZXRLVfJwTp+dnBT8TE6SyKOdYfqRnTbqpvrxaWeDFj
UZPDtfFR6tH3IzqvI0sJhqU7TS9NdhFI0aJsC82fh+t1/RSbfG4ENw58bhAAnTYh
DAbI8DnOLKJwXRti3mzudfqdmfVu/ZT7sZKlJn6J0yTz6PVkLdOWQfC7OZSGbSeM
2dw/TdbZL/EfIqv49xnrWdqUDvNcWUNFPajFGwadtzvfJoDdyB9G13eE1G6lyuAQ
2dfjxT3fz2Y0jCJtv8rGbZxjYlY5PwL9y6G/VQdX0ubi/ibPG8+9tPp+iw0SLqDB
2A2dVnMG788ANWkQr41IkrIKwy3Tm6f9dnmKnh8ZnNalIKEvg2YrgdzLJhUubmcX
HUhJHDYVbCYI6uVJYR+UZtnNTQV/anVyxlP0dcV+68LtWmPhuaZYKhY5HX7TQpJi
9biMSNwtHHu7ch61tVV5Ubf0A1SawqWheum94T3HcxIbgglLsa7jiQmmNwh6K/t4
xk6I8/DaI3oAeAS0/u68tgZGEBP6+PPfcyTlEAAZOnWfBYKlG+pF5fcKye9r4Ny+
2880n/ps1cbTTNd7yb+lAtj5xZDErnhID07qvt+O8dU5T7yj3hPICG42xjKDvkuL
kwYwWKn7sKFgDQPBpt8NJbi1C5ue/ad225WNYWEKtFjD18amfCdLBtKAwQ3og0P2
jdkEUJBiF6uS4PNW1tSZ2tfgkpC96d+EDfrISeXSH35fAxTUTIqvVR52WEzwCLXu
4ePl51XCqpt1XfJ9zXkZx+8q8ZzM20uinR8QM+Ah5UdICCVbSI85NDrv6jp9DZ4X
fxzr+7J5wCjYX39vTREPWsO1DvxWcXUwGwqtxF+V0nnjUlQMzVSElV+C3GJvHW6z
Ulv/baqRi0RsrZrTO9JruWQ22RKdQyMlJogMcj4qZYzym5YLa2xcY8NCgOhaTaZL
CyT1yNPIUDARzzC3lKMieg01pYoSq6/IFaaqyRkuBMjj0VEqJHuAVAh0KPG/XzJp
umaHJ9BAQKyYoARZwhkeRjh/pEuj8mphF6ejKdbFJFob9uDeAqcUacxBAnYkTuKA
`protect END_PROTECTED
