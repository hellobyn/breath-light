`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUAPs7BDDoJfHYiTc3zOy6+4I78rcXm100xWJ77JxJNsk8/QePyEidD8oR0k2ArU
9RbOL15p5/dOHaNi9rg+mSFiWRqJHDCnckQaQyi4loiWfvX9lyjcL7GcnPEXAKnc
raBElIH5sOTF4g08GgwDtD+nKKv+JoCBDomNZhBAoOsTqAUQpYTB7z8DmT7NmybL
AX4QdOepGklfCDm4qULVb3bmQzoDteVXnF0MYiAoq47FG3VbmDT8TDNOgCxIEvnu
SLy6iC6GUnLsEgTlcYk1XDtGHCG8gOqQLyugftD/9i5jqJg4vV0M2twKjN0hcQqf
4xY2ARtTczRRD9Sh0Ai/PYG6BUDyHgBMJ9id1pA5jDkzTBj8NA7YQh69HJ1UaMAZ
I5inuy79RmMkyzgx/U1Yv7BH2uhtI0JeKg79DQ4VXw3xF8j4ru3PbZaWBYWdGj0G
5Ol5/mrvA8xgpGBJDAsqKL08F372xxeHtr+l8DafQXVNpcvL1T0RZQ/xVekwr6Yk
Vk3xu71VIxlJ6N3xUCO2yMSsr4emAoHu5hFREbKCWLKFm3T0gwF1y7yqyhd/Lc82
b7LJnhYv6L0Cx+aUBis4evyYYNBAYH/ZNLoDbettZ4WzZ6oGDlyom16ZL5bLl9WA
avVolND1dLlu3REBDom5LJ0R+/YxOjP9PXZB+JRHXZXcLgkF5AAirXlAAci6RAFT
y7Lb+mdelkQ07maiZpIhHwxLFhgI0OcY6Y+Ue/CC4ApT6egxw4RTOA6mK96WjKIf
dZy1Z+LgayKppg3lL9O9pXnswK4Sq09p3PtSRXWY3F+sK06ptApNNeD8kDSm3d++
RV2/WkfGkemhyCXo+N9KOg1+b+4xZmfwTFBhA0isnuNhLnZjgPLE24BIKXAN2KZX
5WHyLiPRpoiZ/L+G7WKa2HuvI8uTDAFxh3VdgCf1CMLgdbnXJJT119wDylIejWvo
LnLJdg/LVTAQJ8ifTqg/w2aFE9jahh0Vfh4wMvTBfiwAXFINMzXjKYtqF8Dv65fc
/olyhDbp7SjBnsQtBdFUrPjMydHGDrdjBUgfRsIojwpeJLDMVyIHON9rXvTwQfsr
GYgqQ9+puylCNW7Uz1CXQWzx9ScI9zwkThum4f6kqNciZnCwLssalFaeblN5aXyf
3BjPu2gvWnhIba//3cigdYNwuSLtc85zgR5W+QVTQiiVegx2D48vluavanPeQCjq
ujvwhPRGo+3/BIGlBDT+LQct6HQFuRb9qXqC5B+DB6IQg202tY/hzZGystYYCaPw
DNCZHTogpPXdwMX8eVlN0OlUtWGZswHdZvAOc3wZmL6FT8WN4BrZkCK2afhcvSg6
kNk5wEWqaMcvuYGdrHW9+CZKjkequhZGOa4hpCdLMTskJxVMoYdUSci8vymEbMoj
VFECx6k+Z/6OmotM5SWTNKh7h2NeTDTt5JCOBs/8EgLVRZCo96u9c+LL+5h457Cw
CRKWk+9PjnBI08gfqSsxrMGdOTjWZcIjXD9JFHCgrDxHluT61aG4nkehb4CJ5KKd
VRrSi7OngOSPMg1dOJEeSVZWrpiJ/J6WU1ZB/ZeKC1ffQ/J2lWX79Ub407DeKyhX
Z5bpVfvGUcLIvNhktN4EAE0LTcngmw4Sw+MubDBCIgfxm26p/bLK7DYWp9t4YzWf
9MeOiaxivPTu5pqKP1zeV443RSBMaptpFdZB8uBK+BGUz/N6pO5KNomGm4CUYDmi
ElFPMXwFCd513KjChRrqbuzCWQrYIj0Ay2ATKmzkkjMXvFV1X47/JwL9BoufOe+6
TzkJpilHUCk1gva0IWrRIl+ybOR0yhiCXhDpcU111fb5pDLvISNXjdeX7iAdo7ev
P+pkpOPmupwDQgHVpF9eIu0WiLovQgy4jXeKreXpMh/dcqOS+jBUJXQcmO4sYBLV
G/ycxAYHZUb9GbaLarSTR0xUdkKjoR6YaOxJaoN+6AaR5I/dpB3IgFJ4Dd6mZHRQ
yPSUD8Q7mlkkl6YaIsGIFwGcnC4MnrEba36LXF+ambCcPDMOldpjfm0PZbq2KroB
3+XG4zCng/qygoPkc3GrJ4j58uBTvHCNaofyv3yT3RMigcitZnimqYc1gQK3R2wl
fqDEnUiWBNuGmbfm6mjpCaUY577OB5VY7lm2wY5DXbjBjNg2lhafLaBp0YzFHYVB
DG4scRe1wi72r0C1l3H7xLlilSm64caHLNS1CrzQ6b+y10Yu05h1+DW1g7b0d4jF
uaIcHrb7VMhSuWx2PX2Tc9LkPIkhcnHq43Qa2VaLjNxnkmwUvTCqSUKDhePvjnsq
OKXEeyDfzXfzb9FEv7yaYs8NDPJg+lGbirYep4W81jd5vJ5O653gYR/kv3CMWnxz
SjK1KGGPITZbFzMvvNMT3LlRdYbpawzhE3MxcItkJHd0PXrTPbiby+6S+lRFrk9r
yldldyYqJfruZNj7PW/Sr8HIzjleO4Vu1pMJEYwTQ+TOzBgSsherrt2v0/l6aH7R
Y+R7gx1b+aIRSmsm84FF0c/2TypxB+j13mO8DTc7CtjQGKbFcuwTmnhYpzlajxTH
S6AKxa3Ym20qzaLjODoiGOh2P/ckta8UnsSeAAqFLMwmmNPN92Pz2Jla+FiZlzLJ
FihidSS5scbYy2zI1pzEn/r7kc7rmThJgRrnhpdqcKWLk3y4Cvu2aOGnoSu/Icqe
qna4cxxY+Qxfkjj6jmOTjVH7ubHwFHOA56Sd6w7ArV31VMX0qQTG8Bz8xP3uy2Mt
IKO+4OzBCQukgkNQ6xtFPuMSrbmEJJfqFS/ZNWuDfdboO5sbJ+mB8OqEuN+Cezxe
lM1c3jLydeLEL8UOWDPwFI1+cEh71eTJywcaHepgrRGnYo6LxGT3yqq62SGvXZKQ
iOlCRqSQ5HxXK5En3EDtNyKaDeFVypLV6t3vEIejRCvq4eQyKsulDJLpUAvCXdUD
W5an+4CZEGOxJ/FaqYCS/rlwRYT/1PZM26MmMBdPketNfMzAwW0ub1m8uzKyElwo
khK2phNjU4SKNiE7VDO+k3sLFW3WwXVSgJSQ6TngRdvfaCQg77eUMKhHwukyR/8H
VJ7aqGXMQadNnPaxtbR3f3q4glBKfRpDK8ACRykiJ6DGmdlAeg/uNqxURgwehaOy
WqUa7Ql7QRJDXECvTALZm6ja2Oi3oekaGPY8cOSUnmrROawBr6ReUp1x/sWEvD/J
Y9Qd4YqPJJu+c62Alatukg==
`protect END_PROTECTED
