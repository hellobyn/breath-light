`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yzpSar9x0Lo2RMlSTRy3O3d3Tq76ZjK3XtJ2kxLQkRSFnDSpkCECYPQYT4kaHo1
HgnxFvVvnY0UjuGtq1vWXgjGMVe13gFwSn9M+RPSzxHT4oqEFfPdvyD9Z8pByaw5
IYy8fdxBW7a6PXCn8FLTHhfjiV+cqBKMa1juE+xjCOorX87+ch5MTvU2V6DrLT6s
BaBQ4o7OT0O++pGpj3/IH/KxJIIg3t3ba0zd5Gz7Ml9JoGNracOzBiynfCbO4DJR
fQ9zdW+Q4GfiIexzUrJSYHpeyvqzvq9PFtREqHb+dz6CMrGe7I0XA5t4u8Hy+1Xb
7q3ZOStPMMb77PDBGBCzr013/lSs/dusAahLDn9dFJbX3BGoKQ6JaXELCQdf1ATt
N9Ix4oi/Lq1sfLSH1PGm/wEkYKl1ZysOMSjUiboriSci++BzyBFgbICLB6CSN73z
MsLIlbCND/az47Hxy4yOYPWoRCnVqZ7P4BVzTuQIXQn3WZEFhsvHBPbM9qrdV43Y
32xbvL6GREmcIZyZaf8bahTFcUE69ifyfMlJX8xTj898tEuWr292+4gi43IKloOh
E2KpXykj8ywBL8plqLjXpfdgioYS5AVO0ycsTLe3aHSm6Q8XW/wEYJyUyIXfd+RP
pJVO+pDBXmLDH7hHXZ+WDAcBU+xhWPZRIcm8TZLBsIltU+gBBAXHeKUo8iNfpn+d
XE2tZOJMAy8jy8pfjtxaT0ArM7jIVn18HVVWDrGpjd3cr419ksPVyEMx4hZVa2lK
t8Dd9HdomjWFKjA34FELfw==
`protect END_PROTECTED
