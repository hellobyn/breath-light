`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYMY9IjO1oEh+Y0i3IJjgOFfW35K7d1sXZvj6cTqRJpzMY/J0VIuDijSxJwCXREW
HXg5Tb9sf1Nm1Q3QZTyTv9YwmjCgZKBQQua2QOmXyvaD2kynSg1S3MBaHK8hgw8a
ONV3tDhuWqyIeeu5GaFH43qlXioXeHOMsVyOjxAtEPRknjxzaun3AG/uaLOv3fUn
Pd9+ECTj09fICrRTTSzpa/wDRR+ydNCpdWC6lgQ8751MU8CLp2v8ua31YgSdWwH/
8TDKxKppD2VpdDkY0AzF8GeWWzgEPG0zlVxdwZS+y9jJiy/39f7t/gmDhNQ5/jDn
l4nP/0DQWbKbbofWYDMVxw4eDSw8LTMX97Myu+eU1wOAX32Mr2cE1YPxtG1MVTVP
f0dub6JJFDCvNVjW2dCTbpKqAkORoatJHq0prkPXtCzrJi8rSGzrrjeabj0F6LTj
K+tOocl9LWTPuK2ffG7PD153ksNELacV0w0h805D/NrW8OHHx/95bBsrO8cKp9Jg
QD8SN2UsmfaXj/iva8EfKsNkJ4/nlHy4GrMPucU5oEOpKQsNU+Pn/Be3OsGuWDkV
H4QNDBj202suAA2QHlLpGkMuXcUVaMiphz9AQiFKCsPvuBxYFmE9xAcwzuHhOHyb
IrULOiY7PCDqyEn5XH3GNP/Q5sDswD1v4XSFJIcqM+hTB2GRYOK5PF72F7SFv/Mh
Y5n/n0THotc/aHeDrObURyQhcGVsP3E0i+1o+RJy07+7YkvnNCrKbnNQlqWeoy4r
Lbyyzl0niz1/arIXvkbVrnQ9KO+NDjpCWr7qguTjeiyiC0LKiKoFXI798f0U8NlV
i2yPrCyITbtCOEDWvk75V10pBIeOVYE04UqVmKgjKG17NCfYZbJAdueuhsK3PxGb
yS0om2Tid28Fut6BtsLO5G1u2PXHc8Tnsn7ixRXPV4heEzEWvqJr1V3EPcRcsJI+
f13EJNhkDIWWeXqe8PFP8RYFO58lEvcIiJtJq2AmAuTgsy83K66ArMtMrliMGYU4
geu1tV7ASNC14ER/lLDeLRzx/Vl8LHJlMYkkAZNINkVbap49vUd54iAJ5kAAOCTp
wFglhtr++nxKTBU+Hjp+vA==
`protect END_PROTECTED
