`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9HxJYo5siy87Qk+I2Y8qTFiVazuz5MBB9gDSBRQKZUvkz+64Jw7yqHQFJamg1sF
4UIwv+ngvRb+hi8BLSbpkkH95MqIcVOWilBriykNMf/VwJL3z7yt9eOBu7UlTESb
IXymSG12E1Nn7ZcGuqG/ehveWiRsi352ywit9K8dNDW7pr86yRo+axlfhalBKOz+
JlLAhRiqn8rlK7O8P6nlkgrmAJT/wpAjdrgj67rVI6aXgV3ae8ZSepH7v7XlYwoS
ZFW9aHPwGJ6XigEqJ8za6BL+r+hCZadyQ0GB/EmqAViEfWYRplxvJg90Mv3G3Tyb
OxjIEYMX17dhh7fv05AoKn0fLiuCkNHlsGfYmk3IMPr1g2XIKPXYt3ftOL43PmfP
P079FzWKfjxhT9HzKciHR6j7lo5Vpe0ZGTYwVV8aUY8WtvmmO41g8UJ3fUyERwir
xAxdHj71QkAYxZbmXMR54ucJqm7udxf3zWO4r0+k8qom62TK2R6iPn6nuXCROs1P
vrnG4xWcdgZEdUT3A9HN6m3ZBUVKIPJWDVh/CByNRPsvDNAiCyeNlHQORtfoi278
tFmYAi9GEsGJk/s2chxFIvOJSZNOqvcGUXtnh62Gud37pRauC91uKha1LQOJGmMI
/LbweGFCL3ty6H9dlpzw8RAyQjmY8BD+L/R9Uw5AzTrozIS4Kq9I9O+C43NDoMJJ
SsHC9+XSzupPxt2ZxASp86XojmgXBjrr5ttlclVt3IGUxb4gta+WNpD0njd7C6l8
riQW7hLsWchiweLG+fPxaXQpaZ1ByHAtIPDJ/aqFyVQI59itwJj9tRdlDVAVps7I
fmh2MoMZIRqXjTnX0RiycebvjeJH+l41Nt+P8HtHka8YMFYcgpR074IJ4ju4VZlz
j3sdLDEleQinyZ8mbEXnth36Sp5R2VrZSMT2qFfdMWOxHewWxlsxSTPfQQxj/Ea0
icaUx5Xxmc76VdLQTumn31ojHae6wZILvIAS+IN4biFAfxcDNPldDBE6yneK+MCi
9MngywpWybRyEOXgJ7XE8DbODWuieGbnIYl30WeEVV7mDLvVL33FlWATU+swx3oD
svjc5fIWUjIhRcsj9Yd5c1A+kPC7TOZTC0fetg/yGaymmrLGPX3Jig7d/UfztvS5
/Mk3HitbyaKdEtsCjSc7hIvuWMEObUqi2gQrv9l31qBPRbX+Zi3Of27tc9u3F2M1
Y6J+zzdvqLUZNATuU6Y/YiRVq+w18pkLG0BR1ulVmTrCOmE7bSIJQTL3yI5pHiSs
Nr3kzlEG3bZda/wy4oLjeAiktp3xtRRSLafxVaM6bO1S9xGvrCj+a8PnUny9CMis
KURKPXCgwV+szs3MUlxxJnRyWctoJ5yTLZgOpVRqIsSlLkDw7zMl6SoY0w+Tr9Lj
zUuLisZ0aQF+duwMIdjR496QerVpOkctg/CNhJUMGEgUWEAlrbzBLAjbFqJTnAK2
chodKtrk4CAUl1kgZxc8ZkiwHv+ka8Jr7LLXSHx728Z1mTyJaa9cHqoihOuGn3yq
p4rpOJkAXOBfqHSK11ndckojI6Gj3jcGXSbiss4vIbyJBO123cpiDsEXRGtmJY3Q
GSC03eUdNHh3/2i8Yu+ENc8iincgEd6VCi5V+dg/7Ir0mL1UUT0/tRn7wSo5Ajwp
HiSX/MgEoGR8ldtCEbmoUOU60WioyZ70rHWHr5EnhrH0GuqHfyDcL3qKSbNPrbsy
WVh+5/2UradIoLyFjLzQ0jbQAr3vS4yLipwzjQYNHwg01zjA/nRKDydim9/Cwhoz
v3hn65NF6HpUm025CEJVMSN71jdgsJG4rFRI7WtY/TmXf2jJwva+P2/b9LSxkjcJ
orEMuHr8igLjyc0iq9q9OguEPAiBQlEIFHzqP9gJvQnJJVcLMHDxtYZGbkwh2hd2
nsYfo7q+8guq1QgM3koJ/NtTnp6Vw4658RpPhJpQnLw5ad/krkHOpbs54k0Ctt+z
C90GLrRo/vHoDLVm7LzK0f3yJidY+c+35Y71eow2Dduqa2Iy3KL8zs0OA3YOB32K
EYl6ptUJrVu42MJ0YnQ+s1YGkBMzMn/jeXrhl69aeIL/zKCwGjcWZwNrhJl7XymN
0X05iBxDFS1+lGJtjTaM6dJZYn3pZIMoZNQPaeJw/c+fHuKaf7ldpcQM19LvMyK+
9SoDkrzjWZ0nzj8MKbFsUFg3Nydkukabcsm2fBbfYJlDIpySEfIj4MC+ID812fEl
akkzcdwLSkH4Y+NBo6zvD0fe7RHjNY1qfZGthlQWALN7xkKGpi65FX+kCaW/0O5B
QN7SaviVfMWXPMi/cN3BTUtgcPSIr1H2/ZlDefiXXtE9srHrqTs7wn2VHC3+xLks
e1HL7fBkq/lx465NeTCSqPAnSy7fIYzODQdXroZ8IT81r3mPu4h9DwiXTd0Qv1+O
egvbv7Mr7B0qFJD9TTceUL4U0NyJNDGbD8sBU55fJKV9EdSP2XbtCxpsJDrPFpfE
Gn/x1iEfhmr6AWbgOLsS6xIperTiOuYkl7jcNHs4bobQnsDKuiOqMiGGFBMzgEP8
w+EGANpX9eWijNlGtQI0y49ozxhxCsVISpK8uVE9VV71VD/P57MzoghatcLxhBvA
IwTLOBjkHuqbSB0e5K2TtxbR0+sgOdHN49fD/1LfQqYT/4qFWn4y5NXafgRWiwah
pl3saIfHVOUin937k3vbSwfYkB28fg7/1wakwMTg+dkCye1TfsxuDxch+6kdi/u4
MrsJw2G8eQQUmld7KTN9leSTC5rTxtBA/1gvuwy9PJYEBMQ9zsPzGDITYJwrfQxp
n3MFyyx7AaiOIAVIiobCccVIXE/hGvJ6XIyzQzAUbXDeX0p6Bf9qyGqjG9KOFZAB
R/TMHtfx/zLyBYAVSFHplwKSVFEuymNJ5pSyvFrpMgtrNyDGP7IeTuGfHwtla+zT
enonuuOG6E2UWGb7dnZzts5Hb1v10nnQNvfyRwGa2ohH6nV+8sfjA643X10CYaxr
KajuD6jU5ZAvIeekBYZzeeOoYXQLeAFBEVfq0p14npii/u7oaRMAnNp/kBpuq++Z
nCOjwqICVWyu0ORF1y/UobUHqTb//hmOQXZScXVk1743nGms5diVqqjPDcrcAnLp
RKpt/+3oPe6s05YokKjzKjjaR2texunVuM3VXoW8J10aeSIcHNhe5wC3udIA6RpI
7aeOK/SlZhTwF+6sQlc41pZookkk95TuyEDMRjc1hiuagRghafM/2yb2owe25QCU
NpfQCbmMnpYbofqqpzElJjoMIldwHNMsyvwBHJ1o3hes0PwYSQAJBjwIaxF0sr63
3p7iPSqBTpapTxbzzK/BWk9RDOv1z17zPe0D6niiFsK0r47/PmCuGOznKPNPkGkq
MJ8Jc6G6BGe3RNx9Y/EIELE/nWO+I33HcMPcNmcjjP5xpdrzr/RzP/dBh6BehV5u
ju9SdjsYNl49lZ9eTyFFh/aoIt+yt567wJtMUULwi7jVORL6xQY57a3YYhkAtbG1
Ik4JbJ/bSr3FLRdbfw+rdvEuVNPS6QXKtTULiwiyeQ+Wp+hy+K/w3halpfSRv9vY
Mz26V2vbtg8iRejtjOkAJvhKv0ep5K84eQbkMuQ6tWOjlenj4U69vlFLhiFjqofy
8rNQWulAi+QG1lqPBo4rXigg0juVDrbOA6bwE6nxYy9EthY5bB3kMEYrlGOdSoG/
w51jorRumHHFBsoc7R3MPTjb5jKl4MBICnq1yPPkPG1uM4lwngRT+mTMGhWytHqL
bn3GebWUKHVNZK3rw8om/XbNA8xHZmpD++pTU597cBVUtdhbeUdDluNzUSisbTu7
mIclfAGFi++ct8woZVjJYn596POO3nE7p32uyPCVgxjrIQ8wHrohYqhRRIAfpcPR
WBRlDEF4yXVnm+XtVa9uukZ0aXlwFbuqiBS80abY5z/Y2BAngmmvNsvgXEkw0crq
TSOvsgWxKNeqxg9r00lzMTctCtYTRSMKZ0uGx7CiX0AzS4v2hfrrjdqV8YCowRS2
svQcpbbWC0pLhF7/qlr48ZKzIaIZYk8BnTFvCLBsliToJoxjYE+JwXxpzHlaWrKb
jhE91HsNX6GUkMix13raHapXOzWrpE3bhklVEFKQtzeSsLyv8+xwqQIbxRb9mt9U
vWHtRK0n7IeYtPKg3paG23kY4OxJ67a9NlDv5Bn/E7ifs280xPfXWTu/Tq7pLr6s
phrtNcF/PmbKXtqeaOkQyG3OuIJ2oZOt3aZtUmBG8ISDjToC2Jdrgz2Esjd+sqmu
`protect END_PROTECTED
