`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4akwlj16Hp82WRQL10/jt9wcqNL7tEEiX40mFRwsilwUn7uNvhQvGbrZeZpuadg0
MYfjF6bM8phpIO2VKC2NWrOhAXQy6Q/6U8qVd30qZ0az5b4bAqoQS1izjgD27/Sh
z4XjK9ShnUrw2+flLia/pdExLBo5qvQfon0SsT5TQVjrxr89QwsXsbz1ASonge2x
/UeWGzJGn9RQCl5TxDmmLKPr0/SqRG/2BRyr8ZW5ut1et114l1zPTyB4kVIrDMDH
BwGjhb8fo2775xxGE9Yon4tMwZ3xzkpUazHca5otdzHZLswww3BupHS4+zonPNcw
5VmWSHAWFZRbU5eiUG7sz7+3B6Wy+0cJFTPBxmxL2kna/KFslw5hBI+4yaeOXq0E
RBQiBmNKAchGWLUoQHrQFhOucocOVdsGg+wl2UPzuScy6iiSfbmWsCQWFMGN7mrv
tBhy4b6yNgqwhenNjNJZaJ7d+z8y0qsRn+gfXV8U+xesIgBlik/fBET3E3+ZTwXT
jD9WbyHRg4BhToMpt1TFTusr3NKEwiRMgtn0ujwlwRUxKXDdp5iG6qcp3IYVXP7n
w89Yd+uEif+su5HBpA2h3VWeRfVerKvQTLL4jtCgay5TLjljKaq/2r/uPEjGdO8N
y063IondbXz6+bWl4LdDoK4bh+88THSQAUrEJAH5+9APgNn5Y+4oH3E9b+nTu7+H
f7D+SuImGpcvoc9e7ie7rnojxYH/cejT6CMhZV3T/SGgmJIyzpYQt+VOGBg19OQe
cg01D+gJtXEjehbxGCQDfa2sCLnitbjTiFDkP7NKOEe64izZ+Ir/nH09XvKnJiy1
BEY3B++Fr0AqhH/8f1r6DxeX0g+sRO/i+FTKjRMjiXxLqSIxm6jv3ov5oDeqhSJP
g7coZcO9Ry2SlYnjjw890ye6kBre0dcftQR2amyLMs9lUX7mq997F693ArcE9hcY
ZlImUPh//DVO/VsJLUKmyA3BxRJsyvbQramXQLXQryG9f9vygMRNa2p65znNR6xO
JGrkRQ6aHLpZ6TEnVJGJZsClrOYaRcm4x1msTbQKN6yuyRjEO63f9VbVld3xf5Ag
dl8S/p8wM3RPJf+EIuc545/HueaijKhNrm+mOKJaE37Z51OHeU3JGBxBpnzbx81+
HKlhyUqd+lzV+eU6RgfPlye0g7zsFu7NmKZpi5qhiqNNDw3IP8kpjN3lUYATtANT
xg3stVkt/0Fu2PJQGbSMNzVxu7NExo7DeaGzZ4YHRPgJwIGZmCzUp7pXOjJGSMQT
IvlFdqJ1Cdl1ZUvypJo2UtiO7hVYfnd31C5XIn4IxtR7Fj+qEpHJdPN7+tFrB2GC
zeiUJEXJVCh87ZM5adBvQJastgesXSelRLyjZs95D+G+tVxmtzZQW1jNcx0qhN9Z
yXqEak8wnaBzQJYC4dptbRSUPXRfQrgF7CN7Nxz+TSouLsiiLH9rS6nUTe+rgRaH
B/ryMkOkJurD3YFLidRCFqEZYUmTz56TW6Fe39lvBvq3iksccX9S8vD3DpDy6Xk8
2IgZq0ggW7I72+g+NdS/YY8f3M9neVVa8aD9LGUsVGIQyfb5dECCnH4UpWaMBSoK
H4CZSD1mPgmRbR+eD44rLvIyCAqnX+fo33dhDkDVGeqyNQ7cE287DmOOvCe+lkAF
aprDbG9elLcHTxj1Z7oSshvJr8dW9PcpoRCqzVG4ip6nZVjNdu9y4f5VMNMRe6Yt
fA+dh66GZbDTG+B3w00Jk8P3amOGHB/3s2HW6PgB0IiCs/p+2h3KQAw1ziGnsHB9
5pCr2Cl2sMJxflZx02ocNSHv54qY2Gvivjk9tUG0SQXFszO5q1Ntfz37MWPCCJwy
0Y2tN7sE41lL4Q6V4IBH30V2r2Z91TJ8FcOhZyK5cShch++74OBvVcZZ6awUU7SE
HCBl5HZ/5+uQZeJgIKOcLUeZzIVcaztoxndBfMFk6pSmtGD/5zp7t/TxNC9TuNO/
eL2Vv/BsZWdWH2FpCoLlRkvJ4EmlV4n4G+RcXkG0dZ+yU15rSP8NA+LZnceHCv3w
4JRdbsYjvchrcC18CcFC3l3gZ6k7RJbSVnOaoAgfXK2UKpR1RnwmsjLM35+qN7R+
6svSEvL3n59arf/yyBokUTvFisAMYr+5p7ERmwvU5QzpP956pmPH0qZ6dj2XqTl2
ZSOGkKnaZqxdNSDGJmArdNvUtsK3dtWIhYpEGTiVchRgPwA4oGIgZftVvGsMgxcL
S6E6+TW2cWXQrLuZDBc3pQCfBtVeBDVwA9fh23eP6SUyP0wK4zzOE77GboI+5q3w
/9D04f2UTLWqRVARGYtjKouUHmBnYA7CWxFbsuz3jJJ5A/Z34Sq3SUkbX61gON97
4N0bqAOtXaO+mqo5bD+O8DsThsoSKPiLXCLEuHeSAxSHYq1MRm9x/TycKeR9QJSF
Z9tMXGngVxM1AHOlmipTLSau+jO5MEgzuL4+UZbTvOWdaaxwjEhuwhQFW6usD0CL
83bIM5Ni2Gix/fFY/IP4WALMpmW3WEJ9Atjc8lVf90nM87RX2PwUvl75fM892WN6
WefUr287g6LnsRO62yuPux5ymwbGV4HAqY15VKUZsgQtbA+c7KT41VyF65M60IVb
M4PZxpthmyXK4mYxAhK1rYIKffKd0twZEf71SDu5qGBRsSmJdc7EOn5hzjroMGK0
x2inzEzAQqffIFb1H81zkrjJgQDwl4fJ58EG/bQ91u4uVN4/GCSm0NE5c5KVuIpP
Kbr1idRvs8uj4ej/Fv6LqPYaAI4kSij6dJReXIO1W6BepKc87P+m7PTqcMa+bf4t
k9kGbn3F+PHQXdrkXRW+xaTgxo0xzJ41Tr8X1r9/fjPZzdvxEonJDiOhgNyXaMvG
1PFWtMr6NQQ1Pk0ed6+ltrGMm/y9yNWT5oL+Fmwu6dToK7/5/5bfBKDM6lZiZx7d
2LspS1kZBscr9rhsoVPS0KJYBJrWkmnH3f30fAptiLbIFSe7irooHwgtjfS4Ql0M
afjTF5N2YeyTZvkXherF2m9+d3iv4ehhKuav2EFbhZ2AGyLFDUYcZuwGvFbDBnhx
nnozn4w6hRrssFL/DqTPUSWGQOe+/EEFEVa4OZwbNS9hfRU/b6+9VfYPLGStIew7
unj4SIC1BIY6hnLAkqn8voCgoWSDKLva5Rse4dmfCtVxHLHineoAD3o0zWHeAbiW
GS8lP9JTVYCn8gzTg/nOnEbDske93F0frvPRNSrXC7Ke7a8kqEvGS7T35Y5C/GPa
ROnQ9MkWXxChKl5Ovh/UuS9L0e5/lV2zLFPZTsns1mHL964UkZzujTpasgRGMUcr
SY789hZlQQ/bR3cglaBsYBGXD4/RqukEhR0IC6Ag1au8I85JFXa3/J7YJI0a0374
KmN83FqBQcx5ZlAHqiiy1PP7xZgBtTulMb3fyPvt0espmpftMeCj0qTfHKXfHlfA
i9tOxvKbYuQvOfvfu3OEh/0OZA3FQyMt4HbVGOnhmgEXNvbT+3GA5waOq/2Iqalz
MgmzvR/4Gxr/6+o+yOeVSuGfKXnZ0W+uKFqmSXKxgf0wDbhXP+5ZA1qX4x8HlvdM
p20EIqiXfo9KwVzvjTKiu33ynjzeF8ER7p7TMaASfbpG4nCuC0hvrwNZgu3ZeMr0
3pz7bT1t3ua5F59/wM3lBPQJWKN8UhXtLXL9QzlGRrWmdReYMxyvmhMNoOzqSpJ5
dJ40+dv4cKYEe+NNvPJ3EjtTZ3jNXI+YLHsSy4BrifwXh6SF0SLOx7VrMTZd4Fga
/KpAucX4xax9RBrAyIWltrkSakoRyRcnWts+whj0HTNf6Xt8GBG4LZ+RVphAPa2F
1anQiq7wVWC9Cnn47p+kOdti+zb1qWMtoMtlr6//WmWOKHLvIEN388nv/qtehXLz
a+sw2THml2ORzCzqw0WgbBiYrwsw4kRpJEmVoM0cvD7vVZ8TQVq0tLTyIaluoxK5
tG5W6Bbk2meW9uniTSbOmiRxEZAD0NY63AZS+ZCM6VjB9Ng1zrmfPwJ/z3gTAyZ6
boAHaazhHJvJ3bkUg4CgR8TD0GpKncHRqYw3L7y8Dr+NVT+6yyS0Fyl2SD9FuJw/
rL1PD9sBzNVE/4MvtFtFlGjHXYgPWLIJDPoYiNgHIIXHErP0vg6OOeY6MFZwAWhK
5vqdfZ25swLfZKhChNM0a2Sml9+4ebR8aztT/ZIAm/vCxy4uw5IRqUud85fYBkie
1AXVtbCXbQ3cS6VDhcJShm5kXi+4hFwXpBk51ZC2Z4A7IPfQF+FAIVuXpUTiyG4n
VBwss2cADJAZrGu92HA4fQAUKN/Srdcu4fLlN3fCw+Uyp8Hd2sjtWZB9Cexo1gJS
2cEyzMJCJHvtDIENOaLpo4DNh1dciqwgbxRt99anmKDBYsPgNpeJLmou5V3hUFNS
gQafqqjfRl1qfugcd2tpC+JyyEF1ifzn8qmQsdpPXBpNpVwnLxhG5S35QqzDHnpo
Kcyhgg8ClKiux84/nHuYWbXpq1+BzE8YR56XEfveYjW04v9Cs557lD4gzVTuhCap
S9PyoNi1NkjK2OOUV5poolL6UJVTOUiN+yOo/3k6wtuCOhchcOhPxWX9BwBag6qP
pFFhno2egNkDMAagBLHWcG82X9H4sC267b7PuXsytrdlrJxI80OQ5vmXVbC+A9PQ
KBc/VCeGWCKAj6bZW3fUsdG4pckpIlvNJkwHB3yTYmKs4cKrjZ/o2Zaa/Wgr8HwJ
Qy0Jlt3W4zqXdhJctEbTI9pw9l2fGsU1Ho5B5cC85MZ45X5tIqJGANBjARqNkQ3u
zJP4QtcDFD4t/nPIK1xg3njBYeGXRPAl0EnYqKAqLYnpwX4GBq/r/CDG3oWhhVLv
bIOwWvBoTIUomC1mTyfA+W2Z09XUin1uEqn6m12h4ctyu4XT2THRwamIkm3OvWdp
KSzbd/JyKZBIaK0tlOeOFxZ0gmxX2hi7GsGVpIqKD9VgZXHItI21PB2D27Nx9ngA
Pg6wXl6osvVpXNjA3HVlc8PZUIv1zXPH2XUCMX1tvFKRAKPtdTcOdMbr+QtCRsdy
gblTQCyIoY7RtOkmvbH4UQc8FQQEwte4yjD2WVoTg448JW9WiGyOifO47RwRGC5V
wbbKFpFBfglA5++SNTLnN/1orOnYs/TeFNCR1imNqodrB2PYl1J9Ctf5ZwgqM0u4
H1ceThWdwNX5FDWS3OgD8wvCxzhpOit2pWH5SoIYgkHmBYXVgLRJsYfFwE7BArVG
Cj9UUZtJoDtg0x/9ifOdspX2fqMDeH1WYvUO2B0Tn+QCIBGcHHBWzMTCJ5sVto+z
6a1/xY3ZutYb5oF8r+1jN4fe8s7j/nAK9x8RlnBoqCq8MxgkCRRIM1acvFrbaf0n
obT7JVAUF6hWc5IUFGl2fiXCh6SdMPnZUOrQ7L+HQwwaq9G5iunoAKTtJT3hRqr6
14M+fzwaMsKLXbSOmx1XiugbXhdl/76u9QQmHiLakoFA1ECrS6JrAF782D6d+92T
U8amSUfJJIvUl+n1EaqayRx3Uu2SoIaVX61WMik3Of57rRoH0vLTJrJgpMEmgyxz
54A1JWQA8D9fK5n4Oxy03Ewr+730/O7q86IWdEc3cfxJqfJf+evM0ANIbHzxSycK
EGb7t4rSc8dey8gwc50oYWpW8AL80tWI5Y0e5HtZT7FyWOOEgekwvVPFk04k3w4t
7J6QyQizyqcUbh7zLpaccE244/n2VjoLEyZFqKNDn9o9UvBuji9GcnYlzi2ZH60g
SP/0luBS5SMN1goYnGCxvBKOix+uHJ5WkXqTsgRmHbVgHff0hdWt3VklPrt+vHdo
uaJmykWpPUL4ZWR2rhwzQVF44PYoVoAKVkIABAvtk5Kn8f3s4AIs9qaCRY4FMhOK
YpzC6cjAe9z6oW0hK/9rWcixkSb1FEgqs3PL2K0KrIDcf9yTicRMTVFpgBjo/0GF
rTM0ourKuis1NZsWZGgkswKbfLnx22CYABvBcwT8/XdoWsqXBSrdDYfV+HjoqEc1
`protect END_PROTECTED
