`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0oCLTURNeD7eALCVennP7Cwl60nVVsdAPpzdkKgvpwN4OBlJw7UWk/V6wI4McTa
OGZevIQpX9EYYttiDeiY6/VgHq6TqlLATV/i9Ga6O6ocZwybqUFf5jElOZyQexo+
E1HJrNiI957T/PaqNGA9bYb0g31pYxSD87Wq005BCCD9Xy63QMYFphKPV/5+p3wX
HAKfbZgdM2hd2siMRFf738jS9AMqDJf3PjHyHQNAKIALpe5j0jCgX8u/qpscflZC
5lir79JCHLzmYSU4hZ0Gi3OCT6D+NkSIGW+/+9opLdMEZ+aw0jb7DSyesywVJdrJ
aho4ccT+LGI3vbCzoIAjYE9iVrBvP1sUfwgOGAlesFloLT+5sIwICiD9daI5+gHa
WO4Bs+PNpxY9DVK259+uwc2yOqAZaT04RzSZVVTNVWaAhWGO0snsnmnq8rvivoeL
FiRlzHZ1AnaFyDxJtd3ofQSVkt9oVdy0SOIVd0t0IyyI4GpebnW9i2MFPZ9IUVqa
1vpT55+3CGSTuEQC5OkUYcFJwJ3HkCjHyAU0NT+K9PXDhL1k3JO/gPcG/4xDJHBN
sc4mVsN0ZebUmiLuIPYxdQqy6LbqFdwEUpWhSeioR/ehwaDCqwurz0vZmxG5kc4k
dapwoZqau9Nm0tNgjh14q1izppuBTa73o4cFxSe0FTnm35eNFvs/QM/ENAFRHZdP
1pauIBbCp5w7Yi2AZScGdn0QQ0nvs6okjaFY1wNOkJZGncMyks32LDq8DrJJt0D7
FPjF6un505TwtUFiGC9kLNwzn3pjRbVAUzRBPQ9vOwi+/eODboASsA2MPNGUfpa8
DtSil3Mt/JXx3+Tab+ORGUtfvvIipuh7aV+wMtXiD7rlmyFc+dcw3LdktbtsHcs2
RJcQ3G825/4b1UYFp5kVrev8/G9OowrSKCOPCFAXNJHmNlMBwvHnpDycVSHnpyed
JZF6ef8oJI3hsEU8PYFigYpYZoX5Jf7btqY8lS6duFBxK4ODulE4JvLLLcSRSIQF
AN24yFWQjTFQj4i6SnX2GY9OEyy09/jmfINlDKvMueRfl+a/bEDeFnVaGXO/J8R+
7n9n42E/m/YHJ2APrnY52QDicVP0uUCXJN2Q0F52E/Oonj1aUnJYFNba37RWNz4f
OoYLVzVBCnqP9ZB27gslcOFVcRw6HJbaPuxktRbv7jQrRcRStmf45yDrsf+jeT7s
rGLCWPA2d/GRCGatP7ewAfdwt5dyCRvBoFZPXAoePMTyEQjSCTWDzzYXNDONL5t6
T/ptmTBz3Js2e/6OyNdBg05BGNn5/VbSxwLQyQi8b2PLA5ZZEN20EZJEW5RU2JFD
ODgXrsWXEuSaJJ1xvxhNc3SYiYlkL+cTwVUG5KyZW9NoSl2nkqFdnbOrK35LZoWc
O3d1oAMx6Lr/APhueqSWdBH/BpQnFwKaFZ5AQUuNX/psNOu1K7Dg4ZYHxL6Vor60
sG8MZnAIjWUGHAY7MTZFmFkScmmNhURpUWlai9nS3VECGRiJq4NRTupEJnLFa6Ts
n8OawFI0HPshuv5vQBUG78tNQJwTWtsp2p8gIwX2pYOxrVOEOpkDToTq4Z46XbeX
eF/0A1YNCut97sy0LDbi+R5gVmqv4K5QQkwmdfJ+MVe8fo5PuWKs1OfuCgYp74s2
277l13URU/3DuXHN6/bCx8d6UzhkN1RnUst64pqbwsps1WQX11mAw0w36DRMr7Gz
ADg3UHn41jLS0ziaylSDnGYKh8Rt5Ebytuf/gdE17DVarlr+couyJSxmpiS0cOt7
xNZJKgRJoKTahs1iORVVHVAnXj5RX9fnPMDweSME9rLsjt2JBR6q9/5BoOuw5n4W
bCL4yVMfCGClZOMn3Py9En+IRuqqF6Nds+ZMzL0NCvNhbKKnV4dC+hUqv2z1zpgd
4J0UCiXgqxBC+HBSCkzoE2ckIn+Igqu7Gyc26WqBEadQ/S/jcU5hBU1BKgZBqGUM
65dHlxp7Z0FczQyVhUMk7p6h4vxj/oIInFtkPUA3FzSjiivMcWnQvVfIAnLbMOex
QFbxqpeHOz1Vs5sjLb8GlQMOuZeAYLtRLZWPyM8dPAuzuBD+AVRKuHHujO18vmm3
58WRfgr4ReS6gV9DcU5GEbgx3E/nIFG7FKmVLomf5onvuK1jkbZJOXkyEmkk6H75
oFq3ZZ/ymC9clcqmfCduEnMJtMWtiOEHIlueXyJGDTcWpUZHMqQj+UYq/1TtbKLB
r1FyddaBa1ridiwpZ83BN+JwEYKzufYE7pLF0y4ZybNto2Pazt35Z3BpQHyjeuey
yBP79sFCpYD7+0GsOucmSct6N/cSq68XklFAM7E4ApfsYYcn5fdMafmPKYBrzdwd
CQFraBwmfDUv/Kkna33/YeLW0nH8B8EJcYnMdNf1+dbxjX77ucmKvTMbyWjjPtG1
OOZzMw5y5wovoFJyw4WZbTqHm8KXkW9mdgOJ2Z8m2A5BVF2qrGuh0KXGtYHnCmVd
ZiBJEMa4kM39En1Ho71Od2NHfTV6S8j9IEUr9IT0QNc8avpc25KTgrgktFilYptx
lTCWkPfrMe4FNeEHBtkPxDKfefnTMU/ejqyHzUmfUNq6LNtZzW95btQ4Psyehbgi
B5OpotpcAdio7TACmDrAN4+l3hi82Po2p+eo9C7Yl5gyIJXWtgwxT96ZQujkK8RP
vCEKAoWTzcWx2KYf9k4+Rp9icNHGbVNDXpABqXvNm2pfgSBbK8upUhfeLDICQXZ1
cqGbTOJmbLpx+R1Xu1M00GKjX4db8H3ZvP6s38ymkC1yt65jyMgdGwXnETnANXZ1
FpNwaVOqXRv5Nk7ZSLFa9csfsVRAPWwA7dSghDYqGZGzi0jP+3DIKGhBT824FkJC
SvuvzYHPFn3fJlhoN53cwZATq+vY7fWXs9H+dUp3xGyOIPGkbIB5ASnjdwWDzl4E
AfzI3otIjP9HLv9HFuFJUjhIjv8RtlkMBteDW6T4c8o7RPAjsltSiJul6wAIOfGS
V0+WrWc6FHbEuRjgKCT3IQKqsjgb+8y/By2rTciz2QtXocATYXydxk+WCQ8WgoqX
iYv50L3M0X7r8BO3WSHxgn0Xd5SLUesIQoHJGPv9ynTSIu8YOQiT0AVk+LXFsAs3
W6fWwzmCrXlxO7uqfQTgbP5vZyS7FGOqxVh7ctcCJSOUlwMnchQR3O8VnRYsl5mN
/1Wf02f5PUMijn6Ywy5zlbrCCZUOA8eoyLT9fdDf55XNysQ6CDm8MNM/gDkmOn9Z
JVFkLnM4ZjIEGF3mBTPSYYDfAZpE3yQ8Ai5A5kbKNdp1TTQNkAAmUP0vWemd1/yD
v/jAvQ/ojFYv2ml3TuzjzpASj9qsVg4X95E29dyHPviipLYcgLf1Y24/yUjq0Hh4
kizYuP8nkotiR7n34TZdAsznptvpDS+mMZb55a5g2LRouO5XNQ3bkbqeSsRFrS3a
Ke900DkJz5w6giJpVKlzdRafkyh4Mw+IQjrZYsi2sXnzAoi4YKXN5LUJMgEa+SHe
fNvWtGEmoGgMmIJDoniF5lXW1V3eOemHfFTB5mQ0Mw3RvrqGN2En+QF8mxHvCRZf
lFxBV6XXgKcPDGClMrgNO9YuO9BWvX2gO4ObVvZ/BOKh50E57cizF/znsiEgQBbh
IOOMpy5yWJxl+xh07Wk5w9yDwXy+KmqeIoTUSn+HAbxYlHCRUQvoJmYIrp7+AKc2
0ljCXldKrTPcW1P/NbLRjNKFhOR4Ut3e2tywFLPW9V0OaE2PicP/lSlWBf0R9g5P
BsIXUcslZ44ZAdhg7vz4YZwCBT0DaYQGf1jtVH7SzODMgo0nlE4UOTtkN0Rfs53w
6cFjLnlMb7kI9Yyl8YQQ8PYUmYkwM04mJBbJpdN48UL4xZhXTQSR01F4yvJqlPh4
E64uNi8IqpnrApqD2gouuoAFHkAPJiQA8o5HhWLVjzb/SSwLlIOICkCeuWZJH3Yr
CkoPC/IjCDMAzyWcc69RcCFO3tQPT/ydOghZrJOd1vsdcYbQuSEjTQq1oz1naiVA
bqrLHb3DQz2KjX2Xz4fkq4iAifShElceO+Sk3ickcjkVEXco86jQ9O9NP3T8JZu8
105KA23kWxUQezz+vRCQ/Ch0pOBQIirv/fBDF/lW6Uf+UJLUfH1oHg84GMDFxVn9
yBJii0gHBLOvXM/au8cqG0N6sa0jpAI0DpfCBBRYjsismE5X+SRqbsCRU4EEFI3k
UQV8hiJGr8PMq+cItRRt5gX8ssMTCnRwHp0VXDCC8E0rFmOtEU+/dJoD1YsYpCDy
U4z6iumCNWScVm6URRbEjT/tSNICXvFDsl7KfKCL2EYrRlln32HFfIiU4pAvYocC
KYzK8B62EVBPtwW6h9w3RWEijZVe/8oEkQuNSzPNuKcPDVLgO1KmoRYgcl//Ceoz
oK7mVR7V+KBFt5ZI45yVwbYOWn6IYxChL8KtUsBnFkn6GmyF/iHZPWG6vrmf2tmv
7/ECL5Ajf6rAQLrwS6NPOjC0FI3lJHiOCAt4NZ9IFTh3ux69fs+lrzMC/GqYyUIf
oCtiDdlIWzJBDkgwkHNu/bNpTIoMRoBahNCyZ/GnsPcAizQ+pES6tRUIVxYap+Sp
699jVgbOa4r0u33+3n/pT2WdlT+1wbw2k0mVeRq/jONWiGrtF9Fh0gIQjeErshI6
+JDaZP3XP93XkavuhyJEXl2HEAV+M8R9asAMy/pxf4YjphM7dvJxPke419ybey00
hQLAT3Q0J5p2Usg6KfDgUuLAg7M2XGy4YiSVDUlrwYjslT37z7NHZlFs9bpPwHmA
Qf9qaQnoj40bTx0f3eYjDeCEbo5zNqTYjpXkghdTwu4F9qdoyk2tAtehVCqFeda7
dyn8WZvMLLH7WfWVEFvjLTRI5Nu+tq5XRvW2hBSL4Oj/rTff90ENblfqUKlXH5iE
LCB1yd5ksFptLUOPbVPKTmpGir927CQHkJybHwjGI7ys11Ciwb2mABPdS4gy84Q/
OO2xw5n1RakkW7E2NtpfEFL0m6PlvmkiO/IQ6N4l7vOU82RDb9H7x396Wxpczbpx
PVmPwGgqOg+6waPkzu64sC55UEI7NL3NEYLlde0lLJubZQplPYN5JzXQKBhHZTXX
OqQwT74IzEjhqVu4plppTt3Q5yG5IoX43gMdlGqtr+9IKRJDX+DcB/yScCx4a0UL
EquHEM7YmJv4ed/2UuP6DS4zFIptJ6EkKbS0sq/E2rWL43WzydAhk9ighJhOrZPq
114ci/pi3lUB1upbiI0wTr/Qk6MQxhFmWOozfFiyoHLpxxpnFLtAnFQFSpkc7lOz
oTCH+iDefkwDRLkzhl/+prpNwX73uxD1UdpokQeeVYehHGmFlAwFqT8mYqYg9ktW
IwYqEwVLGYSps7acFlTdoLR1MDGMLwQykCA1C1fyAyfLhEKlKEPU3GSZKZ8ZKnZb
xXl25scIjdA74oZoFz6LEitGrj09vQvKgqQgG6gMvPThdT+z6zduW5Jd4vAn2C5U
VT+Dok71v6DtxgM5mdXP0fKB8AsGKze+tw3wjwy1Wsrc6zR9YUdhrNyJuXb6l5DJ
dun1nQv6Wc8FU8q6ndC3U/7w+/TLDvZ08/oQnaLa595Rk4Jbgpp8bdzWIW8w96vr
a72m96T0cU21ON+pFjN+6BiOTfSD+mloh7ebKl38q/V58joPIZQpVoadCsEjGQJO
R/4g1zmd7ivSDgB8q5mJjph8YJyRQ0zZj2Df6IExSo4kHYf7wHx133m+RAnDpKWU
yW8MmMywEt+A11tSTMc36QAyBpsLMe6N5xBAJQ0vkGKa9yP4YZ+fqn+jJEPSDhjD
pOCFupThM6x2NgNNanTsm7ZucbGPVCXddcZKjsfmC7KrSaD4i2rL8c5yxB2SAc0x
WFs/rMdq3HwjLjKYkt59C2pms+ouXM1JmjxB5s1HBSt93/+b7lH/75f/4d5Octn6
b+xREqSdT7sTPK+zyXj9PEXTrGdwhNvFrp5541Caw83FH5+okHDw2t/pfb6/i7/d
+qSBf3vK5Q6r+ee9OOcuqskL4k8BadgFkydUKSuE/gZs3idzvaJLH15fPr+LWU2z
jado5cHDki2i0NO3jJSB5jH76CWIGsUIAYGZhTVe7Z/52C46coPsmPO3SPaJmWsw
f5mIwPeuETV/b5UuRXvcMQRaP/V+vlfdKv5LLAmRiggVde30aPBKDjesGOfZiHrC
Yo9sbnEDb+9zXTg4dCZ+Z1hiCrCieLv20wX/+PRVNgrqjOqWw3bQF7mbOeYhaIHN
nylnGnQjw9L8m6ZTv7ar0rrCPMEHSiFwbmeu8xzOqpPbYNUpcqEYc/pBdYoIqUU3
EgoLKruF9HSyHNCKFvoldpzrdr6/QnPYAtfqO5L6PveFyG+obxCK/4+aMaQwtuUu
dj1TDm5Ha2EgkGTvr3Y7ACyf0jtcu9nd9+2KF8+o9huaQjJUF85SrTtG0IfU3xsI
AFtjjArx7YGA0FRtejFx6y9PLuch3JsmI6am8yiyRaTrLXBYv4m4ncAFOn/YLn+D
4ZK0/r1UU1nEIMj4IgFTEPUctuzGFKR2r1WDfDj93huRfnL5v+ucgFgadt4ei40O
jw/FN7TukQ1lO2W+pFuPUDkomCAULSRdX13W60axE6iJZONuefAIjxvmpholXOTr
XYEt2406FURT8TFDTSw/kNyQMM0AnHO4ysoN0peX/m/0EWg97ksKVYFICKDsQeDL
5s8hUXGllTBzRwmHtiAU5bTXz4eCvsx3rgjoVdwYOoBv+6RBUdkQvdfI33L3Q+Bv
WtKDaNzLQpLlPtBg/CGubYXNyINteSzTPfRG5nfJXpfkqmktGZbWpgiyS9TPCqpf
ivEYaFbJVB5mX8/Rr7R8Cq1nhgRKNPg7c8Nfm6NCbBuVGi97V79AZMYP4dS6a84n
Zdb3QPhUucJ1oa4cudb/VI+n6svtX9j2XD3FCksmCLpK7xae57aSU/wLUq+4F+Go
MRaoSfFpAITAeyc8oMJgxKSAybfvsj3DZdleAQofOwwLvpD3RZdeoA2VG7nN/ZS9
oUbxGUNviRjHohdF9UNU1VTiVMWFWsYtwyHH5EWeX1XV8cHvuWY9HfcP2KX1ri2o
XWUNqYJRokqAdmNXbfWjdR9doJB4Dk7Z/fYrkUPJJlWEFq7awdvUtopvFkbeiAXn
iKyhI7PwJuIxbvw+HeXkOF9jk7gobHZuiy+yKouXSdT7eHiDtQKlVtLuyNjw405H
qwYpJk2pFxR9R0dlAZ+wHd0T+DhLfSugCxb2VqUePx/lbgp0KQa208F05AEpBcDG
hoDXxOG/FAfa/9LLsKsuD0q1OsmOQeYrGCsMyhgsKRLUngrgtjBK9qylaSkRhQXI
FPizQxY7Vm4lgZ/ZwVW4gnKALq/tTIreNCeiQp49hdr3q3CxWARBj+hvCx0wW0aO
vlqMWOyznpvDayHFdnCN5oxkY6eM+bSdXewL7XaqrdbT4kIYnryHnMFWsTmFSJJ6
HPecFWFZ7yxlNpSCf5BGcrbFxXfIT52BouAu/w8my3G2+qXB+Vyi+/z2wyWuE1lX
Khm9rlLX+NQod3LRYGOx6EMQ0TMpVvRUCYSNb3XFxLtwhZCqixiw8ldMS41JXDK1
6o2ASffT1yF8bhbDrAHbrRl17gFtvvChV/X0hbAyHI4awNGuE80PDe8OB+9VSgQQ
JTJF3+BmtXrYoldqwVs/HSPs7+yydQHSFk6wqGg8NJdnMxwp/WDiExeS+3njuPp6
Nv8FDRWw8OftnNV+bqryz3Y/EC69e1FtMzH5OWlkidUK/YaU8AjkD6srVpWwo+rg
of8Xwud6wa5PzAEwepQzullb2qVMHFMJ+XF8vHo2cvYBQtQAz59N9ilKfSyPjLtW
EDT95XU8c3BzrdmjM5V1AhU7WjFbhuI3xaU0Y056XuXysxPCOqfOFfy1eUCjR/Ye
zFDf4oCgHH+w5XD1nzsz6ynsRyAaaAmYP95XwIplb4HsO0xfqvWcOv4ptTQp6lbo
x6JmZYXI9BVFRFyca8+WzQQ24acCwLP29fu9rCCGKenU/DMqYEnq0kjNZTOuaR3x
6sX7ddxUzVMz4tc8y07KgfPYGho3/FJPobDhXOGIJo9iSxWnhuhMRAsVsge2FlAX
8n1qPmW+cKiKlS1pl5Px9/XwIFVMfpWZVswAAAvZCX/Wx3+xL5Ds+p+v4QrWdFEX
OY+RacYSQzRtArHbMLu/+CiJkQ2O7sOYuOcOr/RPFem4o6ERDKUT6QFnGLfyl0o5
ZOgjI9J5E3fTyFgiWJYVPscDqJGoX46u8EyR0UtO0xpA9SMTGgVNJlYakbv2hwvS
vScdh6ilHEMUE764FU1DTtvymhxGFUXRqB8BL08t1M2XuXerdpLAHjbdAjOh1Yw/
dxN7YwJZ6ypPYBPkz7fBX9hOCOwGOIXAWDjCFOhpB7TxdwPIW6usc0pGWPN0OMly
/XTUPnrm+9PtGPUluohtMOtKs3Nrl0Ef9qHJqRSe1LRuq69ehKD5FnLsklJx6xho
Dq8LmXAZ5RMqPtD+gNyVqRlmZMzFdldDXOs9uofWeXpVNUi4iNQCzaONWwlDfuZN
JgB0iGKOPsJdY0dQlGtLoWj1Qsp1go+58kzlfIRlkbYN5EI4yAhBCdrzMg1WZNH7
qWcQ6bk+hPNaRbhhi5aEgl5D5SXvAk39M/XACs0XL/JpY48S8q4XEZao6uHdANe6
22NDFjBO6KmlJnPHHd67LTVAQbDWhP/Fl3YLrOfTLJ2B2Zez4cUehHzrgzFtxQgn
+oRYs0gppp5bi8EQD2Uv9ELs2s5ramlZlIpOmXOlzwcH/nCB2AttB2Z92bv/fm0a
WyzcAHWYmV0jbVpwvMA9KnOKUMjcDeOLd9iQg24nokdze+AtsKn/0ftwXBPZDfYG
4qzW4iWoy7kSchBXWztUbHFtfY5vj2EK0SAOTGXdthb+rCH5aN3jcTHeI0WqzZgP
zL1luC4dD862b8GJkxoPy5xjBdJp20FopMXxX1nHZ2TmAcK25xy4FOgHI286fsaz
h26v4MWBv9UfHiIiN/6L3/O0ylmMSoSJzAIChcvFZAE5r/OKLQn1jsHnfzGkMPR8
S7DyxThaZDzhvbnqqfLRp12RqnVz3chkiGedDsYmKCX2nnY5xzcCmgBBim526J0r
Q+AOc2RI2ZfbQwizWaWYpb27BsP/VXFMSEjqpD80yvve6ObtKBYg4ygMut1jDvZr
8CDgCUOPK7oTXPP3fuql7ppSz6bgguvbAHYbCtziR+mJ9aMBmqAAm0+abBWtfu7R
FwqHk5S/9RFu1oPBhql4NZOmhxyOf5MMduoSdldf8tCNTcyqLpBH5vS5EnEIoKbt
ctc/BtqDNKlTWLGwrXF3nYT0yuhfRoT/WkpckwaMdS1Bj7jUzYBILejCJOwN5Grt
+495d+F7M8DKuSDWlBLzaWcLhYJxmztsNI2wQOkLXNA1MxCooKoylUQvOSns5pg9
587BSdLxJxJS/RkDw74yawFkIkPnOmQNAGr7ChnijmmoeJc5udbEUsHYdqrapf8K
4lJa/qOtulUA3jy7dlZma8GoJweS9HXjGcshRfiiGQLZ07iGyVqjFY0SBVai5a3m
BxdzFEZX9FUybbM8xZxkBlrQVcMOt7fUMJvkEs2+2xQL+MyEvj5SsAyjEFHXYL+A
jB02Sokj5LTet3FjfhAKFStOP+ZlxvJjbOcS7kr0bg3edI6wa88EHtOVMU97YwSW
ci5WKAs9iBQY+c6XNlbyuSvIoOlG7fUdmQYgfIweYCWmyakNZzoqO0/SB12/D7de
60m3gKeEMuojLuHOr59IjVkHklf+ahNYWadSzRPqjXKN5NgeTOKsWSHNFe+njyQS
fmbD0GcjMOxnC0P4etyDW5OIo9ngDGPgxtgn8w9wjY3scIsR1RWRCl/NoGir+kEt
sVxevYvIqAKoIA37QmMgmXCyrqzAFS+N13DGUkaj9zNkj9AJOTZ/tI6OgCO+UOfG
Ltv3fFKYLttXPghwBw7iOBLm8mDAUXAs0o0zJojeFN6iEpyOUFBhSIdpY1wkkvXs
6kamA99p98rmoE5VT05rzTitFggyNIoPEpCM0o/5dQjxsX/w7L2EQ21xQr3aIeyp
URj41Zu0J3TT026Pe0jMoSHDBwBecGqIm2FMt+760bW+k1IGZ3J1eOpqF57pWsQC
oPWepqjGiY6mgTJhH5s0WOdlYiuDyO6FFFwiLebz+pnAY+N+3/QhFVoi6lLGHAvb
7sij+JMBQxIBX5/2GUuQbBEm0n2GMhJY9RjoE/0wCwZWUShQvyXqQlO0ekmZVV6a
h8XATwb1ITQ+lhzmRERVtYbu25psKZD98u93zb2Ing9vTQWdPHNbQpRLb1UkjCwz
G7xpNjF9lYJvtpzQJId6WKPEPdHrh8PObZiTs3dhYuxBwFBRFtgG01zPq/CG5n8s
/Q//IutSwPMigCUDFMIYHdyhaTtmk9vSzMXWv6f0aHgf17ktzDSA/9HKF8V703NS
0NLDONGLpruLSoGwwgtzintxamJHw4SV+RTS6hS/acBmbjjWhqG9fo2bMUww+7X7
it+t4tBBrz9TR417fLAxcd0D8zE35PhT9T6PHCWL0brYkksWtcr4MO4B4bQN6ZZJ
QaXK9ZITdKrxNQF/yNRgKsOkHGRSGQZkP/pgRyTs022EAtdMOwq5ems+psLRYvOc
Tnaph2Hbrd6FjPF2wZttQYCQoXrDm+1ExLBT6T4yXz5OOLoTztisj+teCzRGvWax
SMk4xhTJiSems71OM8vemKR3AQYs+SRiv3wloOV8bfIpugjWHfpbT73khoeKvBPn
rLHf9Ka02YiB+Zi/Qp9GRoWaZ6Yfcrg8dtM0sOE2zjG+O+g8XsxqC8H+GRhT39TX
HGl+7MmLrIqzka4ewvxfVaA349weq4Q4j/KjQoFeKB+36l1DoCMlJ4gDMCg9sNXB
4VXueBd2/Wlhmhmks9Ib76xcEHLeBJvTFMS99hAzKfI9iORGf8D/PoEMgMB+LUAG
D8rvC6/GUV4EPwN4G4AXZoiqngK9JBWT+L4hYUmtxSe0TtUYDU4dlrT1WOukhuUI
jMUOcRugHg4As6QX441f8/aJNSpeZxWlFkTYp2tuRW8wrrvZgXGpTSRlOcGbNXLV
n0ZxCl1HeTNXl53u8xl0p+JOUei7wmD1sEvieyXB047C+IByJmKdbvG+Ga4fRaz6
LjYaOitme2JUtOdJ9B1rlR27c20+8dyoZIFKUzrXkhZikclebPocpt/UIQIYLcXe
vajLWaJMi+PEhGm7xg+Iw4QvvdX7z5d/nA3RYQuazfNaFGQAJPVuXB/V/LwR9X/p
A1+GlTP5Nhstp5lhDuANKrPNESwIyyENFP8QUW6US4d5fVjSz/Kb3ry07wxvTGaq
BGC1Pvr5xCbfYFi2rBqHHKp6oUUqI1Q9s06OBkuDHVAiyXLLtQOwrB9u181Rlrkp
xDgYHMAzdPTdJVKt71Q5MogIaTb+zRLMjN4y6MHpb4COgqdTuGFzPv8GKXMiBdil
l86fGrKTnvTrfaGQsGwuXUZFK7RysKUsR9F5UfCMalbIzfeO3RxQgeCDwmRe0L4I
GUxyEDJeVv9cyt8tpprFa4jbYRo+DNrvNPWys00wE62tStW8/AZG0hvepRpJCWQy
4fTClUsx4+9tGjLUD4KjJvNquGyim0WTahIAelGyorvv7R4L2+B8xw0jxrcPhg4p
T1WlOCyGLQKC1WyQP/2Jnc69SL+CiEXsSXnHK6crfhyJm9dY8LCnJAeFEdRqrGWy
INR7ev6pT05gfZeKs4FEKeeT6sYlLfPzsYPJzeTN6cZSpFtwgggHbJJ63+kXzhiZ
7FU06VA7eqxXOMyyGgLWM03ig/BILCpuqGGRiQsfn+nf25gh1s5Wpyn/vULucD8K
iSTB3+bSohotS4aVEBE+5DYjnFNUp0rG0YpJw+hkO1wnGDRUMluCHmX/C2ZYeMh8
r9UlVnEjwdrxy74vF07AmrReASIFlteMJnOMqX47iwxukp0eD7YMDtpMiqzcOKmZ
9q3R3vyPBEcVSpTOLOV8xd0N45XEUnGGkBRjSUvnSa62vhrtvfkKL54/i+cA0ImC
QpjA8Q6x+kUeX2BbPj2Vk36tLpymhMy0sAbF3Xzem5oRO2VjvqAZ/8TkIKFaxJ99
7EvLXjrWeeGhZN5sJQPTPnBLfQ+h3Vw/6rkgbcbbokI6Z9hyQQbzVQXvi/IpJTjD
sPSAZdYWuPINAOwMiqZ8vFHeyVO6IAkSrwJHgCkRXxWStudjFctS/DSPxw5HKliH
oKp2yLuskYZK12Zg8khM7+06JKvZz+rKssWjc9WiAPBRtXUEZW3h/Rb5OyuLGyAd
WZo8/WrrOEFC2HPy4YXme4wkItZYFb3ee5upj35Rd9L4wMPKugl97FxH5l7Eg/vk
KosybVRKcCLurxK1F/aeWaIlgeslcCnBuWkIGlW+oGOUSj3BFt7QQh5oBWHEUKs7
/RSdRKKDfgGjcFuYEAE/No9my2MJPeMrkLWACvCFTXwmsNykphPCBZTEjP1eoaSB
l8ZTZ1aS6NdJZXnA6iVLZzxgPfINoIXQasAExHTEiMs3kutuyICYU0VZUtx4PYTz
cUEbXDQ4vsDQTdoZNIYYzbt/kE60Vkxr4KZcTin5SfC/OEsnNnUr8IjgQnHxBwTc
8AiKjDLpL0Fm7NUn3dI9zrrIa1agltc6dNt9u23L6dtcxd3gYCy000vGk0PGeG9s
L62mQTNejNTeAeQSyUd25ba7BVKMPPaNpXD0bR+oWMHP0HA0OOGn0pErd2yZY0zG
EhrED598wTYYe1JUsWZypyEEpOHsuMK9mOtK1J9jr4wsiWIh8mWlniGNPjMUNhZc
AZCsH2xMfNJyYMbGc2Gr10Ch1krKGcWkgMpxquXd9OLkRmN8eMqb+RRg2hJSzCYN
x3uu2LDh/4o8isst8TrckcAp1jGTs7BMUKj0VmBVMJXp4e8mpKsWQ/eRfbgPSIqp
kZ9lI3sMSYOPL1cd2diAQvtaCjBARwry0jHj8gAPpZQ88LQ0n0yX1ekEXEUiA4V7
nGpxmvw08s/RCEOvLcvwc+gylYXu31WLIAoLz8ovJu0CTqoZcyHPllSbjlHq6O8t
IuOV2lcIVX4Udlew77A3aTComPiMzVt1jTznAaHj4G4Lf6kUGy3QifVs5OUW2eX1
jlPd/NTtSVTRHNTfQygN0oanoifCTgcOgQI+ILcuZS0m2icFivpjsxtXh2FwOaDI
qgyjTjfyHc9T9IipVB/3Y7sVZbU6aty+DLQ7sQeDTQj7kyAXNFv4ArhNM11x3mcd
OtSzn5yRDSPS0K49AkgUGyvzcTXjAFc/Vy49TNThQ8ejO0ZAaupP8IvJaST8myFb
7dSw/l81MfECmQgle3jptQurpvRWIxbKmVICx16sJmGT2qfzJxpkIZ7E4HSTVcQq
DHEvf6bFI6XikHGNGgs/k7CImRAZyLTXCQMn6bjy4BeB+TgzoPGhtoYARkUfEti3
w16gdgYycfHykvDmv7BAaTvWgLxz9lvTyJADQEYpP/UZSItGJRttN9lObVUhP4Zl
d/UBMgv191OoL0JgVIDx6tWeD1Hq6rU/QzZEkngd+T+dcULuNr6swrxjXjmfhanD
ijqN/D8qgg3+t73LvyZJwLKynhcq6qJO9ELhpNz+2wJTWL0M0kopeYQRBcAQrmWR
5sj7m5WA4vdJ04kVoTF5C7avCrzAsBYqSnyzEae4LymD+rCwjLQhppHQISKYqt7s
lgK4ZoIciebgv77VPUpKRKgiJelqZN74CrNRpZTSmulZ/nJfhwzQXdZY4pvNWFj4
pGgRbpRJihNru7b7PX0hEgCGXG/HM9GTzHGXibWZea1+I/oOKvAMfOXMDp8rKuKQ
dtRsmAn4WiKtSW1nFJRIiWhPsi5oti3Mx2xOJCMqY/O8ugzPPt7TYab1SzZSE8IX
qKr2rC2LV5Hq/EY3Mj9nZ5sFssU0wNIMqXW0ecEDR5LXg4A8PjphPYohwuCmiwYv
wgRJXV7Ts5dMQQjwz52V3fVIEyBv3PF0/61feMj0v6QQu+5F8B14KEYeDCOxHzW6
/jjQ6d00e7xtuXUSVe9/npnE8+IoD1rXZmc2kvWj9aoNk19t1RBKSMhxoxKKuwTm
0x6zKay9MRHkPwm6rk1ppMI98ntGC9nSJ8Eu2M4Vw5zs4SepEIqoQ9hAXdB6GGiA
4SYFK59PFiDTfK6vTXD36BBgvgtG5BcPbnxmJbzg4BcNOJeH9SF7Xgg68iy80h/S
dFBkXx1CK0bQSfZyUDf42Y51oPBgP760Wtj7j73n2muqjcZ6xoxGyUDxh1iuRIj6
o7sADAqh7hBrf/6Ln1bSRA9iYKVS+PLU0iaL/n8ARQBV/KS27xannPDr/EFuUwxq
17tJbuNQkY5+TPsGCEqS1aqwna79uBHsVpSUn0tSPzuT+GCowKUyrbrVj2aUZiFi
Psu/dOGK77JCijLutkZOudU/YYSPJsqfdu5Lupies1tI6YZDrGHXv5JzAmGwaGws
XVZw9HvbZq6GRZLgM4AHtw1HI//Pvp7MJg337pLss4G5uwwjl7lx4KbyUbSIiRG6
Kf6Y1LLvRCCHMXa9PuTv73j0xaJ6uuFpoVzEwFQxsQsEp7pCf0VtOc0MLvA2O4K8
QVowL4Bft7dcOhONRmsk4MJIkame5e6WlpqNeX6HFQJpYGmXu7gwSIBE+9CVHW6Z
ss8UIkkw7mLc35NOhwHUbIw7vGzVloBzVHr5A2gTlQMFuSsZtlOULmnrUmlelwfE
Bam9qcLsNYOo8Bag7xXasfM0DraOoXzs7/8T+TG/xNwl0jKctJdmuWEhz+iXy5ut
+mUfZqrxh/aFta/C4Z2Hie5a21DRbIVVsu3XDJanCqwIUYc7XYOOBTfbEG+KyLW5
PSSyXbjlhQr7MIU8NbLMoNU0y3J/Ww1NLPZslWegjDUEhewzuftDFl4AnaYfvkFf
wZnVepfWYZZfMBBlK8V8x6fIOKeMRiGsoeZFXiYn9RTWeJVzG3wL8VPnleIBVacJ
IFBWLanP6jknRn17mIb44TpCG48EK1mgueZCSBoY0iOW1alFqLis/9EstednhO6v
fkDOKsbNB0PslRTlbn5lm1TIiUZHUkLiPWnZBZSA9eiHpF1lJ9qbYhpIv+2cutuy
5dhzB9dd2/pF1Ls9LWeGwUsKH7uWBc5j0vLRXDiwRGy5ZKImDS+AHXVrpVUnCtLY
Sdv8we0ltsji4l+ICVNpb+O0rBgUp1YYpenjceFu2KUfC7U3zE97SWorijpRS9kO
ShCWYFuLkP2+t9ijQHAcNwUA58uScS54l4x7Ul2LuHhzLpTVonP3AEHuR7OMWzXA
Tr+AvFi4AoH+nsuc96qlULjfJzgFLGUygz6PhVdH1PtTVLU9vJlL/rzlZgT/vjbN
HRTZS1BjzOUDDK0egFlX+2hMyA6gBriV+WA489E7s342edq920mZSVy2Afi4TwWm
luCYHGuJ/TbhnmUMxzsPaCWYQkZA9pLBU+uOLlPp/714JxIIyke6ncOhN8ZsPMW3
hue372k26k3i4S0QKgwAIW+0w/fLCJDkC85PWAW6SA8bnPMzqxMNrEH0kptQ1fqR
sNTwNfF101M8Nl/9xCyLjK5OJqk/zkKWYyFmpI62pnxcMZmsbctCmLyBcRgZDR1Z
kftaS+8ve3CxdU/BsN8cpL1A2UpM4AO4vmoNDtYxeOLAgs51luKnFk+hpxj8XvTx
/XUlvNXfJETmrejIYny3fgS6dImR1WtSz45u90pZQE7kvxSY6U0aWmclDF0nSVAG
xJBPoADotBfl5jC1MFKrCmHIMY4QwWh3nvhZx0pLJFZxN28YJuxjvmaFazN66tfe
H23W8V3eaVvszaw8AH55NtcUuXtDzMxHQU3ke81Fr9aSo23mozzPK46e69Ulc44i
JShBPIKx0CWeu/+0KGWHuQvpAUedMlY0WB1gWy0vq47RWK9qVcoALD/atmgvk+n1
XuuFyxXmTyIxJV+SlpuIsZ2mRJMDheqYjia3p0fTWGqgYMZ7kzA2gPcjRJNS5SqW
Gk261YVCPEDFjt44aOYNuhShDCeS9Q0tiF9mRuWnAygsXmz93BN0wBfWYE80LWph
Trsp0jS+6YDFMreuCbNZuuzdh4d8Z0uTrr/tEsuxJDArp/xaTkXLUTmx7P99gMnL
WrKJAjQs+5nxBFxqBknwyeNcGaabYdJCS/ekUT0MbbILYQQiHTLy5R3Io1TCwYGt
NQaRcCLHguyl1LdlNVid3xF0ZbprzxemTi/2+om6v87xhRs9lBbsCz457G7lLHNj
Olgp6H/DiE8qxEp7xshZlZ+FJTcQVPa8dNjlV3UL7GODMcrWJmPLnnfAYxWvrabb
1NZO9igbLkrrKPmfJQ7Qp9ftF9IyS1U8MeFI46+uTDCFdShMpl4NWrxswGmenPFc
JqsIpPaMd6KFZsbJba4lhSdM237mvzWJWe3K4SR23z3NkhrZP4yCd1YZ3VwE6GR4
D5YIzRB82X2+TDqopb7wXE6Mwq3MPvRsYxU3jWdJAEdzcfTZZWPcDaFymb+w0+Ae
COkMvbLHzJ/MgWiTn0KW6clzYOluPbkqiOVJMGMiszlzcQqiHga8yW0lYg1YOWiu
EtkwPMAVgeJQXCYxTE/6XyLzFAcbjPF5xbkwWRLjr5K22n/uM9k9Rd2ThlZ99QOz
1DFD2nCWlCFKQpC3g6mkK2XkPl921tPAso7fExH67lcB3bX8whq4fmdztjTo9Cu8
ABxcE7BjbrpoZrKJnkdxiqpv/SB1bEEs5Iiqj4Krlb7nPfNx0XoVqLcwpKlFsxE/
NZctExvozCUgNv3sZPyVDgT0xK09+5XmwOv3fRvYIm7rkL6oDznSFUrqGi1gub97
7XvJ8wsl/Eypw6m+mJZI+aP5+qp71rybmCXLhX+ZVaD6YzzPNIwsTJyLpdDbfYbN
ZGTaHCQV7poR46SqB1FPbnz2TzJqwlwqkJ2FWR2UERmnBThYzmeon5eDKA2gGNC/
ibhMC5T2llQXLaV1c1oL6iNviRxjvx4asiPm6aC8hJ7tMXH9Ybl2VBjMD873qrUq
KuRoCB0rNV3CdbWrK7qLaPy8kkHwlCFK0HeOlYQ9tjPLjj3MAhCQhfPC1yrxB4x+
+Hsr/YY7VgNW+N+c1IYVYteLsa0BOwjIQM4mKRbElgXAgw57KNf4nD/vkg87VeQy
3dNFQhDL/7LsYiKjx7jUY/Z850ssVH3ODMQgaa0y6C6XMzaDPsbO0lBT5meDp5L+
C0E5tk7ZvhpH4tlJqO1iNKNCAD7T0RKF3TOyPhYJWhlb5JW96dPcKv7Peq4saD49
62Hpmzwd7ls+UbfWXWEG+w30vRffHmFY19Aq8tchnlgP4juUMaie8UUll4wy5Y5X
+lzzaVxZTSWsZOuf3PgtrPn6oq7s3x44knUesP3lcQMmadXzruUB3lXhmQ3p1Xng
24dHXsve8W3kcwLkrTDC6bzX2/LDuvzcg8bbYACNzvj4qxDFZjSYZ9x6vwRubfmo
dd/tCxepwze/pzhKgsHVliC+Ob7RChT6s9LeTotDH+QzrDFRgACC0vwqUfnyi98J
g4ELHGe9NYr2CenTZVbQRSkmNyw/qgAOl//RVWOHzmv205In3kPqi0AlV16xIV1y
BZ+Y/ikdE6OjBzkZ6vrfOytZIvky7f/5cCU/aa7P7XxRm8BdP/aNxO2ktVLFMFJT
+CQnl8MUeAbf1py25iUFiTE+NCxbXaC+ZwTXNNudfMCHE894WO7Oxufd/E4rnStG
ZRpKujrEwnCvQkwdcL8Nn1Fi3p14gR5Q3Fe/g36Nz+xrrWKJU6+FivqZ928PhQJ5
lWASHt+jxTAdbqsUnTZnLD9NS5P77juK6PmCX7hao/NKdKS/edyCxPD4J6B2Vwlw
Z9eteGFWDkHrZOCiKlRFnwRqUI2RIGgCRtc3A1q3Lh1cePAgAsSWh9d4k9uPKbCh
Vt9+BgDEuPkPGiA9NYr4K8XOaskTeu/Ft4jOtpzzLwVdTrnTUohj2iT1oaE4/spL
aCWUVmqoTWpbbGkgsNmvkIzcefokTpY2jF9eifmaqYE7bLrxEtsEv1sKSrWPwYbb
HqYGKz8O2v7LCipJlU5jNtb2Y7hQ+cqASI+GxtlzKmp+4kxq+mFNywtRbllPX7dF
6gtbKt2KS1pdtg61f5fJw9Sbl+U81SriUcCN/oqqqna6VyEFsXvcJvYoXW0Eoph2
GC9BZGSwKf1/CciixG5NmWdz6xdV3ZXcw+BLKbRc/Rg3rn0f5CrL5dvhvwjfzVdz
UzgrXuFCF9Ae59NK5mOcBPAwQx8rUDManTdqMNXOOizZaA4G2PM8pWzXlCWDxVQA
3T+TJFPy+oOrDDIulFxTY2/y0dFqvEqeu7qRYx32mN12rA55XTz/ETJJ8tf5oyZa
r4xXrO6kuM2f9TLSNyWPkfE1mdsthEKHKnCuI0lnzsDtAZ9F0v6xhzA9M/Nl/EMg
WFwLI4uL338EuphP8LRiwJ3+Ss7ycWXc9eQYYmisoX6nX7euuUlWUJVBFtjhxweS
AckUMVJevDkDX5KdTuuRqkfh1JgxYRmlPgYaZfgYhEl1aE7MAEoA1HNSjF/NLFaZ
42R++ZIJgFffI3D63uV3eL0PR+yvQOEgbyVv5KTqawtqIe9JTJ1lZrJikUmuIwUA
TtvdODDaKD4hwGfAr7aEwl2EPLrAAAjti6Rkn4d+ujZKWOUP1XZ7dOCRXY9dc3v6
zuMnhbw4ET8cIqMT3crazWASi+2GQP+SzjJpfyYtvThf8GfezXFxICMbLJm0X1/D
WXY70U0KnZIeTpUnzSgLT+usL8CIScR6okQTXz0O9R75cDG2M3ckm5pFfF/txxOb
ekJAK03JAYk32LakDtz5yqyhbOnTjvEGTTU0TA7muts8k3hxlw28AukQuNcfK1Ap
aHWJOsV9o+J/moFB8/aZ8Mjt+nkTd7/xO87l3+g5DWGjSmq1TGyV/gwlOWh3vXxb
u8gcku2fosDSJqiwhLEzWSb+BOFJl28brPQ/kQfYWjFGW8DdbT9AKX2mHwRi4OhF
hMn7DUZu7EfAOPqMhPTLr8jXG7+s/FAI8J4cRIgxqQrZ47KiQY0hTDVWB5yVEQgg
prJbrwDsBHzSzeIfw3z0ZJKAaAEwEvCun5iwAeylZiZT8S4byJ+V05c+k/a6oQ1S
tOdTNMC2fIl2MHecrKsnBOzskRO5Sy8wmeqa3Bb9nho8cC1wGlgnM3bQMZjLTSsW
KU+ZvR7/S5Z9/yIcMq42EuFfN+7sT9sL9uY6Suz1yDIaHQeViJbJrbVd/vSlsozi
ZwwhHI71YfFpZn4PU5GT5xpgNxyoCmGTrl/RZZYQPvqIHPciElFt4wARVtrWMxj/
qNB6xAt6pFE6A2VUWBq0KZUjhmKnrQi1A104/cfRpYOO5Qr50I8vWaum69n2RNNC
+YXVz0zqcOMRHnm2t87efeDi8efUsVvPaskiqbQlSX+aO0XklYKHuMmZ6gMauVbA
eO2I4YqVU7wzIwqxucE83Jy/zY82TgaepaIDshoXUZJyjba3aJ4Au9+jWxhsaHWf
Bdc8AQaSgOx00Sn0vwWLOV9UdIQ7kwtsjDQ/98fPsCz8kNqaseyu+JZGhMyE91zb
EbCPlIQkn09T1fkblRyj6XLKyDwcmtRGHbqSu0ypYkVGYj2jO6D5iKE3NzrqQ3rP
s4Ag2QgOP/UU8H3vDmRIuEMzN2HTOAwZlCk/3whMwlPt9QOisrlMJVl89uRozHsN
ZrQQHFTnycPj76QDdcWPIY/MriqCk05TV0cZNy/xCOW+186O2AKgUKDPn9/ahoTE
4Vl3a/gJ/boQNpltsCBjsRFvhFJCvnudc2jG9g6EtPyaf4VAxKM7IUMzvrY1Pyrv
xoMpK4WrM8bx8HmVnourO0pIdjIXMhx84i2SpNwHYP2wqdCZy0a5WjIJDB5W768g
BAZa4xz/q2Vj4pz9V/pknZFwiwkhcff1ADSnArY/uA89fQbhn7DP4V6iukV1dLmf
oIYErnjGD2XMztO30pbjD4/sDGGUehZ2o1FzQyNI0WJ7AKMyr/D1K9c5KWoxevS6
S76HFzygZbj345J6uDVCR3VO+jcL/lwLek8Th7otPzjgavuHnHqfqGz5/Vf6/iSD
pfxYARjKnTdijmXLLGdE9vobBP1XPlnuvWkuxoHzyCd/yygoB6dZ3PaTs8Rxzsoz
qITeWBBcVRhalwhB3JpidIuFwRT29UfMiLNdD8EjYCzjQaPI51yYXvyFfPvE6LHN
EEMvOmalZVE1ZePtsWpUXTPxMQ3HBJyk5rj4ESD+M5nrZ29xC+VFeJUh2mTLHFFo
XNadLJvSqxrgGbqXz0H/EbGM+rpwEU5CjkYLNyanzGwaIfB9ArncqGR+ebaCZiDn
doBHeKTmkuV4xm9q/NOGGCWC/RMkfmUH6XOnSlZkE4eP2Q44H0pAPQzkfCFNCDqr
hOTjU/croQuxRaoD6JI53TxZLrxv09zBcARvk+BZL0kqkhFmHlt3+vtjuBrGJGOu
9qhIFSO+o5qTr7Uo/Nsa17S3CgwTWhMF2181Oy5ByC5v9smTCfb/tFpcfA5EWZG3
eFnMTWn92YTomuawgGpsr08Wv0KCIrEJYHwAg7rrAbtxEjRuxFJYaVjpzOqIwpsJ
jAxcXWTknTBDZ44Z16KqlZ1o88bKIyRWaj0z1Chn/Jgdsbw8ulNsuoeJwJpY/mnO
svy8a2IYnTlT7ldZU2/g7XHoBfrNOqfC3THYX1Ua3Tzhc7YCipT2Uxta20c/wT/y
AZ1YkvNxDFL4b0ixHL/yeCD4OYEUF2ONg5PwMntutdcbMljkpM+90hIw5vO1mHDU
2G/zsR0lJw/ySHi2etRBSzgtim0GAlusWBArSFSSwk5oi+phmDTnM0J66Zm09yFV
E2LvurAgLZFYnfT2nvH5yeSNkHgsDkesZ+au9HjbSKuCE3/dNg2ns4oilgFOF8da
jNuXWcI1dV1WZIf/BlMABszPkSSbFMN1jkT5zkpUbIYXn2E3TEO91aq6yvuL7KAS
/I+JHUI+GFCeN+QTmMPwny3GVQjXbR8tula7BvVmtJoQIrYPx+mO8fSWtWV0/tDa
fOk/H/BGlNiXwZ4nYIiS8llNXS/+eFk+zVyrATzXoL4yZ7RCcreXLrlhjzw66LOf
ztoW0Uvm/amcJNDLd09V3AE07tC+dhhYsS0e0oKsydJPAbG+YsfMkELjaWGs+tan
jtxqlxy68vZ/HZ0iyxOVhIy0sKRqOMkL5kkEkwX0vtHEptkZuPv/1p65Yt6ihibJ
0P/cwb57m/QfH71+O4uBvHpiwcu+Kj5bc8H+X+EvHyJp+vB+GN/i5V/QnOcBQROg
yypc3y0MyyP/DA+fVOPD8CAyDUcQrOq9/nDDt59H08aVzKyTVnsj+r3i23xO1zLX
bVs5NfUlue1ehUxTJKlMxZeVbsCq288TfjORikNacuRbMUYIqzlIPkXc+gw5mhlV
X0+spvddsOY1xCPHe0RlJTMVU7hWDccsMkcM6WYVJGonDEwnx9H+sGg13btEL50p
/6n4Lqj26vZwZmkZyITQ+/hk7oiM98y4ServnZdPoc68dxe1tULI47Or5ufLRy/3
4FObrB76HVx7stfYq44xmTVMmb6eUP00TMtqpcs4RLJ0bfwvQ+SzS1q9s6LW5fLM
Aia7sTT/UU4xxuKpY6DdZ+3Rz3mTvr/QPjY8HdSgVoaBTl6pJm7grlkQovtmQw5a
bCQ2Sb4SsNunGXmhxq8wHQ9gDbUx6M3g17NOy2khTpdb4WZu7VjyxU7RDni5br4y
/NVoNMrmBFe4E36W26lWsZVvdNYuGGe/JWdj4OlYeriVVkrmkLaNO7k8sg2knXwk
RFll9SnMQ7yw6JqmICkNOCrzsCvByNaqP0Nz9yZ8FTzyTDaKGVODRPK1fNRMFXND
0Fa2Od2+B26kKaFBE43Hr9AVrmvlO/RjzvW8liETDVIYlQHK8csz7q4B4apRImlu
0nqBSSxV4/7247IF31oUkKWI3nNGhazi+jGYFPgRbTSzhXnleumYAntiMDWH/H0a
k8sYDW2/s0OsfvtQJi5RjC+NemEwFAjlxGUVl6neq8a68klLwA7iIw5J0qBI/1ym
U39jJSP6M+Go7MGIZTjUA2i+EJQD1tO5TvDAcm6Zt0g3amE+7KqT7h6bwQMgmqoB
qTOV7Z7V63f7zfMZ9OW4MSGh/Plwx6KQfgirDW21R6mAOCX62Rv7EsWWniHzvGTB
flTKahF76iq9LLKSqT1n+eqIBUFKXPNTLm0wWZXohFB4z9Xm2+N9r4Lecxc2vH4J
Q/+ZRDSsPSkQHZmj9Ug0V16bE8JLK6xBWUw+bTOJ3tFNtcMAq0kb+cd3BwTfuqe3
bxgxGR6xJQzYGYKWiGWXDeuG0XIqaTK/U8ISTu+63s0CiFDK3jsVmMntdvtfjmiR
W2bygLtr3IOzdbgdmK4fWeOQaJOaUQOS4x1LEHs+nOE4pVZ0aX5R93HbTJifUUXR
+zAjeN77eQiYUsUuvHohcEmpXCjcGv5K3Kq76pfcVS0tbICgoI0eAOudQhJXZSsr
ysv6vwnYQMD/Alo2FwAWV1N53Og0JmXnJZ7UWRSaZHUmGd48KObw4MYE4bNQkao5
JN2Dy7p/TMk0c3rHCyH7GOjOCEvGcLxzeUEtREPoIrj5m8fqP78B2T/iy33pKx2s
zA3EQv5rmtq3GtAvAyySCE73Pn0az1fwm2zJI9N/gELLf3Nu6f+IMSPXkhYZ5lj5
droWwCYm/53Jjzvzt5H0qdIV+D2g5IdNQphFwdZwyvTWDxixhxmqwDcc7qRhIWPx
zU2JXZQEan6oRTisErBXcuybba0SpMBSsZMkPFaLMl3Tid08QJM6z9PhZq1M7rsR
UzpiypI/G7C+DpdkiZzZfWkxSqeMVoxjMUkTG2KBQuYbsCidvTvSeTvaRABoHyVE
2ik06dvNNHTmZq6bUCvFfVinyeCSRbTk/eKkXfSJjXdP3Sl2d/Uj8+N08rnOPp2c
O/6yKMKUKnEVRL4hdomzf2TnX2e5MAVo4wo7MNMSOYn2Yfg3UCm3rEHzjz0V0hvb
wyZ0+F1Rtkf40K7iXCviIUUzi4vjk2Ghnmc0EqRPXFoGNUt75ybuzWiur6YR/8/H
XKVHfqZldLcoFcDoIcsmTtuQpAybcf1wangrPCKSdGPJM1KKoBy7gU79k8ug/ydn
Bq868JhL8ckAa5pWCaCuuGZYFuyLI52kJ6bfjRaxbXqKQ/2ws2BTj3bAOdqedbbJ
07pJzjFE8kUoHxwPQFKxNAkZEM3IibGRtcv5tDA/P2KigL66yLnKyFLaTqACSNTk
vJPtBeyvXJDb1P+tkDsj7rs7Kyqk5NJNm1gTkOndURMlJ5kPNg4VxY3cgMHSBlgI
Q747U3+KleoDZki7SFFnncQatSAAnsRNZRNwdDUo1Ohp35EL1CsrchUeE7wdrQoL
Bp2IybwiUyUyX3BXKRKPcUF3w+rYVaHmezPIOaCvo4zfXjy8oFm00fVKnNwnUhpD
dOST/EfL3WQUhvzg50972/9OSK8MXShQbC2hDYM+a9OqWIX6nm+2XkMe3yd0u11u
ca9S8lw10odc7j9D8L1TD/Hl4Q22HVHVf3i1H2sk8V0fV21BY6VVf5XUgeeGLbBb
b5ITcWCzq/7k5CojDg9R8HxJ4S/YK7zoXdQHVv706iO/DRQ/3ATicwzarOeqLtBy
W7Uk4Eeq263tpQn0dSgK3P9n4ziGoI9zQZmt2z5W7sXJ+oh/v+1Mog04Iq6CyB0T
coLOCWPAaOBLiPt9tpLKWUOeVPAZZ724uWEOlwDivzrDwWtjLiaTHaT7ZJCOCcnR
8Pw5/PzlKOHIPMANLZpZ8HRqNCGapv7cuABfij3fiSJZsTCG/qK6uv2TKTqjIecZ
G7Hj2mJKi7r7N85soZWP9H06b34sTID2cLnFlxi7vIU93Nkje6so1HpVRlDLTn7a
QC6MvK3g1j2pwcEwFz6GPESQS3GhMxb0tXoun0myECBmE4q4FbCAvnObnCEjZRnq
HTBNzJ+BfjFMltQPs63lgju0C57LWvM76cLbY/Kuh2c+jp2OPtgXQ6hYqZimFF1O
GVTj+VYa+0a7bgY+NHIVS/J9U5KQBuMFCImqqvTYj98y8S8ULgjYsDH1gsV98u4S
tZFUZpGxtDt/os02yCCRP/GZBPQk5OnsgEKqO1G7q3/TebiieT563ke0WU5Ua8bx
7Gve9Coc1Tubpnp+b52vtpzvfNuVbdk12ndHp2KSco/BCf+Tq9GBE8dgCbWzN09F
zAA9TT32vCx33lXpVT2BKarO7YKztxAUvuBg8/Dqvk2oI2nYQExNxqWUjoTLSxPP
spaBKR69qoY3sQLqVVh1IRi3y4d1cvLQFxKH8zkRfM6KaFhtbtMggzjt5hiJpQ0P
4oVE0y3fxUuv5BFqzSqCDiNcWgSG9FXhNEJDwoZR5A8wqyJSCG+LhmnPQZnwTaCG
KrR0bSeUhfDGtjmULxSitgvilaV3jekjOoIqnfCzKklPdqXWODdma3bV5/1YUCT0
exutrIkaVkHP5kioKTGuFSpqPo/CONCVYyCItC7ncCBaYGZRS2RtFZXImyI+On7c
FPJ6XLfrdSKrLHqC3+u7hTEiOYLsUj0KVZqohROXik1PNXdHbhe8Bz8HByqeprmT
kd5dZg7ssDZSqoWPm8A6G29PIXw0Jb68zUXPftWXH2HkV+MWwJXpZ7OBMdlYOLU8
8V97T7JiiRJ7FEkwzidvTXvU69ztYbnQKc6VWZOvLUTE1FiyOqP/BbkiL2za5/Ow
xS0rpQt0A7F7SZg//kunuXuNPTmdQFxqYbggllZKyH+u4caF8g6CDgq76+KrZ4NQ
Qu77mKDbQc4Qgj5UaeS8dqCId/Dikd1BxnsLeCy8dcUX/DV9thwMigATwjkZyQX8
f2o9YRBwCIl6pZgs7VeUCnKRiBxb9mtdy8p3/PjbkdpqaW6BWdLogUZ1TLM2dZ/6
VWMSGPuq80E+jY8D71vbqVCwLdSTdIZtd8V2DupapxPMOuHKBMNOCZaT5eTJhoLB
0UZMoY3/+IyEbC8HkuVcOBiTRJWu/qtzfUEQjUgKRfRMTbidG8W1oR2wUslF/WGX
Y8tJx8XilZQ+DBer8d2eN6RtZMFZHzq9UW6NluL7FVt9eNlwgloJzX+BZ9uPyXXn
933O4pDkd52yMoOy9HRHMkzmAlapgmqwf4qVfhX8TR/l9gfF57iwbWi9xClXSvNP
LdlyG+kDLQX9EH/kQ3PsoHPgJ6ECEb0aI7vQhaeshfsW7hatAlBdnoxkcvBjIRot
Cx5LFV+zDAfqSllOwXhr7nDYIZ1Ym6CQOZ1zV307xlFS3yQE9yTViF8XzhNpP+DC
5iAGsQIvEwEbRyZJ9fp9ogPO0bmTpdHp/3lZKR/3ka8WA7nbexjgmefTsBDfhqSj
1ef/EiFqhMI+74opnSW3UVKCDvrOYj28tiEO7Ec8OU24kLZQ9zIzrqofa/8p6Xd3
BLmLCh07XX90EEkivky1dBl9BcEfg1hJEXeCDbtulmbbcD7ZzoenLdEsl8my6sop
CNsoRiQgaZiOF2Q5LbMl1LI59brk5N8g8T0YVLzkmxwDopgw5zXZNTEgDEBDnBXL
xQRSCxBLuW+1rrM4stPTqZsdzjSavaITgsG3/o3HhljLBJwUTtMIdyeUD0SUmP/6
Ha5d+3D4/h0C1Wc7gz04034l/qp+H+tmvPM6BC30yGTMTn70Y5mmWUdESbYcnmbr
K+ZwXwWx7VqdZIW/omRFDenA2ig8sPwGFNo1nQ1ELq+KeeIecbWjT9MqBILWZzYG
MSAtgdRQ9xEttaQriPwmozZRwlhDId0QyvQBB2z5Qd9JypRFkhaO1nJu786k3qP+
btyWBeBWeRy53MxaVmU7+kWKBWF3D/6hgbkE1pL3nH+m8iEkSU5Tw72f/JMCT2F7
y6pBfwVS1gzgJEClCsF7sco2z/lJLqyHeq/EBVMRmuzZtHP4Ad3cClBHVE73bsaJ
oSOj4qlzSAjAtQyH4a2hNOJ96Rp/6Na7DuST9dFpg+V1VAg+YbejKu+zkZsTV/f4
Z33xqACXIQvCR61msWCTTvRWK85vhWH+nnP9Q+AfrbLxc4TFGEBD9DXSn0nRsfxB
kZJhaQS0zFbnSbcz2r+mZIWIoDSuwvoQ0QPPtt2FR/xp/Czm3uQS2BIbF/kga75S
qBa8bv0e285Xucqp9Yq2LzzrK1ZsfvcYWI/hk7JKYJ3G2kVgv9BMzHr3YiigU0Jz
pBNB0jzLaE8wLrI94R3lJrphLhZ3G0LbTXD7vZldbp/vR5XyhLYGGMHRo2WjnSvD
Z/3parGKB32v3E3NP+Ta0kVatpnw/eA/xCG3/LYh6ANJTINPXJKSQ/jIWkcUQ1Mk
ZYvAICz/BQxehiCjRRdvtRDemJtA2T8bMaEdbc4yVRww/bb3eFEfoP6r3z7Ib78H
Fcoflji3EkCaBc88YKJRLh6kPTXwguUKiHD/BcGLUwxQw6cnTWOpGdUTQg0edGtc
o3uwQcWVB4l2mbBUI1pQILnJIuSqjiDEVgXfyNnzOMPGZ73XxPiCmVprlgYEHvve
+Qf5U5BsOH9+PI1k5NBger30GFKKJ/NuDXwkjafm4X++gNIq3pW+r2q6goIjSpNY
TCaZBh4Do9MEso7VX4ff420nPZRr7a5wzs6yhxk+LhLQfZ49KjKPd6eCurdhtpvV
JdNdUdIRoifioJxj3BVws/7dEvYgoxi++jYveuAOo5+y568IJmOEvGOVJnxx3Y7j
8rHXqV77MahoJdN1d5Ekit+FUcMskq8qItv7Al17CumS7A++qsKYmAYkpVsoWPDq
gy49HdplLsC3Bsu/cxS9G313GM2NXCeDY2HvI2TJ7xUf7nDxd4iT6a/50iLJTLhY
+0NcREy8Qqh0fiXmOiWAi+WhRHXc4e+c5ST9u3mghDBu3vo42nhPXmU++lH5jvFW
/nvMiHJqKkgGamidQtIKVAtDZrV5lmH6Oarq4wH3DDlWNmiXOMcod0ruBlMqzv5c
Fk8dq0sZUeNT6l4xyuSKkHOVMo8DnPVCUMouMCjbRu8aSwFIDmv4ufrR7T96dIXa
AWsmTL4H3y9RnJub7nzosYj6PTyQ6pJM3s/bGKIOsU40GbAGYHtnymdL8cD3dE4c
FqAbN6TQylM7NJPAsWigFK/ms+do7uHLs5ztr9YUXakCWrpJWmP5aREse/GQoCuF
ZxduetO74LAEfED0MdTqN1Lui7StjWAAVmO7+bkhVeXzPFJJLchxOP+IiyXZfJ0C
UV/3QAebdFxbU0jewVyawkCQOxv8dlsm2I6Tx/EPrXn4DAfuUvg1gnJ5qKjMXBfR
6dQjVpS307QymMFlBtJSM/vc4+mWGLnRt//Kqkv/ssw8DmAsRAjpKpOyuLez7YRL
zuaJkFFH4UHobgyn4yONKnt5ytkHpya7edZc2YiVMraeKOjIZewlqkiMpMPRvaDI
gFi25HrxlkmnshDsgDWBv52wMAKnhaXN/3qgJ3favtzBna7M+ydMMrWdmEatUa1N
UNWZsZ8HkSiWVy+ONjHo5XkWdh+DhvLvZO4euD8kKKo6x8KD9jVDJfMnPC4GyY1G
UX4CdZ4nHnYW0T4qA1iP6KbOtR679SAmcTUb+qQfeqoAPoeaubI4yxU12e9WXr4j
nx1oYMZyqlQUAkLayb0Bg96taPj+w48zAngKii74UtQtpGZj9ELhqXvFhjZBwz91
RWJO/hV7rLet4icsxfXfQ+LBDYzKTiMVAcqyIWa2KE7N0b8WGo/KfS9N+Um9RxGk
Lp2GYdQVNmVEU0IdbPkqW/TPxg12gk+GNGuylVwMIoGHn5CS8SaVigM5R28M+6iB
ELxjxborWNcVmwARdc47xNyACWQZwEMYoJSGlUVtzPCWUX8N957+347v5sEos4G+
89aFnuMYnkGe2XVN0+f5GyBBnVjpeUUyPQz2YPc9z++emMaxGPnzKYe1Ivi5q8js
H0ZrDD7Tgju3qii6IQJuyTxNE/Rkh12r7sK5ar1yeniJGQ9eqjH1wkNoFdEOUjMH
IotQ0qSNZf9SO3GCXO6FydalVqODPvuMG0pp2np4nRyuNRXmva3dqxA+6r4Ep+0l
6L5F/Z+ggOrvheGDt8yEhpPaHz5TeLzMKaV+lhHGiQTFcc0NRoDnUwTltITtFYSY
bBBVADPjHySUQJKF3OgtnsgG5RdJmJB8YhuZHYuuTD0qvZbyARU941WjzEVyfPex
hXY3ikpx/TWo8cIFYKo4qsScjn/DHwBcq3Xf+d5nhg3+PSBgpf8fby0utr2NYrbJ
aPcH+BVGOCStjzgr3MqkbyAR05ZKT0QUQRnrmPH5srVW9WjgO9h1TGa8Ht+slOaN
pt0WiKKb9be8Yzw/WaYfGsF1VmJ6u2TFiODzbQTLRmneGc+e/38b+Y9TlCDinmhJ
Jhdy7t73yx0aVSSdWmXb35Hh9GyaSnSUFUjlIK8Gmdz4Z3f5FnmWm/FOIlSA1YpZ
A9A4HgmIzb6kTqiyA/KWfDQK0CvTAvjfpif9WU/3CC2ndS0UkNGWOx1L26alyZNE
Vhv8SXT1dH8Tpga+yKxTkLEFReg5dV2o6KQNPAd/u0RVwU04W4XxXmC6V44/Q7Co
Wl58unFeSO3u46zvbR5TqmS0zeP10+BExL79Vegibj9BNk3om4hn2j0Tt1b7HYEe
muZONw6Jb7fTVinsElnIR3kIiB2q5sQvwwRSryekhS7FT+E3Vzg5Kttn0CRb6yE7
1j3j4+JbobBRUo+coQjuJ+LBAtHL12QYgTxKd2kXDNQAo2HJVHBv55dXSs5zEcG/
iImegSVmhnZ/XCjnkmrVG8ubtuhjESedZI8bwukOgy+DTFgkSC06GOfwvwe6OP9M
EM95ehTzyE6aK3uAS1RNg2c3DA6KLhS3Q/9k8O4mT2kif5sJndhJ/gqoc0xrUl0T
7lgFU/rij+yLYJuMNfbIgIAgHIPwecwJaYU7s584JZpNshwJLVXWRtz1GuQwmYmv
342gxUN5/tdnW/xE2CdB8JddJC6JdvFT/yyPenu8+qmYjv1Roz+rnKPBPhenO5me
Vy/ekSQYnJF2P6tjETYSWaDpyYn40K1hg4lx889oIsmBJu+Kt/p+kKARslhMsJdO
wNj6Jbz6F+0cL/VdbgVtcLOUZ7pHcsSH0FkS8k/vb8o76OJWon+v4h/OmNqxzuBp
9X9kSIWdr/5lZspddE60Tc8WeAdHwPn2skAo3iVu6Ate4r8SylJzeO5vzcLkDiif
jcfX4Em0o1qrM4wLuyCMStfNbVa13jLVmp7J+4BTFqrqittkYzhwqFd/5d0+oBda
keQgUYhri8Xx7h1hcedZMp0L6d9sFyyY2RNspfw72SCnK4hAg0yCl/nEaVnmyYiZ
h4qn4+y16eidQQU8mZdblNAhgAMEbS6vrd4gG76SNfDg7FDAi0JoPN4O4a5/HCaX
c7jZ/bqlZTFyBddMXMd+DPrkzKcneUviNEQS9KsanMP1Yat6VserXSQRV2LFH1Oy
E8A1C8yo41Xeuwxh1v7ns7CNeZ2Ctcnfif8r8vy0BLmM63MYT6T60cKIlJLDlMNs
QEsrC2JGvQ/tYoxLU0r+ON5k9ZHa7TCIg2TdNiLlExEnHwtknbGSdfRh5EmRJbNH
DxCgPB2EI5UPnbw8uERekwhQ785VICkbQULW8van/+NTfRxr4Q7r0g5i3yOseEzF
FrOVYrzs4n4RlHIaogE3Decpmj+gY7JrGyydx0XBSqNoh+YDYjXVRqXJpYFNQZs8
QNIkR8cJ9fnw7vz6hV1LtPOQlE/Kr6bj4QtSNVQ+Hxn1zwThNIddItj81j7NvbH7
7gLmHE67hKGhTigIEbBiGSRrTEcyjRD9xKjB9WJg37He8Z+jkd6kbbj2o6gzBsTd
f2TxAH8RHiM+6fQUr2ptqMUIMvW1iSJEAw8AlQUoLBfADMVf8U2vyrzcWGPZRKRS
ulDgnYf+Cbyyy/hiOQe1VIL6/TGXd/ocSOQ06vyXWSdVLxtO2JHT4dprIkJoP1K0
rw9NEtLU1M/aQWM6a1O99U0bjCXFrH+32BbpVDZtUku0WuO2gRujLW56slRQRDx9
TRhwQvbZmb4jBVjIGJgWoAyaKXJu/25gN9meTaOwxq3u2qr6EIgtfUBkzwcbLJY6
xPbViddvdS5pJhD+TpnvqCWbjAATeFLC2VpAsZcdXsIQ/Gt22mr5bBLUJLFxJ/Wu
hHEdGXSjuHg5c7cm7kw2AataKczbvJ0c9lEmdJgCvPtNWgzZ3JG4p+6QDcZ0EYZu
Wbxs/NriMQ+cxFI9jIPx6ppKTt4racP+quKRWg7zZfaU2FyqqVULorKF7BmXSHCv
E9j1hQNNFpvBDwFxz+JxWcqggV0qAn14/O0YGfVO7hAA0GxHDDqK1C2t5ef2hpSL
Ve0NhTDbGOJL2ki27yXGXH6SDlRGkIG8GQmR39OsRz+XkQ5dWo6a8vKbGqU4wL8f
NZvq+6m1xKogpRsBr9fJ1TayQZ1ZzGWs7gTO/anoMSDcW3E4oUaPpfa+p24juQUh
pSIyCIhqzTmBGFDOPJr24i0+itMEuJDpuQGjLixD9IywMdBZgA0uF03dmbv46WEo
vwi3Al2QzPZzv7tzz00SZbV/3EkvvRJ467hJnDacsy5K89Eqxtl41Efpz/pRNYB1
D6r6R6QV+3OSzOa4TO8ze+ewLWKdUmAsiMAAgxJ1v5hJiZFoBtx9DvXZsRSCqRZV
ucpStjtfyxo/dri5qLPqqhj5/8G+pVMiDwXrJ/84yoMhggQKPUPanAusrdvAui78
5f3RHF3YDJLWpPWVTJd4pzRog0Cbv1GEAaThCdTAlWTLX/IjXaBwuZ3Bdn08khbV
bl+9apy6VVcXUn5frLP45S3nPwf0+JR2L4w7eMuyMe95K2kw0krm9pcfHbob3Ft5
lKcXH9EHZXXd9PSKEGD05luUYCY5J/91OlkGNzig5kv+QQFsEm63TQrI7FUUEMap
oAosq2QHSW/04vGFp34OCCOwsalSXwKlD/lcTSS7/eWVRyz0Ucdqgn4Vg3abcRWd
v8UNFbdlfzIwma0jZE8ETrqAWPuKjuQRMs/FcEkJzLd0RfsnEiQ+HTLxSqHkLUIz
qxPgBwnLZk5P1iwoWOJcXdw1CxOhPsiNC+r8tZfqci2vBlcc3rLjpUvTOFPT+LyG
m/1hYMln802/GbCyzNgdoCeL6VCe3Vwo8nEjbuxgcjupmazMqmnU3Chm8lzMuI2l
tpNX0+C4bHh6JpOibfmrxiDpD3rRT/bjziPna+HjORVj737yy/QIK/rYRAvbsv64
TemYxv6cVnsQEsNusGZW4iXymvN3qAoyz8e/2rT4USIKSUU0XaqCAyCCfLxv2hnK
iVIdjw/4Z7R60wa7egEb8uQBoTiMcAAyloFCFab9TgdHJFf1mhNjrvqugMygBR6i
bkAt4MPf2a4rv7dC74umi9snP3gbpG5X5LZ5paCYfI25wMQFCOLMVSPWkuS2nfIK
KdS1MhfKatL/Yl6vraLYBxdQI8YIgVUpUrmjVv+GCWu0Mx+paZxsnaHDu7/pixJQ
hdeRrob/3sek9BqlGzJeJYGvVuhwLrDScRoZXpcHwOhBzQDidM8eHCb2lzWydtM3
5Nw5MchUoqZDXqYl5zsRZywopY2KzqI7GtZAtvGAq5oZK4j3IiVR9yQLOzUnTzBZ
b8lZJnVXKcbnSgHeYFbHjtth8DBrkGr0FbdDYT86AMvv84tDgqAsbf+PXI3P1Re4
HA2lwkGLI4XcEJDn+5M2C4jQsUOwFbJy7+eDrxilx88tgv07lhex59JTWDTXE/wS
3q1+oyeEL9/sn3hBcwxZf8c+ALI0TcmlbfGews/DFWFUfbuE2r6wJF5HjFw1aB1u
OiYq5fB+CPdXjyXr5J2Tuwq1LI/YTIcs/dFrHcD4QkibtjoSzphDeXWmd/Ev67s0
xbzCFRrdehWY0QQ1QU+YLakYdFu2efhN7VG31vPihYIF+JaxlRj8cusAsH1C+Tnk
JNJP7zYgC/KWAmxWyEBx1I/4asILp5vW60JBaZnY6/NcMlrgp7C9hM1PEIfpmjS6
MaP2zKbp6irwficX1LatNpnwm3fuXkJWCjRUKQ6Pp9uRD1U7Qh4912JA3IWZ33AY
PhUahRGoaHigaclh0lRH/KKWU3FujeEg4BMOkFumLT8CswCN007J8A/7Z6slKrqq
IxEYAikMPb9Khg/5qVSRKeuoTQNAaA8Y8SY9OmQwlkIBDhQRaEsLK6YG1pkfcgw6
y3gNEq+E6opu+4cdWtG71lRvOzrzTYhzRiS6mWsblQsBi6WO7zUM+CntjpRn+fhe
YRT/bKe4UVT/Atmez2ggfScz3waxkDeaaOPspcjUmq0uiK/8WwiPNIs/zWXB7/GC
tsx5C3P2XgcbCZ+hkV4YGrrTXKDO4tMpCCjv34NRolmzYST0LnxGfl/iuYzbei2o
pLTftsswUtxnF+tziXxeJnicRg9M5aLS2lvrioEEx115pbjW9jc1ubShDtDxRYVY
5V330N3mKSFzFGpeWPs9PnCdsIA6+0kyY6qp5dsdS0AhEtCRe3p/zZZm2nifACQw
+Ch6oqi84ZYtAlQNpZqGcauvtmL10iyHDe6e8PlFZl+WqRQxXzZvkFyOC0wGT+/m
o+EflfIioHlZjuFtmsnlgJt99qmQmJG0aJUr1OWtOKJkrsXPEntEoX2aoc9Vg3kA
ahYOvhR75MQdVHfu1aNQGJWgWJ5NYA/o41+M8WPRKduqNuvuI3JSLrF8o36mZKB6
SJBTkbqi8HLPdtEhHu8NYi4hSzgDEyuRFXtxY9zsf/RKgelGjPHguKb6+v8Yh8Ij
Mopd59GuGoj/Viwd9WALlXoecTU01pu1knPSY1BnfrEPC9qhFTRCyVq+NASKPf1w
+P55BIzhzYkdqgD3H63oDFg8+nQYpmRorEzhhNsic+fNElBK+7vLtvYR0wVYc88E
2SCLGEL1eflZO93c5BpjHmFA+pV2MIwVkghI/EyZKY0Oj5y5a5ADn/kZa7NBU8wM
IVeC2PuTdHJxyB7OEECpKQgdRgGI2ouhkVMen34LpLy6WlrhysU1qcelildW8lbI
QuJi6FsOMlSlxLhHYj5oNE8jOhKD6zLRVhjKaZ1UkD94Tl0bZkJeGCVRVlo+ifAH
s3WcLVY0gE1/ZaMh1q43AawF2OgJw+eJwrDYUvv2pr8y3BvPDWJVq/UELPgy+MPY
WJR7MwL+tNxLmrvUXQnaNKjD3i2T4wgOb4XeTX6yD/6hSK5C2wWh9dGRfUuYoTAO
H+r0ayzBtgYataJoJoFPiI3+04Z0c/7+EtLxO0mCoow8/3BOnqB5poeh0rkQOQfx
FRBFj3BezNk4kpgK5Ka4a9WeoseIELvQGabJAml7HyvSJskfAcjawcabUWi5cEHo
CgLM+Kl5Z5WRJNDlovka+p7y72E2FwG9acku18z+4zt/bSEbBjN8712Sb52OXcNn
z5XY1IXSUaMnmeKvMfhTiLTVtaj1wQGgpGzDqc7IhbBi0E3BHLslsinPWI4FMe/7
u9xZw9rTD0u6oIZhvSDqNQYWUCJEb26rUYcxVOKzEPLXA62jAE8g/ZPxSp0OBr7g
pw66Dl9Mz7dYHglp0+ypQJmKXEA+jVRuN5bAApZ25CJwCopWvwaJPIW18A+9eVsN
kIzAkZY/pgMV4yh3dOIG9yA6tDxE+SXPHIexUWaRpyG6wjxxFylsuLGn3ER9l5rF
3z/Yy2r9XUI7XsO5rHJ96UQRKAvBsBtSsdZW0LQ2gNAQP7lgYqIM7l7zezrAp3yj
/OrU0kemWTnrOp+pzd57I1f6wfvWVpnLiW2LhnED39AC84K3+Y15xkVmpsTX0QAr
DBs/6bbrAIjOw+4mAVtbhjOv6KVfAMLBLgid/eYXB+K+/vnUEipqNmlmWjFIIB2D
VpseCycEKG8UJt5LsIHZ6x9R6QyY/scTI+nzAlcxA2HUCgj6e+D1k8Ro8taFvnm/
/QvaX2K37qjfgiTpLpJt503KIoM8kY1+ZYupMiIS4eq0Fkd8v80VOEu3e6Npc6sD
2X++Z+PAX4BCYZeQVScqZdHwJ2hP1AH+nTULUBbqaKr5C1eBst0MayzEpHlyvMrk
TeooOQJZ2ir6KgDHNwbmtK2DYteqrszhvDHfs8pyNZhZ3wUMCxd/A7kP0wx6+wBJ
yHUfU0DJLeKxQs6DDc9/6KfkKuUG3e7cl5gkplf7eq9ZXWFFwcf6JqpdaALDnibP
Uty4ivw4o42kEeqalsitgCLxzSTEd8iIAHtIeTNiWtPzTnNFa5mHD0SVb/+UpC4Y
UywEge/RU1jr0UFsrxeipAgrWqn6I8//uHkwK9AVf61jrjvyMTmgxc5urJQaPe3j
eEWMsdoEJ0MUzJ/T18oNXCB8+Fy3RagVmFgWdPRnYC/8c+E8D0mOhC97LGyX+FKq
Vkdaw4qR1A3oe890VfVYqBjAr7rOCiGxggyC0T039sHFbpRQx9g8r4ov2r8nBTLr
0J4g850N/SdaTGc9lrwjlXqCYqSIk/t0p9vtMwqYRYCrzQ9PHYrOYNUT1+t0NlGX
FZEFfnPf70DcIywOhigFaTV7Eop9vVuV+JvN/HymSsZwwcQ2d8mRjZtIa72yMCi2
ilGO5CgM+PGpISKwSexDrGdenA6t3ae11PqGoH7+dvSruzEgb9UHpo0VCvL/DE2z
/6PdUE+70dAviKoO+e5f0yytS0/TjwwvoCCtyJhemHWLz+uDc4ShvOW/6ArEcRqq
manwTXUrT4mKub4bFqLxtr6wEC7ogn0bqlJlUzRiEqKsjz+4hyThOr92ua+6crB/
SGE8q5Bo+XhLv0q0qMmIe46xVRnIZYe106LEDm3HAFWc5jT94lHw6N4q1wxIrBn/
6+U2dS5H7ic1hJIZUlIkgXNlcAV6OI75JkyxyEAQ/Nmrt6yxKpTSdko9RvLTfsDx
3nYJ6sfSzpf//CmSEACpHLt29pg0/9AwWjVqyF7SBhz3x6UYOXBlSZrsR4Tz5rC7
aXLo2MqSW5g061L8003HSaAAZhBrN/z6YDEWpwdVE5lBDxLrJ0Bzj/rge5shVcpD
VuH+N+Va3GcDNX4R08QwaPJoJ8Zmju/ZKsSqhCsXD69HivAw4XEWPY3d/wPSV1OB
SqGILpVpZ7US36W+K2BG+SCxq8PXkBe84M64hJZjerZ182KmHnDGnmxYMj2nb9vh
jRzomLmnVySi73RVGJyqEOuppfAeICJGOVM1mKSt14Ld6SKO6pphBfkWUodMb7AP
sHOmpOUbp4/bofFuzoL8crnqYICrMMYS3vnDWWAfnEE6regFI/IuUJ8Cb2ZpgQca
AY/fHBeceEMrSibQ3IIu1yIjzXEFAB8eoxu+Bqj63hUf3hu2SW8UbjLjC8+vCDex
abwWxiz1wTwKNZEe8OmfEqbSRoQ4/jDygF227NRtU6jqa/ra8vNgC8JA5vrA7r0t
sBesf+QIy80ECXrgLq5+rNZDIih3C2vAKfnfC8dklL8xOHh8h4Chv9B8zCZHycgM
CoNwun9BMhTipC92ItHxGamTTQo3iVwSmhRughNcS+M6w0NojHghwQUzy3pTkVyF
zBCPfdhDx/7aOhB6thMD8dQ59fp6bwMJZm6BVxbHTH6WEWF2zCuma9XnY8QNW+1H
KCy0Gb38SWrxgSYSc914a3hFqcS8xjga01viJUwid1DBaDcrOxbLvfuHnL3MNTEE
mmk10kab47VXhuu9QDrdMVqNB/D0pZb4pjv8q2JZsQZp+cH9eDHdxH0xHk/8W8cl
XiXYStHH4Rm7yIAZUHkKyROuEb0JWDrglXbdpdLSTH9DZaf8oJ2IfoNPg1XMfEVC
U1ZeSwau3BC+SicQX2cdXn3LrYdJkVUIT+NVQ3pO68SR5mckXxg9lfWl4qGDsund
gBm+09TBnPG9K1YJyHwPAYqF3hADPWaexvFYtwta7zdB+mwfjR0wMyCVchdqVYGN
Tj+Cf8hIRbQJwl5eJQBtaefdJBsQ9MLGcq3GkhL6bRRYAT+Fifb2GhtyAlFKcpqK
lIaYu+swKtsLJyx0/2lLWQrYRyAQvyS6B95E/Jbvx207Fvau1FzinbRAwe9Kmdr4
j0n3NyM8sRq9gLTV1RJXJcDDvCVxbEvB+ut/IoE/2lwEPHRSFVjNbnX+ub/EnuEm
PMmiIZvtXb/ViZiyqDs8+Sr2AGIqw0UIM2UX9j14nTvmELOyy8WdH4o/FxM65U0M
DxUJajKVO8K95BBCfG53v5gS42gYhkdvBiaWwo4j0MqTMw4i0ANG8cVKPZmqddf3
+puKCIaywf1lYzZ3WHDnREAqNxDHFSs5pXKyDn2LPME/LmQL/Am8d5ZqNd5k0utB
R8gQa53bLiziB+Hlif/rwC2FP/Cy39H5MOaR2WdgX4rgCzM0qRaH6D5MuF9WJRm6
saWPLqiXaZF+uEX54bODIygx56+NGvdKH8CVhulScZ6VMonoAQMyhTca0UPTK0fP
aRw/r6eIFVpS5FwIijfXbNDbyxswegzdWG2WoQnESUuuiMT4MIasqW+ARuKALEgj
pJdpiATJT4XGS1wwjz1h5LuN7Djsnd7oCxEwMOm+S8O4gfGHRpqQF6BuGExHJREz
1rUZDm+PZNVk+kom46ci5zcbUeYvFXNz4xxXGQiwhZyPiQCCQ0rvrEG9xNUnqCVq
AihfdH9Zh4L+tg4WAIPr1slTnfzDKeyUFa3SiLVsmLygy8tRsGOb8i2Njtq7Gioh
QiEnZTZuuRA5h2qsTaGp4fVOFU4DLEIVzjwgj/QNyfc=
`protect END_PROTECTED
