`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4wbIy8PwCX3ygERPIy5pxZRON19PEBUKpdn8HrXMuh6fia39V13x4RBBwGQV53b
oR9FM1qwrbaeKoPudbs6jhgZFPquf0Bw7ExVMGlX//9BbJ0+wvz2vuDubAeIvghS
M4OteqcvWM0P5lIVuksTM3mEckMA3t6UwSpNVdS7U5GRiCc9I59twRRdJxt0fYzd
ahOFhsC56N6EzoD82jDk0UhhBGQezp3TqXQ0NFccVh61K+ewx8qNkig+biNzb2Hd
MbK56P0OdqrY/LOT0SGcSqgfG/uKlA+mIfwJtNVE1KekWER1TEW31i4D8/bzqA/U
yHvjWfVkuLcjDnQzzss7ZuRHONBY2yowh0uToAXEcQVwCJLE46ALl2FOmxEnk5SM
OuamTAiUDmHYPDpxfFrwdwljoaucXda0OHXV0MXaIE5hzUvNiaPOCfZs4PLludnV
qnHFJNVYyzIW54qeLZ4Oo/PlAzMCWnb9eiieMuSNFqXbelD8pG/STwGHG8I4GmUX
AMll+FlWSNwDEO7BCZahw8ZSIsMAfivNkGSrymwdVCEVJtx1ARpLCRE5iD/V4qa5
KPUX5Mg7jOKiDxr3cMKWYmWAqjZnv3GMC+VOYjmGNG+3J8ySmHw9oaJ5HVu3S8dr
nRtrA60gix+nNT0etoJoITsABPBCrlAJL4JAVOU8TpgqiBqkl8/CgEcNoqAtYJcr
`protect END_PROTECTED
