`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bs+edIh+hL9WjVOIeajaXJZaF6Vq46+uM1V/X84DxzkTP7A85zi6MnMtqU9ZWwUE
C+WWuz5ACjrHGmgovthf5E3IDCJLGtB5s0/HrdEDwI8yap1E9ROtJEDzDVmKXdW9
5WrZBP9hRJi4yd/6J+vocIa+NSllY/Xs1uVuC03qQaqfC3VdlqwgXh6Xa8BZJ7J7
TyOhJPoifuH5kxcZWbyGUAMqAVSVAIXSsEZbpUTvM4SS4kZLq2m2+LHsT/o+7CNn
W6T+CjDN1+ICNSL9s4pOxbo7YmHcPn8VLkJauFll+jk72TvEgcmstZ5FIpbV29x0
TppMl7VbFz5RyPbHU/KDB9hp++XQPqBhFD6G0ApviOW0SIK7V8qYhplHo89wmbr+
1tQodaoWWCCC1BQUS7SUTtkLCkn4arldkCRilfBkQAafucPnpkM+3BPkttyPvevy
JTfAD4PE3GzaHWE367ovTBRR8PgwQYEzfs0WmGaDrmO/kYr55YJNwn96uTlR0Rg/
U4JS/baLpM7IXw3s0FGT+JTOpDMRK8xAcTfK2P7hOHr0lOlTIpP2RMoe4Yl98cUo
ng3VW1Jxynnm6OUgRDNSBIxLIAyb7ADadCyz6k3TzB83xUM/FW9MFpEuotf5x2LJ
RfmianpzIXRMU7r/HJ/CO88jMTZGSROxM83AN+4DPUEa2jlQySQz79Z0eYVLCrvW
mwhkgwDg7svcrw3K2jTQPLZ6HnKnSddAiOYUm/HQaUgLAF9JJRuSWa+LK8KxO4c9
OjHdc/o04X5NPhaB1ltNvd5pVH90RQI3uZ8uJPMC/tktGNy0ye96oJgVJ43HTPEh
QHh6rzR9uJM9AJ4uUizjrL2rWjtmhpwkTXM9kgKrlAwk8fY+OHre9UZBWnK+jtlt
tH5qxSd6wf7SCVQ2iT6gK9OF0H3iTc/sCWhHoM2GzNzx/4GHMVfPIJzVOMpy/jrf
GvPbHjzD5U196++tYn4SwfTDk9oI+kK1jCaA+jMb7ufR32xd6jsS0LsXeilItVQ3
5N1Cu6mE3U7+0m9NSOgvZZCQmvo/iMCZBUzyQcwGKeUSeLotfQv3jHZMXUI7lCzD
3/X5U0CYfjRIlfim5LGRcVgBJS5rs3Epf0nz40Wbpa8iJg9K7kzbrC0LvDidvzjz
UJBlsMkEVBwOrBHjdzFKQBG/QFBu93ekT4MoMyCfyvGArUNx/exjio90/Xwv/+r8
i40ZmoTGUjJBwcHNSL62yZ4Hl1evknzFf4yXYeTsmFc6JMDG+/krE9DYgGbyzR9y
nYFxn5lGzYI1Rq7Ejb2R5o0fTDy42RkOoLz47oZyJFBonwgeJu4qUrhRij6twIH2
PwAIAhcrRsdOn8ZQdmfiUgmobQnuIztfx5Ajad9qTW4RDDODCTX2pEiuKpXbc2gp
RFFM6lwiIDikhecMqjFy5TkoZXZO8FSg56p+PurzjEIHsNg/GcFMXLqP9+dWWd8i
nPb/y/bj2V87gNoUsDnASCsuaah5on3wcQuPL0kFzFwZrwSDxmedE73r+3iv3Kk8
GqdaYV3+Iw8UIbomohVFMCAfnjBsgTuR/01sBUi0965x2NicKQp4rOgrrNMSjPca
8jPQoHgfztF/5rKSpWTDvFk75LhWP0XeakZAtmb6g8HmcrLpT4YMXHnBnrY+v4Zs
gtG5wqHIY8HLYkiHp0EnbQ+FXG7j1KZpVM42Ih4Ti3ggw/vrr3P2mV2jgyLPbzLI
2OQcLuhYmJYRrrtbSg/DY/ZBXhq6eeSOVuI1e9v/Ylrfd4VNYzMb1ASl5OJ9bVt/
lFHgh2SEHky9/e1SmiPjShAH5CN6p25vc1gSkWwI1CZbXsa9QZ2pF0msWNf0jcqp
8T7MNv3P/eN7xdAaOsCElDPeF30jDeu+3IX3UnLaQIL3u29s0+6X8+gwTTlX6iD/
W4QAyyYddJ5MWrTNzxR0Mp38ZLON42EbPY9NKGv0Q4yFb3wur3a7E6F1BdL375Ts
bBtJBH5nVkPN3pHpXlSwFbjyDFH4xXXgYgp5iHomtXFF81Dswd0xDTDzVIa10k66
qow0+eIlSvO3JvJoQjSXntsH/vv/QxdQQsQDEWIOw/IyLf2ceik4Ks1rXcJbUALB
XdpAqrVk2SKLpG+9h8CA9Zi9yhyAdVVY5hDfmK9Q13USm+O87TnpJ3WdO5Uy5HXL
3aD2b/A5b3/1iBxreXRqltHsJqbrR+uJZTRMmQ2T3AOFe/KL602hJl+0l/FGQjHf
K1W5Grdw1Q9bTzncybS2PpCX3Mu/9lilPdMitmMiLv/vue0re8cmY19+FGb+tBTM
5xx3rZWgIKwfEvhzGeqFhqGCSyjG9bdZZAcotojJy6bh9VMTsMQAFq4YKzrzgPfA
w8VSAt5jBjfUf++0rzyQVXAi9tpSLd65xMD4hJ3sUd75reDpU7jQ2CEBIx97g9Dn
vHbgg/SJfRVoih7uMEpNbN56e2QE9j9jeQjU6o060gZWHDjArPM2nI8fOz2lyjMj
bTZnB17Z79Ivb16WgYjzPInaRb0l6P6kwvZN51ZkrQMTeLwobed0+CJV5rjAehWw
ahLmAVAvKuN4tGneQ0FpvHFRW6yHGdoRE77MqGXKOY9KiNubdbu/s1Fv0YnHdM9s
6NY6FCJ8A1kHrHmdtKza50KoNX12ttXhbClUjgRRKYTNKwIq/msY8DefNpycv4Wc
`protect END_PROTECTED
