`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqCWwRfHLVPDbNt9xcXfYxpX6knjy/lSEX9sl6BlhWXDp9UQJCpTtTnagddrPZ8Y
o3cRFj38W20uUcexJjfKeAG9uIrVMKSJZfDvPHI6A5PO7Rrw2KBIGy0SCF+BnQWF
Em7FZp5qIAZh0V5F+U8GsAKg2l7ZNPwWU6XZnOS/nM5pJNwEklP/Ov8N1dXk1ggd
y9zhcVg4TmgN8UVvA7ZiOnhx+xS44HSdkucmfv5+MYGa4AzTHfK4enWpQqIqkmjz
HrPc62jMWmPfWWCQaSK76Lqqeq/zuSxqyjcnqgi2dghDftsmXcHNqUmYKj//4A2s
6d9GgkDfHNO304wAKgcN9uBQKPmSg61MEHjcj++naYu2K1bJUl+z02KZLH9aNHRE
5PMRh2i/86vesXlqx4XhxRYJ7S4ju5htUaDfBf2RsbemZAuvygpwOgf2ZckfBChM
n1zfaxgkZ2BgbYr9pQqKycyHFNPvs3WL2jkptGiNXcEZbo40q+iBUO/g8lEKH4CH
wQz7ITekrbqLXU6/c45wv//FSVzf+Y2bZXIjwrP1JKSzIJxuVqUMm3SzyOW+Lehw
EnSmPcI1qvVyPAZhegLP9p1IeQIKrnhKqVNDXKPhMIo=
`protect END_PROTECTED
