`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQnkDRZXkxo6keqsSOiKpg7ctsFPqGUZm0hTswhGKSn3AG7YvpyuHwEfbTLyB0Ej
hOXkdCm6iM8bcStBGmjpeWArxqmwX5x56jM5pFeg1cgK6BKSDebjq38Kwznxp4wU
9KanxMXkt8me/yFLHmkjgSqdDv4rS73SjL//MqcYLadhv1/bFUdlzSX7dqJ4xhpa
1ji/u1JJR5FQzgh0QueE1nFfF+S+1wUz48pIh66VYlEsa02ROQJ/eorn6Owm7uxP
ZhahILJAH8mUWALl9OLNVC8u1S7VNRpp/KsMVAkfGp6yukAEaaXAT8LpjL26eCEq
O3hu9Mq6dJlNbhh/5SVr5x/PfkI+l7qn9uXsxf/u33QcI9gsvE0jzusl3nUYgi49
B+HthIdGdRyJuMD7VxBWOnCOE2+7brh50/r8a2jnrxMhxEl0rlIC3ohYZOkC2i5q
fdZJUFiPC4ke9zmf3AomY9Zc2TCqvhTJLfV8TXvon9Def5cONpLflBIbGvontugg
S4od9/E65ETQpCR4swkNvabCvtkLOGYNT4WW27IWl+fgYL7hTOxe1kjlWMw7HEnh
6pJqpo+wQcyUsxQzv1jZBMopRN1B6qpVf8LZ3H5J/bvGPT96zc+PF1nKRZWh7SQ7
5BszngYsnrqaV4tcVMzL+MHEc118GuIef/Dugq4gNz8H6+rsGZmv7VsF7Y731sXN
RpkDUV58T/xSl5bkGR8D9Y35ydvuItPb8l3h9EV7UHG91gLuDa4OUek1IoMNJkpD
LoTkJfPjrzRU7xVKC6HrilMP1vqZjiEouxnv9fhouPZbbqV+IcMlJH9Hml3AQz7n
n460xSNoyxxDgcuduvZblXW/Av4XtElOE6Dnd1Isf6DghhQGUXukefkcWJz+FiGf
4z7H/06n2P1xL0mSt7N0aGLu4CxfudGXhQiB6irutO46sy0ScfiRfAYFKFGjQ9aP
bNu7uM0S9+U59kKzJ7hpecZRd8hYSoMoRveLnDGFQPUg8apPHuT6UCT15UikFRF5
Phci3ASDEum2xaPiQsPpJgvo+n29oFxOBnLzjF4SzoUmeI4kxTuJdE///Cy9ug9t
2l1djsW1EgKMTUQNkB9ocgfxcDueHj4vQzXMDsaGAohNcjXe2kGVxTJNCIG9OVBa
6nI1z8Zg3GR4JBJfnLBCIn2+W9wtaE8pBd1+1x45MW7U8bhByi5r9Bv4a+zYiR0K
/mue4ZquFZIGQOWC8hSPGNCSeVWDoGbty7p5eAeJvIIfmtKx0Kd+lmQ47LpsQzJi
WkhCY0LgYKQEErcnJVLVwhQ6+B/QTMJrePrr5RwBpZ3rbQ+8ZpIOtTh3mLLj2iKv
0lpvCalksYZCk11wcRwJy+7lJXVS0lca3Adak8JqKIgiPIICdBgTFoDS8y/j3yCJ
nKa8GJPIuc+Acj08thA2qYBjQqNTDZHKo98n4OepB7O3T/J/ynR13RCso1PgJWSU
GDJ6PDeHOxFnyYYgRsMBXVuyObN6uDc08zGuInRPX1S0ustCPbKTWrhn14glAR4l
DxAXRLg3ektb0/4Z9emtszEkUIbL9Wa/N9oBpIOxgYFKQ5pv6HxiAYldJzXM2zCD
/dvq5oRyd3OCmzkrmRUb+Xym1UKpDqcQYESs0c+z1Nz0o500XEvNnoGc0OxaDk6l
mRXJWDiKWDwCUh0RCDQq/4VYzShLKEoFcaq4XDjiNCh81M2ivlDuIrb2r0PNlmws
F8iHSmdHBVYfY1pJFjHTNnG5w1DrDISiiK0jemY9tuzqKDDuhBDH3T1B8hD0lf59
U3Hci927lOFFyPmBj6LCJkBNCwBekBgK/kxok2Q6ug4bAB8RtCol6EERG0dlRLKQ
oODoYfnL4L1sYzsbLM6+odoThF/MbWRJxoAyxPGDdj/l55UXvSKfFGJ3By19oASb
CRMOFozsrfD6VhyUXHsklePjJ36QwvqmkFzfshy5rQ5KQQmptKZ4HZnc+1z6G8Fd
HSRbI6/skmbjpsgfZ1MS/QJMQdMkbr8rUGbgLG3c49lfGmtFw02Uo5AasirFr0o/
EfL+g7S0TXZfhXrqgBkrbyhdLWchx/DJQkGzkFq11Ke0qO2utiWHR7IbBu2rm/ry
VVSTxsc+lux4gPGqu7eJcLz7FpbSZ71Cs2QR8cXXOF/T26UZMSRaj3PzXCsr1C9o
22qL/FpYrswd08SPN4Puq8/hlVv7/ECOzAYfuD0gtQ2VCKQn0jfLObK460zHBv5o
4jyk/ZNg2rOPYp/pCkBtbWlsoeHiAZJtz/l9HQJ+lOfNNHcRIhx4ITDmUD/3UXTP
CmBYhXHNHdp2baoPNSY1Y6PUSiNK7AUfFjDty0tBgtd4FDiSHGLbYVd3FNodWRX8
fw7vKexe3iicp5zrwMmOY19CJKuPm7QmsmOLAZYy6k3b68el5KgfvZYQ3VcRzIM9
nH7cS5Emk82UmDL/dJYuNr9BSnA1vo4n07g+shLruxQ4xv/H0g+Hel3z5ZHO681L
9a30FfuZy5ITYcz9T5P/1KpFgtKd+ELtvG6g4E1eDlcBweTrZTfmwKXpQbjci+jW
mn8UoJt9DgElAQCnrhHVNdaomZ3yulxWkXa1PQZRZ+p8/rxvzqhpGEZvJe9vnOYJ
9hHiWpyeDXqxzcG7B4zstF7NdfLWVTEaW9LSwEPrk/7RODTK90PuQcpMfDY2rmeN
ogr//obB0emFXj1XFQUe1JCs5Lz37fQkWqQj/WVpPS/Xh7i0S3czGFU63Or7EneO
YGbmqxD2fbGfTVPV2RGXaKsaruXRmdXepT7QXZP/i7ljYSj6HlicbMsMinXEoyg0
5x4vldls4ysalCIn8/5tA3BQsEX65usQNzqEs6p7A0hAMDbZ1HNeX1skPeQ7/gcp
J1/FVjxt0DTiiEQ0acWrXIPIVEUYgU5pPuJ/2Sr3LDuJrze3BhxZ+ix07aNjAd+2
2E5OPdWzXexx6+R6nXH/03D5168Q7oqX6pDs64PnlXUxBV4f4lW4HTW90w/JT7N7
96lOUdDfjXKQ1hrSepr83/2+pWsSZEyxGR/WH+tddXMrMsc2nzQXcWtyAowUKq4h
8FYS8iVYz3qr2buMAeHEBJMWUk5IYMLuZa5JGqFJbC3P7xb3ZXaf/BpPLzxVqoss
cQq0dVzm0ZZyfcAYUTJ5k4VXwcp+QTVenx2/Y16rUdS2tgI5vXO8dRyG6LJqLhmC
kNGm3pCA1x+zJGg3QXbKRGTh197HxDPOnkWn8uOs9Z/03/90wClLrJkPFo3aJWMe
kRhnhvC+I1nUTClC+sjLcliLwWtM/HwCO/jNgcLeMyGW4VQ4QlpHX3SoAtANf4iU
FjRo9qUr1UwnQ56LpCoYLH7u72rHefCo6byvlfzI9i6Exi6GrlAiNbOxj0NPgq2H
XOQ2fRCRAvC3aljuzCdZ7IYPrv+xFlMgeniUi2/8EIbLZxDjjZtcXNZgX4Lp+s71
lIu7cYjzhlMHAaxRk+aXTHI2HMu3ammUYCL6Y6j6DB/gG+VwD/1GfMeX/e98jXBb
1kX4hsA4SL4Dz1f7/KLKXspHQwFXeYCugmYs/eKJNJh50+IosMZ+Kwh5+BZ6Nj8T
P4DI6cVikDLXvwJ7GY8eRi81Phi9Twsa1sedXtpEuN+jfT+zUfcqEcpOUJrIStOb
n2D6uM8JpOqHc1RM+YU/hbbRFRgWvfMJZ17Vm91ZbKoBRCBHvbHowuM0xiJrJ9XF
O8+VthCCk+pPy2nrixj+hT09s+A+RwPvlZHfTPtOjBKhwPKTTzqBRNZL8A396jM8
KXogu0AIBq1O5Zxbc3esEw8o1X4auHZSLD3Nf9d3501N3jP+Bh0oqZ3SBYeSxp6P
5luTWcKgDL0uiYN7rRrTz4hBKC/a7PCNrsyZAIu0Kpm9tKD4plSyBfVUfnwmL9e8
qkLb4an5FEbj4gy3VkaL7TryazRD16Z4igl5UoLKyo7h4IYNyf9hUapovkiV2jsL
m5GbOWmTzv+qV4RjGUsVwt2I5G3B3jouKMkARoWLj2NlmrHW6OT+HCoIVVNS+W/S
l3YhS6mUOone79c3zk3fAXHeqt0G/Faz57xmH/5pV0cLSf1FL+8bXZz2iQsORrOR
1RgIBjovBi2PYyhejiYcFnLiqpnwqkAz5Y2M36OT9xCevnL7S9pz49JcmAAHxgkk
GVHpQ9QaRE7zISKjsb+dAjSoKxkxDU1JxUpOdHKjb/wCuI1RXGVo4j/sJ7oPtV+O
fypyh7pw7Tr4aSBHqaU4tuJ+Y9Wt6JGNoM7KOgseLqNlRIvK0fcrEK47YIwnZfAp
UtpguqLT4EmV1OLUOTLAkyufcmaenVjLeF6o7nYzhWzCpk/0IfGUtzGWG/qq3nkE
LH4cTA2Bzse1ub4ixa5UiUy7Qc+0x0uS3CL3TaIT+DFbJsftcJQBe4lKFtD4yuZ3
/udZGrt10CQ85R8BrhmxW72dciw8uVkaudL5S9JPRKYMp0O2QSYH7o7UPzLIkskL
Aepc2OIr9md+ukZjTZEeOW1Nao1+eiMVLcsD3DvHA/L4+AIDH11hpOaeipPOTNmw
cgyYTDrh1vw1GssT3qwgBA/Q5P4SS9GS5RZ+hAiA6RFHWaiwRKldnna6kbY3+XoI
5Gex/HH9z26djgA9aMEbigJTYmwy5CUFsYUFvJ024phZkzskMfeYbZiQHHBAhkqq
VoiFT/C/17KkYZGNKrWd3WMVQjxRVXG0P2X0WD+VGM3MXTmyvaGMKrudm5qCu8SO
4aD4QeWuq9CNskOoUgqKBWHuCHrUHba+E67qxp1m6xkIux+DmPE42KsezYoBMDsv
OQk++VsghptMLubMb3YPUsDlDAl+YoDOHZgsR9Tx+gHxpmnE0nNzSfQOdCCXwjTn
q6DrLf0xudivCihP4Ix6v/heiHvjWbfRQRurp2UZYFUDZe5twRq9kkh7Dks6ukHT
KS7JSmKE85Cm/MgHRYywjikXibK2UuiivgrH/WLCJJM6SbGMKs9+JeIA+F1S7Wmr
nJ0O9XQKEBYDiHCkbkw/pvDzCBoxlistM2moDIr+rc8gurw+Yp39DNKVEzLjeFXR
EgpIqF5pD0SGzz7PXAsopxxsDjMeZIPO40LvOgYCqbokLUQ7wceMpF45ml0n9f1P
MCcCmaxIN0FluMbi2Zu8M2D/WMWnbbeNIR1rkBrXnJDGUnmajVA9h7LTog52ZOTl
F1bMo2wP7zEvnuoBPAGTBrWEGjqUr6JZ76Vs0OeICxm9MtLiXsZz10VxTTtP6TGJ
MU3HGMVuCds8ahYi4YshBs1iHmNb8PNeVDFZPrXzsIfdmiX7DWRcrlac8YGznNZ8
taJP8cmqxKDoJIHztOXC9Y9PDi9xGZZM/++n0ma5Y53hJMS7IfyWDYvFCtsT3Mg4
fZ+1uFgxG43S01kS8QU4Z4FuyvlIEoR3wleb5Q4i3ZKIvRb5HVzN7h1JN02DYrYe
pNB1EOSmmi6H+HIYRcn+uLcr4G82ceWbuNFUD8147N27jzNahbqY2gFsxMvzouJ3
TrEsNMJqKbJHYSNqCUlYBt4ykyrf1Cu5YyKiX0WtcUzDCRatRetBROSHOCX3Quu+
MKWWtv1fXnh8ypMX1rbVq3PVaoOSfsXgtpr2+UZdqDGIhJjrlcm40KXwSrEZ+qcf
6DG1g8StI4O2aOozmiLOBg0ifNvTSuiHHFKuHVK5gQVqBpHHUJ44P4cVtJHc09M5
OCToRC2dj2hh0/Vc7+CjtYZChKv9IIgOUAFH0kj0RHUBRGbc5lEcXKiHoh3c+5H5
iaZ8ze4CJ1NHchk5qrRikRnRTF0IscFHXQcgflqPi5nY81p0I5bq8o3tjdIo7mLP
ZSPAl0kTs5ANx2To4Na/H+8GsEXiv9MmnJkRGTKuQ5akHyGni/bXXumFi5zUducd
`protect END_PROTECTED
