`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1X4WMs1twJH+t4Eb3OEB0OAqS05qNgT8EAK5Tt72laoCQ9B6t5qWBLYNt2pn135
x+MSUwGt5YID9wfHS9R99YTI2FRcFT5rpQoAaiKbp35DDyWfbGPTuhi4RH3mCJDs
32NioPYeXyEOgoFb1J+EudERvz9Qv54xC6+vJAJfXzO/5tZ/ekMdiD8qUVud76ou
moUguZWxn7eYwrm3f+v++46bydNa3fn/qX8ukjEGYKUD7ve+KgxoKnqEDgBNumBd
qjUBmbfQQTyCkEW/uGxUNUwBUvySKG5r97mTEYm/oQpoQ373XRI/vIAvV2iitzL0
wg7JcUpWYIGsT37MdMeMRnLWmgw91e4jr1JsXST86V+Yp/bqGSdtnEBS/+1mHEO2
eelJC1/cvTvtL/cCsthcEYRRISKqvCzLqmXmO80UWTAxKmvKYgUevn4OUx/n0aPW
ZRcvMHO2bcA9+5bvKSY0SJK1Z3w+GJfSnDQAPUyoVMriPN9QJS/J/dVLq+T/8QfK
NgmA1RTP95i+qecBEpRmKOCS1pMSXqc8XR3yi+SGBepvN4BPFIC/58gdgPpOgp8A
l5VDFWciABiI3ts/Yexisf0Se/AY9uO9mPXRjYE+ZMcIYBLrNruFAUM96pNjVRCv
eL54i/mThuD4QtdjklEKmADl0P21Wl8DuDd8IV8Yjuwtq1HL8bQOJxAgxVvSIBzF
QIgIpuhpF+uwlGTyCcqN7Net/NmB/XxDiml0u1IyoqKhODfTz7YWknAia7Cykgom
pojQA6rydfPP88NpMUoBFw==
`protect END_PROTECTED
