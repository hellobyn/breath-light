`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2tACE+DQNvxyK1e3GROTMdEfKaUThjfTEzHj2h4DIvDzprSUR18FS2sOuWmkOnKy
R68pisXKlLzam9JkA3yAl9gTXkkYXcaz/XZ1ouXB0YIXi0SbNhg1Je0fTrp0tu7s
Xuz5pXndGplB6GfPY2txjSKZV8Fm1oQnk4irjmmdC2FVP/C1RuozZ6wzl3AVjG/C
VsSU/Eu5liWFD+V5XpkGbKmp2Vu29wX1YMhkUkQ+bAidskl+x81FkXA9qbg4cFJq
xNwJUqCbRnQR0kOXJDY9A3YH45EY7+1aLfRsQW27kzAgW7pVhqa087VgzpBPl2kf
vpoXQ54GEWU31YeItNEJd6rwWWXOW0DbmCXhru0UKtfiQ+ajdDujWWInA2nItEiC
ANqS8l+hzW1CX9XS5ElCwNn7bix27eVcgoWgBc/OVNE2Hnm3Zqa5MRu0YJyslfRf
6vU5KnAPnlKwwOJbvkATWkgFU/6c3k32ycBWiH+LLxA=
`protect END_PROTECTED
