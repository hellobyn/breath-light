`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yw9cn3L8deXFxm88BOHXJZaePgnMBJikfVMYGIjQsITqUJN+suHoxC05VoEKCI7Y
r7M12X7GYxBJgLnKYeyZpwoiR7cVKCOloyXUDSN/JXz49QDS1f24viKpERYInIoA
qWTjLXPGWYjYkxBY3BHwD5mYdsiLtazoW5/nuV7YcGsjWh4MReTskooxX5oyHj21
uhJK5CgKYQBIiCm1u8odpfPU+r+EnXd3e8O8hSWoTAbzxT1baJ0fyiUwvu+ZInfX
Elxxaq5EjjlBYQqjrm30EWiTUoiRuDVdk27+JNS1sLKnhr+CSS2P72W8/XO3SYRQ
sDGMJJENCGlWchUT/JLThWHqqSZDMHfN7zoALrE1vNy4SqsI9QBKPlaLC628dVxi
wulMUqfVhzVmyxpbcXx3dXS+gG49QxsWtXDhDk1+mA60YTQahSmsK8Ker9h5lFBe
fbZfk0PkDfLW6vBjop+MgwcClIo9UASZA8/EQfQiL8BnyPJ0YTRVzivYdWgR9g+L
WMrjamN/tRNC13LfI0z51gCyyQHRegpQhwCCfb3WKWhBSvbsWlCUHai2QyIOrQGD
Wnoukc08e9qbXW0quL4aJKMCRo20AX5YozDdX569DE+NgzITd2c0krYMBaP8SnRc
gRbbSZSvlI79u/bcRLI0hbs0M88ygIlYjsCU7iMDXBSOgiZv7RsWj/6WeUrM/Wmu
bXFucHjlL4Duc6CcEkyl6nl5oX557oO6UBt5XxL6xeJ333ZyQgSNnsxP9aYq37GF
SrDTF9w2cofspKDXEJDBlREoYDVqQ/UFiP8RSruHMWqBWDdtfVWBpkpFGK9diWeA
kibJ7/mZDbj9OXYcLTdETZOW/deTJ6sDvr/0N1XHUXQO8KwaZ6ULJH6iQZBWx3Bz
Ciras4xkdN34nAVMN7FbiAtC3FxpI6HrhBUWSwkjMD6uNffIzck6xzHXuexpeNEV
J51STTsUB+iRfVYuQ+oUZ9vzAtLtd+2hrAQ9e4EtOc5/1c+f8eaYCYuRYzqUe2dH
+d75pn2/G5IEmqcU2sWvG6A2/snB5Ip1XfehfkkMdOkZviO4R7spQtwa0/raxxY+
7d1nkQQnoaBso1Un8RLNReQgdZlhYsAYM0opZkZa1pZ6YBS+kO/stBSs7NShO7yW
OU9kYQhjZHhhbVxWKMOyN7+cfOlpSdKowkxgdcVhoJtbiXJSu9UyqfHnvA9gFcTB
ZRmzH8uDpuK7l+MQuLcPkBmWFF9NhXx5X9A4WHXNJ0E2aCsSb0fABANxY3JbGyH8
BBYSO9aftO4HNinD4+tAT+V2oiSrGNQzWUSvcZp9NcZobNNRIWfEkhZzxi63cM3/
iopjoUm3mPzJNV+ymQccjBHlI0XVV6v/3K/Sb21eveAGi3DYTDQqcYL4LnrG2NUM
jFxHFyaKA3dZ2qXWoBX9R5PyqkoZzVbp3r8E0V22WRVfSjMg7ki84IQWCIYiuhK6
fFBH4D4XRi3FzGf8Ehr2bHb0w5MGhTzVHeyjKRwcIR4KamPVVVmnG4Rapc/Yuyyt
M7frpziue2w57/BsFBHD+F21OZTNKiDu7sZxJOq/tj0C3WXiVOnMmztAOiAmo3KJ
PHt9veEiQnnf4MsI8nUS+EqOa+tSfE3zOTigrDmB+JLGcWaeQzaP0m4WEZwFxVXL
nB1YSXG8R/LjJZD2TipKoZgGyhtdqnx2x91u72VnRL6IWkuiPB+NnLcRMl0R3o/p
R+4pWD9rMcdYCYW4iAPirh0HimHyMk4WwYL62F4q5FOVHwo9LliHA50fKFG846ZH
DPzVtjkRriGBhtYrrOcJmjc0wC8RTEbVab1XckQawzNn9Z7qsDtt7/uJv6JC/x3Q
MaCLoBfnlCNDgdBie+PdBy7yZ36yNxMlwh8jPgMGjKnKfeoBbyIkkdgJhM0gkkoM
3WGLP2FE9bLXvITIU75nQkhkESUp3re6nn0R0P4PeXYM/busIU3UopOovPxerEJZ
rXcq/9Nnh+cA417T2KKgROfqhTwP1u1qfatpaZgkhYqXbfdCQbh05ZfDPlaOCTsR
MtJ/LSnMyICK4bZZVWjdoY2uMzVfOp+es+gYG3Ikq73vVy5+630CEFVtBxVJexG5
gcTHUEPOnhTAEzd4KX54Gg2DWKqLqA3fKutcrwjCFaiQINFigg+2AsL+AYuGnAwy
U993rH9jjpXBaGMznwzJCAB8XM9DI2Aw9yeCpzFzvdMwk7Gu5giiZK52MXEz0Uo1
5ST3k9LrHejWohkVVYjl8Qe/lw3n6ymC8okR7ZZMutjq4GbAEJRkc9LvADYMqegk
rUma+lfB+JAH7c3WpWmryieM5noYDwUqJu2n4qXMKeDmvjti5qPnV4CzxJtV6iX5
+bUdhc8k0UxPUbGLfJcy7DputUnnzy/A18mzggp3lVINHFhOHKB15Tr9QWRi/RYL
ZCghrL9cdNKF23MplIVmiUdDZk04VHoEp2iAgoBJwRZQp0ktdjfsGkGSBH6aYsel
GIEIciyuR+e+ti2Rfc7tbtfmm/kaT9KLb6wQkIJmOxYsoZuXOGojeUtxlzQwW3ft
R69ezwipOqc7wVQRQxwWdtbh6deIrKcDBxtbZlAVwYFH33bEz+TNZl9nGAj2UJqn
xvtl16GQP8j3b173/BoL2sPPeP0I9K6e33PF/J/zTLhVBEFHcy8p6t1VPzH3T2CK
UstuxC2X4BMG48rDk7NWFfMfe6jj9aNtaFgQ9AEjVyhjDp6kXxngzyhszlqRAJX5
mjCZ/ADzPVUEe2kDyyog7lCCI/eNc+tPMUPgyHacd6tbg+Ja8HdmpK86LG4mO9lI
`protect END_PROTECTED
