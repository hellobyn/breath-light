`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ue8Qs+DV/5caCLYkC2azycuioolROkDiSwgU10yHTWkzdQ6ORosvCIB2PUJjAf8R
WAC/UUhoVaVddk9LABpCT8Y0ObNM5FsTukeeKU2gL7bq/ISJ1EEI+dGbZw40OYBI
5gZwjSZE4Ubt6LKqA5IX7sfSrQi1Zuw2Rt3YKRV7XKWim/lPlbDEXGHpy3rwB9VC
j24Vgmey4O3F5zQsu0ENCkFUgh2tzCtXHB7xJFhYh98CVymUa02MAwnTiKlGAlik
8av+5hekR+CKOq/tR5mhU9MJ3BDFH5Vo6yGqmMuyYw0CKBCW1pdX2auOQs+ImYQa
0Qa2Gqh9lu8RB21KNjKsgAajYIdEgojJonlQRvCpd5afQPgZ3RLBba8HVD/s+cJm
+HGg5Zseh3Cu9ioxkO8PQk3ffhbSFfuaZH/vbThkcZVG3waLJCJKwdboaop2r2Ji
/dz+//sX4C+UvE1BvJ5enCqmSMoDZxWhbxIKy1d3pOIKDe16RMdfh2Mf/h4xVAmm
KmTzcS/9bP/F9xgN/oMdaA1xI7omy40RzZSALV2rdA883Ou9MJdTcfjd3VA4T1JA
IxOY0Z9kOlhXYid19CUOCGNulGCvmVtdK5AuwNPSUZplQ82sMCzzn3QVfOkt3wFb
FijVu7jmwBQVke7ZaPOGv3XA9XozqxXcLlxT5+tt7Tg13EXyD2nBpeQrFuRM01DW
07L0VZVDdXnpuReaewpBLZ/W2H29eDffcDUUqZRoCrn+134aJW3DKWLDzxBDe6Zy
lPQ2RRG5Gymr1qtPCRWqaINjE7YNSQYsmmVrDSIu5QR8/oM9eeWt4mp4KFAyk2rx
`protect END_PROTECTED
