`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prrxQhx+YbV2V5wXzr4pyrHgzjqaHO+kg7beLsAIr6ZrH78iGCLnB6zkvdBp+s9d
jGQexmpKiZPOurj9sAuBzKx0uNEmXKil+XiokqeNFRVGZqpgG1EWYFboqwNQ0J2q
f7wQmRb70Nod++q5hsk1f/l3lbuZdonYwqKHd9YMboJUwnOlvV9s13c85b/9Htfi
e4svBlbGFyhQcFIEpXBbC2jx5MjwRSHzVdqlaz7vL+PNkGI+GI8lSEoGmKm0HWil
t2QEJE0oiP5vB5MEiwC9OV7QDKn/eh3uIXIi1oxm52NZlI4yeVFPcbqFHp5UAido
UiHKEwwymisyZzRwRODTRCtaYYPuDGfFxFM/guxKP0yfIGjXQR/7rrAWhFYe3hua
dCsN//9qdtZ/dp5CMcvV+m6WBmOcwFduezKXHDB/wai7SzCHkP8Z/RidVt/uQZ46
x/1wjUcNq461gFEnoITiJW8LFJRvIoxRbkVPGgvlTlLe0vUnOpepCE0y053gjtfN
zUpXh8wf8HdcBhMyrgWLnHPDXPGr3NwcOkZ3hVJgCLg=
`protect END_PROTECTED
