`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SfMWOx+bTPTjZ2X7QNoTXqwrDRvaqFP0yUuOpxAu94bDGnS8ae6tKLj57o8pORzK
c4TLXrTXYXUHPaErjMK2a0Lf2LvPMopapk9Wal78uZWMi1+bmL50Yyz+X8/pf8WX
e/2tsIy+Cy+v+1dImhYuA2Wsy9790BDRi6SE9z/1wB4enDy4vtIf7o9P/c9U5t5M
m4zbKDg+AeIVIeo6tdDj6waJln4cYqyn/Z3cEWog7khtuDyctvmZZVV/e03G45yB
9VcmU7wpWkeAz3ILUDlBnbwCE05M7VCw0yDi5cISfyo05+L2s5Xf7chHtVQM0OUO
yjyYmBZ3qShSAN2OPBMxQuFjZHikhkyzJ+hfcko1k9SEwuJpDnsJLWg6MFP5dIjH
gL4IOEULNyc5pOQscQhNIi5IRpe7pja5k8Q7ZeH23vbs1BeaTcyhJfFZg/r3diTu
AAyCEFPUdmYVinjoe1mudjpzIh+Zlj34WF1ktkT3V+eRVXOZqZuHc/H4foBU/6lR
UT1WZbNzPZgO73j5a/QhgQzey29GdeADkcRXgqiG1YxF0+n6qYu8m4Lw4p9LJkc8
SvtaDSiIWozDCG6UedbQ/okIFef9t52MaNcQnnavavLMTjhNdEloVhsU+jtQ9LET
DxEZDBSPm40fJT/vjkAsA1/zv3VXWG99BcLlpRGmSgmD/SNFssQncsSXn5xbxgn8
r7KdnWqy8QAooQl39PxhsWLCm8DFhR0WKrTAE33GAFV0z+beXYjb2+z3RKjfFIk4
PHvt2oTNQIgyfcjejwwOVBO98hSGAn724mD1jTFUJEC3gq4aQ4gW2iYiKKVim252
1NBnaEc1CIDtQv89VtMfghuOAolEj+XHyRIDOJCoNiwSLO+uDf2B6rA9PFxzWOF2
eUpHoQjTZuH9SaZtDTkAMDF0Hi5EHsqRY5yRXCcj6jqAPMSzzss68Nl7B7rX7WkD
WT3LJ8QAR/hVAuvRHmagiBHCzfy1dns2BTIMg5QWqDqYueD4iIEm84hrvHPvYChR
nu6IaKJdO+wQzm1sQrIpwGAO8xhQUANQFtCVn2FA4PiOx/lgPeZfpnX8fALvgcir
FcZ8+WNUsm3YGNFCF9Bw/5YzHmv1INbXuSfsRAKmkdxh21xbRFqolqbeIRv3ctQh
s5p5Z3E7KKCkLUhEzpxUK4EJkKSzsNozF8cQJ9rVuW80htWH2+4DB6jBAzHr2hNM
sKwBDDVRgZKMXitbjpC/VSDl1gQHEWjkgi0eOpNc54XtZuorAPWV0o8PMD6mGdhN
RNS7g6olMR7KT+dC7dtA2zakFfdZXuAFQ+OBmgCi+c8Ad+zJ1VKx6cs0BNirTSdA
6vlBVZ73hrpajKtgBM3E5xUA14Mt1wn3SuEY7rMZ6QqajxANEKddeQxfuzrsU094
LVNGIDz64k1NDOlowi/YisHQkFMjZfEB73pm0h+/TdfPQWzZfht1xVZoiRxZBcSE
mjJpNH/n+ohthqpEz8FwPA==
`protect END_PROTECTED
