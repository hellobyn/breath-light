`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yr+RxPdQmKQCQv0wcLFOE/3yvVbr0fdA9x+D3x8P/aCBiJdXkJ3YmEEWsG4Zslk
6ftqrOUDamRgVZL0qGidiIpVrdOGG+T2NjGzaCOr0ERtuEFZYOIjVMB6thzpB1aK
kiqHt+ZD7r0r46wOUo45lvBRuhEdnVQ8Ttbs60TOqo2bJ1cSxGBSBKjxxzVqmUsz
k0R6YPPEcUOhoXCF78pzozqY/HZ64i8F/v1gthCFoMdpHTo5wukOFw9TW53ZbZQB
U+AdjACWZcc/nAKOwGzHw+VOI8+aJYVd99cq7PGahgcNO1Fk4D5atje3SKgiku0m
ugpltq+CKK4diFYPAEmI7WEpNhFsg/KtgAaSyt2UyufzqvLfBIQvlwTTvF1m2eCN
5UnaN3zNtk20Zzl28KQirD3uoLFnqEK4RhvMmhdvCmigp7IAGQZqz/gqmKfdO4r3
B9oD6I02/zCgvkCK6RmIbyupKSEde37ksSSWl7mEhNZDkzkPiEMPdEo78xdMmrJ/
Me67hpQ2PWzm53wWBhEuJJsLfFOD705P+Jb0I+Ar7wksNaKHL0bgwcWJdRnwlPha
DG2ihz1cfJte7JCD9YVZqtGQMVf99iEoqTlZJo1XYYgBkr7UOEIqTpz5x1kjMoL0
XFBjncvmYRpb/GKIUBWztqvGv2bvfO97iEyfD4RN/pu/zFK0FLY7VhhLnAAZBzik
ITy3O2tsPxjQB96Ii3aJpXragvwpBfNY2wvaY/AugT+ukqEeDdUAVoMmRsv4DdnI
8bQDnpgDer8cJPdvy/CrAkLzrZiDeA99AhR44PPgLfd5ida4MAuO2adSg1pPE0/f
6UVCX72t0PtCsHxvFpEDsn1pVE2nArajvn6myT7ERJkUYq4C2SvXpJ7qIEI97EPf
X3bmakRv2ZgAKrDnHlz6d6x3iwfF+YW2CvGpSUr9BUw=
`protect END_PROTECTED
