`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2meBAq/f5ODPd/1kqtxZMzk+nNW/7JIFXYZh+WjhoDwMGrovUFiR2LpGOI3D/P2m
nF1MwX+NWR0XqJlZCer+Ff1oaul05k4idPU7XiZ+StBgTtoarbK7tU9T0NzKtcD9
QSsyzdY5vzZt368bjIQtl9/huydOvMfvO0SO5TS6rGzj/K3I5SfisPuFJuLXoIsy
dZLDQRvg9WcUlCf2pbKzFd6YN/5OtDyHPNHRutJPHnjPrENMFSM/dyvhagVwLnE4
W4mE1FEWzFdXMgWBgUljljre5UCW3+WFjY3qHzXwSLahqrlrONfEg83Y6wz5LP3J
cMq29xzFwimtvrHY5CcLJ9hujF+bfbBoLCgHEnbOpOUyFR1i51Shf9m3PQDE2RPK
JoUqkVU+kcQbhyNZzTglWA==
`protect END_PROTECTED
