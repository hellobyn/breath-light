`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
InA6IhN6b+KvMpIYob34zzgjPbC7QAZjqiBxHrBsBOcjERwCzpUNMqwiJzHgfBFl
5iI79gi+7lugonxe+UwtUVQy06/43ezXC6KhJYhcslZS701cJQOPUNoHaqhYCkCH
U+5IxzLzdkcRRSTGPYXerdxuzZNrboQ0lz81WVM4mPR0dXUGNEx5R6XQXv2LOMA1
SuBlZuQ49thS9rSIz5t26hqbiIcIQItGWnjPrwpqQv7HRTHKirwUaS9fT4v8TcMS
0C9nVOcDwImvRseJ/F9OnQLIp9+hb38ErUJu04YCVP4/zaU9Z6HrCdtzYYBUcIhu
j76YoRCzTiHacS4XFK2PRUrdHcxfbQGUSqjVQBAXVKpQ2vUWLGpds9WXNm/Hph8l
l5FF8n/mF8+XQMQJF5eXWJcGiXbZIopLLggJHPmt9hBdgz1U7u+h+rhDRjEhRL9K
ivjRb914V3baX/9RDIddgjH67u1xEWe9HMrnrxQKNApOi3+OdbjG91VpGePdiikj
ocMI/2yKRIKk+wZf+TpeR0Dhsw7qlceJHGJ4HK0ElC9vIE8N7gITuoielJ/C/tAH
LZnDcyXeSKet6EvQb2K7+dOHs2NnB+GSdQ7ALDEYub0bN0SuqpbEO00YuB2cbbvP
23OF0qHPuKkmQ67bFVYPJTlLc07Yb7Ivmv6Mo6xdgYzRctUlvoRmMpCGj+RU3k2V
yD8RsrEtPQCwPbTh2vLP+XqFCQsatYiKBnfan77CR0dMGlOCqZsd8vYIw04WKPEF
x+IuoBm+it/K8TdE35Ki/xxhzsRBJ75LV5OBSXEHoGfcnMdW/lxtAzGPiAloB9N5
`protect END_PROTECTED
