`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6H9FqPJuH5Fn6Oi0rHQj3LgEOspay+pS1ulLMxbDR+AyUIFfKomKkwNdyM7CPIO
VfNNm7aXwNOgdlFQZct/r9ZhhuB1qd5bHEdm2DDKwOUrB2/T57UfiS4SsJRDjTVg
YFioTpMROiuoDm7HPbWXdCa3h3j/mF37+uos/zV1PBUjLemYDmbz5LRtR2kgNrT0
HysrC7qd4m0Zaxkij2APg9aBowEfaFdHG2cIR137nAxXuOAgzBj48uQnry/2NCsL
2yiPc4bMmOLZvOfMEHZ/RyX8UciFCGnA9nbnxID0Wa6FG39DUPOr9BJ9PdBz/qnu
6g0K1z5Zi4CRqjgiH/XijzbC0RZ+lh4hatimOZCiwQc2ZRWbsxDyzCXvIGhZuBVC
B8mHDfl8XPuNmYmwPbAqhwYUFrjkb/WbNXZfyXSx1tGUFdPanEm3mMBVH7Rs+WnA
9MuUPf/e1mm5Mt9ktApmTwZj9em9+bdNrli7Fvu5Ht/7iLit5yFjTG+mcXnJ9bvr
FZHXEXn7tKsOk2L/J6Mnt8RHSzoMGWrFQW+La+UnbrJtRC5uEJ4XVCwCzapJT+cH
QJ9Z62I/zURbboQxNtXa4UKNlNHe8UHLmFRgex8zwpuoowAZxT4eU1vbsYLSbqIi
1KU1XE7XuAh9RazNRlPDDHsF1H2whG0YQ2NHvbqOf8g015qcQQbTBNnsKNpKD6Uo
3AD54J9cQQvbYM3xDCPj23iZjiy6LXZYQO5baYK+Ge0WVp2E9dVKtYNCqgv8dpEw
5pJcmHIKt9hHLvNp6h49Pc53/ZCmIKPnNrBsnd+aDkcxU0JpJPorhabtOl3o+5+b
xZKxtqBaoSA1GgwP2byelS/Hec0tx6Abx2fHvLTYetHBwMGC6odvpsPGUqeRNOWA
adlZ0XXooC1fuxQ5TuEH89ik+Q6Q26tuVQl3g5rRJ13AJaod4Mi3t+87xUsF3Z1Q
JQIjHFF9AQDg5a2MLT7e6T7b0MagCt9WeqGQZ0sEkBBJlCfw6JbrejqKNhbEdkJQ
gxIgKQvh/i6mWyl1BQAYMcbN7eLS/vjo8mvBaggnO1mShMVptMvr1rJk8TEMyZSD
NKk/3ENnPPjsTnP2r9yeX537WLKSME8+cmPGHoK/iUfnfUV8SwXCDfp4QWfWm1UT
RMILUVyA84jHl9IHdkqYaVwsOhAkVvI1PBU9LVufSj+ofzmMNVpafwfo5goPrwXR
H0pyZQmLEgV2+NwqNaxrnCMK3DI66HoCeVoWRwIF/nxf983x5yIJp7yv8/dOO35U
3DSrQ2yawJGDq9Zc3CSF+UUaK1kVZaFcqKucf351kn3fwVCf3S2wG3G7BVbprjfj
SewwmsJkEYqqRNwWCMXjWk5ahugPSYIMzg3WzF/7BiSMbGoOvBodNc2CP59FPf1u
ZbGRPm30ztG7uWBQhZ4CZEax6EZ2+qnkHHE8+TJaT+AAA0I63omS1nXnTs8/6IDB
Jrnx7Xp6ZTpDdz1QuJKZ1JGnBUT9b+QipUGjhuiXOtXQedxhUIbWxxB+2y9/YWqG
u5IGJfirJFdQH3l+0ViOSxlRKLqkKZ9MhGelhyuG/FjAbj2+jl4IV37hyuGH06kW
bCyOZ91HWVtEl39UrvKz63ybZvi81YR1mU/8592skAYINOa66LrIr8ZQkcH4KAyy
Tsy85Q999haItVOrVURm1KTz0b+/sKIRubf3H2eTzEmRuUnsdulC4nMnlISVrme5
Byz3ev6TrZSAdgwqA9oixqCyNMYf58zg11sCyVni5/uAwTOAAZxk00XqtDeiD+JT
mBna7OwexmznzMgcqMrS/LYH3Qwrc7kjyQi76QJwwFoww0KWYQKKU2YE68XcKnwL
kThocL+Ox2bkSkr237WRxVifvg+evZpSDKB7Bqb3umqUG0xQwkX/bivJgiw+zjsD
l5vv8hQ9JvRj+dhZ8kmKbPfVI8SacMCc9KzkxFLZC7gTHR/YPqWGcJDjxRv3JtUH
reR89AOHtoak8xvpFczC+qbJy9oLoBxQfD9hgAcY2qWey706lo35/X+ZMSaCdbS0
fbUHfloPMt9etZXHfX77w6llYlOXX3YCo5kgTEsd70hRYMUAshGo6EMsXTFPDRRV
ul8Mj5HNyKEaFa90DiM5RLLulR2FItNCT6kK6p2T9ZOiDSN6GROPVjwFfiuj7HnG
QmE7O3sSp5vtv85hFTT7kPYUai/+LqBIgnoYd8tnfEQ8OtbRgNwt6um5jZH6FBcz
qKZNZlbIg/8W9F0i/kuQytJVnS/b3SKW4m8FSjyQhz0XP/BVQkXBGRn/pAruaOxI
jP5BN4scqZxhaJpNZS1sdmbT4HYyH8PLOWJDqoaX9j4BfSZVCoa8dWUN5ZzsoB5N
uVW3PyE8VjqM7Xt00XJkbh4ksXnL5LgG4E58qGNpwoSDSmETIXcmOeI6gLReecl2
sadRhALV/KOHc+u1te81Ie491KzcJHu+5k0R07fhNIBjw00/DYhnT23WFF2OUWPT
U7iaFW10JLVpBwAFNRS5Ice/vOBkVOT4CHPSEChLL3X0MlSp+90fRW1BV4Yu0x6H
ir1ecdOOXxuTuBDYbjghSoYrE4pnbG+ES9rlHNX1r0tsFKusBmkKsXtGpfDX1lIG
WUv3nRHf1uQjA+xQ5LUOW0XTeqJbs6RjDQ2LYgEzI0pYJFN2y/yeeeGhUYimA8fl
gflOvpgNamjemae4tLEAzxn3+jTyqPv0H//33pj/dOHrlTTMtqIZsakfsO0ijjwQ
ICo8vip2I37Xmp9bB5bj5Ht4oGT4/xkQa0U3yjBeGXfjRDBsEmQt2hJxpllHllgi
R9pE0c0v++Cf57djXj6Iz7Dcg/1d6yeEP5K20JpiG9csrHdp7yZmfwD0/8ZpzuTG
KXjTKkGEMnDqyI48FjVHLhQvGv02qL1ePF7lXEjmzrLjVt7tGr0iaQxftLdwc4of
SnQRLQluL3xvs8NAFOXP6GeVUqOFKWwAMtkSO2mpZJCzJPDpgK0+7CGr0OGPYuc+
V5PNi8iJuFktOeYm8Zm4YTsVp3V/AB+FatLe/UTMA0u6K3bVCmGdQKKHHPNToLOs
I7Uxa9xXQrpBNZjmulP7cDtrf01b+mUyoWT0KmC6OrIfCgXDXsQeR2ZX74vksKjU
anZXtuYeBdgUwyYVLiwmfkyJtxki7+6FbQaUgF13nnn6R5sYpLskDZsqrz1SsGRZ
Jj7vNUsSWq6UIyZmwd0TFvKbrbvQzl6sMtEY3kw9uK5CXuiST72pKdJ7tMGU5Pag
9ohxEGFf6vB7/O511/aT0p+pL6KfUXpW6Qm+38KQTSkv284Ba04gSOqRmioOduc+
/EK43j8HjanPn2IlbFeSq5KFrA9SZr0nUCOxF6LTLqHnZ4m3HuXqZ0Gym/FrH7xG
o0Gm0bc5WzLAd1Qu5mwAvMFGpr/hbXrfHCzJ+JiMYJ2pwFQhpNUarxb6m/+tluzH
`protect END_PROTECTED
