`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpEskWHCGOCGSMYzYWIIi4nRtNXB13d4e316guLkEfIXUAP6s34kU5iAk/PBMcyu
9davQG02yBvmIHR6uCc54KxJL+g0L0NQAF9FZYdHQkGTsWJvsabfAH3WWxve7c7l
JcrL7PAPB0ZMB/99TBzi4CdD6/YqxHHnrh5tvJslpGr16ijfp3s4omYyxoM1uOfT
Dt7vHGh9i+oOyIxVe4jzPUevlFgb8Jt6Ptt6Axcl0RYZ8IPFucOMAbYTeaMYp6wS
oaR7k07q2X2PM2V45IbcCvR1bgVyA2nnyU/f0xqHKoQlJT0Fz6qsfa4iDb3+ypiw
Ly/fMAy565vWdMaiazbJjVJjPFXBuL0CpEG45fI+0Xo3Zp0dIAvkGwNLQMe5+nRN
qoS0pRgDl04gqiDXgy/MiyVSVNZCv4+f1/Hl5W8CsOjmF+QnRj1Rhyyk9THwoO+/
35I+ZsQSOX/tDpNFAKwYgmCTv2rSzkONnrg3zZwwG+4O7rAqSamTZjNlOKwuvAY/
/9f9pIdkKLuo3Azmgt92euVbOyJ/c/PEpo2PqDWRohGjBwKV5O98rvUo/+bVbPz0
3eAqbowzp9yNwRIBKz8ln/ayCQULRFQmlJNtC1nXvrswqiWus+C3X6PcJK6f4vYw
wNh1YRV7jWvJlMJUzVOw1TQa+XAhKmE/T3NcEpklSZh2MTSijtWF3A2Sec1Ax1uw
XUnKLqRE9RB6HJ4aEWisdL3um9aWumeVEiADxJ67U6nwmsJpxonZ7g5uu035dJkn
Ba741TVzqcI0TUup2r6b9lb0qiArfptVD0eSHhxzoPclFER+dwX8oLDJHmkltD2w
+hYY/NVZh+g4v0EhZvHirT8Y6yDmJ8LkWSkYG1nvM/+eVCjXJ7FoS96N6vsMMobY
3uDgib34UXt87QQhM6X2npqOFSsHvVo2yZEnG+mWJUjM14TA55TCDLjVi24V363Q
cOfiM9HOyvj8Ws4bQjGu5PbW537OHOyekqm2/mqVC+JIeYt67rx7j4pgo1kOGQZ0
RYL708AO88r352f/9VClDKNL60B8Ub9CySym2+K106Bhuv8vFhDTHYFgr1cJBFPt
KUWpvfBOrpoU6tBsAbE3Km9V5xeQxqnVIhAxaBqi5pGKW7/3kLKeql0o3bgK6h3D
c8+74y2Ze6SO2j3Xkadzy4X2bVDmO7D8yYXTtOeqENovA2+LV+1b4YhG4tn7TKIr
YsbFmbRi003Kk9yqA3e9NxPOCo0rICbubPebLT0KcDz+r5zaOkR7hvVUZzcnGvJE
vGWkqBdLmpyRtWrUBWtvStbQd1OfndpwYf+I1un80IY7qZlxyD7BZOcX5EI2v804
H8dTW/Aw5ctsztSMmAqu4XhiGAEZiYgVWc4gyvlfzJLi8UyJtjKZJvi/6GjjM4Wb
L3nARQ1dUqtRa1CxrvSALHFzah9ECV71+NBi21mXoIYInfV+zJpQv5yMYjc58Kh2
YklSS+UGdy+yndIq3Ys7nXbvNmEpfnST/QB3yAd9LY4Ca1L1uW3fTQcNyEc35+fI
XP7SMjeD3Lxfds/SBBaQDWVpna6rNssYtiYyWuGhuuQsRvY2Q/v3hdxgGjgZsz4N
v2/TVWM6IdhxSrsKwSAc5Lum16eGHHNnqxvLNrdDOCjkk+NCdMNa8foG4NtLvJ/b
EYKUNamgXJgKX5dCfgFS3XJs2gUP5gUeCCfC0xL3nR5KDo1N10foWCE7MLb/Dma5
80r807gv9NuqxkZ30nNYOfV6F0ml7Tuyrf7GRX6f4mDl02+o7Kk3W4IyLEaNiEFf
XoBZEfn/uBr37yeGmbs8srYMdhot1q7SjldFk44R/FihDrlCuqBEWu2F/OFhCb51
yARgnbb160ZxcEtNWGyfHCdkZ1f2ptk37htd1G9UYlWd0eIQ/C4LcplTT23q7DWj
QRl5/NlEIcBsLvhRq2zLnoQROfbW5JtbiF+UpuHPChcazyfUSrBTp/1wxLYwXZGN
d9KbuhSoRSPpxLgEY44cNXRgIgvjEdjsLXONXmpLukYuhq3lVH5coRjGnyxNt1Ea
gRTanyyM5TXeocAf5sTwE5l+1odlpyMvtAcMBvaJeZas50oRcPJQy7meV6VZM8U+
yxTTTx6wfj0dKF8dQMM14rs/tJCOtCvpA6quBd67XupkkqeLDmNlteS7FA9tzQt6
vOnC88SXxyWH2nW36QlpOZm3Yvi85a12M+vi59J7YtrqgU5Rbn0stBL/sRMp/C1L
1ToYLvmmO+15ImRFkWGzKiw2ZRQS/zT9G4jQN1gTX6IFbEuHBc8CWOKAaVFwakSk
DD+5QoI4fCkAzCZ3JHBq0vSm+hffoHZN7P+Md9qFxDu89e9I49FL6nYSRBxyeQzi
A9x6vTktNqJU9fpgJDPIx//tK7nYkyCEYMOZCOvhpjZ528hGTXT30WUptYfLioSV
maXZ9hN24PVJpQWBLT/tsWqB/nwTtFrqy6ayvsoDE8/OBHGsZ/CajNi0hjzsjIkv
HnRCuH3gEoT75MsBKm8FGiIT3qe6OrXaZHZV8ZT5M/hAJ8LlsuHkZVBg6qj5f3Tp
65lCPWHh6+TmJ1jP8ckRhidnsr3UTdCxMtuv1uKOWnyFbHjJEIbFxfF3TNMzvYkr
ag19sHyK/XwUqPNDtTCt1wf/BJoc7WWr8JfTUC2Co134DSXVUaspgLD8eZkzFpjF
Cm6FH4eCY3HVMHAhjGJXIMLuZJ8kfi+9D6frKvkuIHCF5vCVjRrJvMn5qcPFwG9u
paZdW5NzjnDBAFrZsq/iOHMApIYEfq6F6hwcULetpSoZThM2c8iKgTW69C9CkOqo
SnssikebNB2Utrd/0wy+v1h4qUtMt2gAfclCZaVSlYa80LzSKfkpzZ3xN8fnq9Bd
2aFIi7mp4j2U0eXFGIfUx564KueO2TTlQXU+Ag0Hz6APd4iON8DGHmo93rTACqCS
6xnzuE7i2paQKg8Kr1AdnRJZ1dEyTq2pnfoMB6FQw5nhv4gmlgliHcd4yST4d+gS
M+0c/nsC6VRMFPtktebMLyV2mo5EjcFUdjsaI8IdOicEVJPzfXUdbKMDTANKQky4
cvJ7eLJ4/hXKnTw6qp6dpadd//KOTb5DphtULVVZC7Nh5iH86OFAjbot8X2ino65
XZ4i1hEKvJ1JRnBWNcNLUoOEEoZzTtm3Ph1vJJ/2dZ0l92xi+nj32zidY86ufHSd
pF9TvvkgtJfI0hQmXDdpfztThTYVvEgPXIQzdZYGm16T7u251qQdp5OlMyZueu7v
mhFha5BGbOOMtnjpT1fj9Q7kgchAdmU4xEGziCvJ+UMUbzR/yBQG6fNikW1XwRHl
0JdMTKdbCIrShE1ktIT5yFwQ4kEsJOVswL9Zol1Z6muxxy2wf5xDLmf9AvH5z15/
dOVpEb+1IEVqfDmEiTQ88GFvdJfKT1kfktHyRVht68c92EYtroCO0zb/b1BzsEii
E7XvnDnHGQQZkX1/0CTTWT3wo8jzbgTaUitAMlHajcsez7Tca6RCoaUBP32Pgcn6
7eWS/Lckx6mfsiUIGoluWOcNXyA5tCHV4JB5UvCnRVv6TvV91jdoQtZaAdP6ZIRn
L1Uy8Y/YVn+BTQ/JwnZffzBRjAwuNjL19ujpYdw/w3msykzbwzcRxgMCv70hz5m3
sEvOLLppb5i+I6Lp3fUzorZvJjRm/MzYeW4O2tg/74Z1ErtLqtI1ti2Uzjk9pX/R
370sYMess2edimKc2JIjyXFQMM+IBGwtLM1NgKFyGJ7hlXvpZz7qho5JPE/lG+2v
5+iXrFtlI2c5R0kldS0sc/A+RCKnzP8G/1LsaQSSE8S/VCf9mZB6siGsyseLyOir
87H03xNe18Kq3/t9ccb62MZyaEwPr4awaOK0Ec17a4oQm+l7/475jrNGRiB3LLZI
hct2/UOAQXmFvglT6v3I7UA8yVT7S48EWAhVX/DE0CLxOg1AI7kbpbIdCXCARZ8t
LeX0vmFabz7vtGTD2OkbYbj7USn2l8kM7KMdEzoZbetB4A1z6kwaIa214RiGbECc
rMSsOMkJFm14d8w0HSd+5yxx9TQUk63GMEd+6WQ38OpFQCxuZJBiCKSE+JQPgNqh
r+fA8bamTp7pcM5dxnNojgYHCXTE/2qIeaiQs4VEM/ka8MQ6g5P1sezVVyNgpLzv
WiXE9Dx7gIkdR3RuJ+uJ/KnXpLVKfOnDV8Q45ZTLhTQdbCjDNPIdqiRW1CsY4uox
elCKA98S0xtsfxjbsa9h539cSCiEi3DiUveUFvt2khX3LOKsy3Sgq0qMz4gBhHhw
flB13HcgeBFhduMBa6V5oG8VwcIWgfZRGMhO+V8v7P+PK9V5LSh4U6PBheGNKYRq
yGO0t8jaDX8E8+aJUdtJovBF7N+Jli1C6Je8Y02rKA3W6dWT4x6KlyESylKvhYNE
XF30uSq7mBygjVK2vn9GeNacYhZRU6yRZbKpxQ8cnTv7ihBXP1VJxMN1TK7iu+hJ
l1rZ92TomejtnwPHZT8qAklGp1q7bp/Pq+2qNRuk0Gqlf7S5W1/bm4WWgYAvUnri
d9767XaznABzSw5lhsxSt4HJrnp/VGfhvZE86+ikXqeLJNN84KMSvHqaIHvd+rw/
OkMl1nd60jJChSlkivA2ktHUOMaNfcNQzpMcGmajPQ8l48+67NAkU/GD8pv0hUmO
Nk0a9T+PS8UGI2dMPUdcAvkfhWk5O6RNcz1ju77FDtWXJLITVMIHaYVOOpO5ISQf
ou24Pc68tpnT7ZbBtG8kKpftspayjNJdpIxjgD6jliDsPxTAAA0PDwucG6fM0+r0
51CY1p6Jv+fk/5Jqzg3Shhg/+RIlI7D9WsWSVKUflEEYzmRw0s3HvSfwVGYj0g4n
J1RbRBzYpaoQrQPp7veHd6I629E9m2rgYPzwyVTw2pnqYZ66Ifu/U7o+hanruXKD
hpaSZ0bq/Eti8RBxmjl+wOFn9L7KInoEOD40lH6fFojMQriFjxMVwqY9hM0IB+TA
dEMCCHU7XpNtUfZGWSJ08+QzX96i6SrifSUCo5oxmtfJi15aCqxwdbyr1oa1798/
jqIDBTR18+mr4Tprm76bkxacyJDhSFr9cRnM+covTd7ImmIwE7pXqGmhzhrknpMc
4d10Re+wKKzOq08dmsTopYQgfnxHSKkiICCx1VuLVysNEIchK+Ya35thcX9afKAl
sDI+RmiDipQ0x9UxPrG7EtWpuWsMxcAeEaAgLjMsxflnUg4uyiXWdsd07vF7azri
rYf3Y1xKfgfWZQmu8GU06MK+1C/rqgKEbWoMZrRCRKprSQFr3h+m7eaqoWiH4weS
EXTKZclYCFHzde8pM5O7EaDBJsnBVUeGLrgC5VzD6Y50aYj1uZjQqvCa6EO6rMf1
cQwM6E1JlGsaC1IWx8yb0wcS34nGcOjI8AYLscfa0NwFiRBxylizEBEAJt1wzn6/
VL0aqdi1RWbzZLmrPHqWWexFz5KC/tb4HtxMDC2kFhrD7Dxr3MY1hG/5umfTzujo
HEDhVhDhUIRQVQBkD3jegOzT3lHuRNpgqQKmUc1GvyzQmVqCIfhxPr6AwlpxOLxV
krsPgDECN5H1g7B6FsXJVE7enwWSsKyRzexx/Xd1BoI8/YUjqeN4S6JNSL5zsvg0
4JyKhxq655adO6BDFoNvLUjBtrp12p/F8sODKuPclHEl28fDgFzwb6NcQVI53Q7B
fprf6zc1DDk4cum+6K7h7Dgmhc6RYLbCcFp9Q8UwZs4q2JeN8/jnTR+B4FyRIETY
WoOGjQY8EKBKzmAb+TJ4lWM/Np8hBs5ZfKoxT39k9yYu93gF/Z/ZyyWqQBVgeSCN
ucaJUixEXo02xOIZTExnTZ3Bna2wLufBmO0+BqjKBX+/wjT2cvQz7+rsWk63kwbH
7XTrib8wnriyKE7uincUeTlXe6pBu9crhueAK36otOfJvNSTf37vGTkCWL47nGFU
TPMU8k/zVOt4kPx/R9dE1Ed72KdivYbtXtvCiJ6CiebpmSrWodIJAJWibh4VknOK
jC6GZnM8ix0rXM1iTc1+iIR5/2keTLW3qYuUN7n0CXiAIJr1TlrdvrqmHBuZvgDG
B6jsjG9SfVGhodAcEGv/u/kBheXiRo327/l8zUTtCRaK7ZaYTDyejdXq0cS9VKGZ
0bCGTXO/iVv/x4rCfbS3UEFooltrfuzeeGXL531dqigJGDuKlfAe8n8ha2MIH5nm
tPn65UlKZLKD5UwYzizirYsfSmKaujBmHoiflAOKK/Ahtaujo1QW7VI5875giJOV
Rj9xSNBNde6VOlqz4MkUHYGJLGo7o/NXrsPxaFcM5jRIS5gL1kx22HmzliC6pg1O
e6M5+qx2Yc1d2VOqPanePnN0Zg0BTTZgpx1IQUOR4OjnucbXLXUYqg/pDNH2V1m/
oN+iYQD+54yFjc2Bd20YzRXEwWQj5S0NCRbj1F+JJNpMITC9CH1liE5/jHh6FiqN
aVZZpTK7RXNLtHm/tcyvGTePgbg+kwYCviOIw/Scs8hRdC3Q3ZmkPb1PeCLyYA9E
vcwC7dz2n2GwF5SCyiPIEk6xzGSmy2OEGyz+6gIpj8pn/vXSanseDRlPV6iRk4F1
r7i6coscjiekMTdqYhLHAnogpOkCsCLunZM4joBk1fRAaIygCXLtyJyqMYQO1F4P
VWkY9j3Lmdwub1WVexoNhumWpOO4pZmIy9QxwP1TaVSSXr/up6XAMeb83yPe038l
F/knrp1uodKLXSg6t2ZkCLBUxMjKu32yPuYB4lUQnUzLMgpfr/RW47K3+e6YK2u7
9eYGiwLhPJzcyGQgISI1m8fLlM5yEzf3n9wHeVgEGmVYEEQI00xySLYpZUuVjeLv
2R+6UOz16Bxsd2cA0rRztNr7Ja/tTZB/cdbKUkeiRTPpwYGdxv+v+nDOexMRFHWl
Q75fswstzJhbpoBHTkWiU/1x9Iy/gxaOZ+eJ38XcBEtSALwoxD9l50xRh6orWEVO
poPd8BGi63Hc2nSrBIdIUukCFeSWac1pY46v1a7IYDt8PauhIiyHCBhhO/LnJqNI
fiC9AerqpQ15kUzHyohmc6n/C3dOQHWMGG0ZAu4XabJ68c8M2m5mWtr1+pI0IbIs
T7sZFeR3lG/eJzBX/IzPRm2nCJ5WcrOOSq7VHOC9Nyhv0QYOppd3G/w2umsOaC+g
KZLfADh/O1Zu9GxtWtagt4XgEsK+byCm2lUEVPPbA6WPEB53lJoJZWAAzTO4VKPy
t69N+7xEjW360CdSG0/WZW3J4w6V089CH1YeC1qzIAvuhtmEL62s8DSHYitB0iYX
eQXSaIOT8PaRxp/FrJI53ETfi8XE85oQGr773wGCA3h1gc3NCKwyWIpSl1hfMdZT
bZHswjKmZfBg9Iar0EOb3eLmme7FxNfiC53N3LVc9vHtLFuEiqlruIw0i8ZhJhMI
s2fecT+PCgApa0FUs74FfDg5uby14Xc9UraNS5IRVlP6o8e3uH6pVbQES1tScz9P
UXcBpYhxFxvhzIJiKLDik4ICa4AovtE7R8yyk/Bb+x3sJnWZsUfrabHwNCoUS20G
5b1NZF6tKVWTUlLW/wesGXTbI+d9ZOhJC9n8lzmudNGhNYziC8VM/umsDv1Pp6kp
0Xp60i7zOwRXRK/xUmO+eGtmqhd9ZJDakdrbpSPylyfN31EiLRyq+O/308mLv2Vu
qzND+cHLf4gAeFtOev7gsHNRWhayX+C/NcM/f9D0OZBiwcdhTJlVMasEELq/yTZw
s6UbzlmogDK1e6qeYJJ060N1JawRTVUFFmR02w0sTldBnia7zwtkw3IJgZk8Js7/
6Nlz9lkij7tX+oZaD0EFz08d0sv9gKVpZngtIiNAtrVOAjl/hryZWtccmOKDs/L7
KQQUNPw2VRACSNtao8+kCPG3ICbjUv4eu2yQQZoLpBc03XTIuPGwV1ingoWAopGr
/LFAMbg8KnBh/T51V4v4Q0nA+rPLNkq/LHCcTV1Efssxj+idql36/+zSrrzEfari
l0xa6dveyfuQFZfCdZ9XzwbxYdvpj1N1W0V89P0l1AD4/3SZtgMTWpDQp9ePZuhN
JG46/2w7oA2IlmfifQL2MQZocLSWlz5RCKcuvlfU5yjUKA9h9C9Z04YknjVDz1GD
DgnOlRNaQVZUQEIwyR+ZGwe0tv9RIyBq6bvENfH5ZqDCEZOLYdRcLQdlTtgfVS3p
6OCi/4DLlb8U/Cv/hKV3m6+ZcVHJfsgyBBHcLcVxDviDhykHd/yn6X+WjECUYKWG
tFWA4plGj4muZsMKvZBG/gJHobsTgVE9UXepEVFZ0MCj4lG/U5P+KnCR5e6vUsB3
UmkAonDoNCHXgYbo9GA5CRuPZzjjMYUwjX/3BIlCdEbZbY7v7Z5t2W89g4XgaYep
CC+OuQjlAjBufXS8hNdd9yPmBOZApF2r7E3R6+TpgHERIc+O0AIHLZCEhav0e7Du
GWKBsEZW6xQ/xaL4beVFJai+qbO/6HzE9XELo2V8KOWNfI/1w/biaTEhXRfy7eSL
s9oug0iku2xc/sOJyG84xY2k3aQ5D7In3eOqjDZLL/BhahtEXa8bi/AENtYLHHTt
WBxcPtQYIPd29Y4V8p5sSj1j31EucA5WkRGkNrFU9AJwb5xFzdG9YlUnHaCDedHe
8QYJrQKqBAIy9qrBnx4c7F6HQfCJZgVlFnpBdfsSN7U/FbouwZ5QB3eQxi/G8iwf
b7dgzdSs3E+t7770z41CrnOh1X3lOBMek5SnpNUUSJP9fuYzzQ0T0JIwhUj8sdbu
2pnh5DyPLnMw2PuqlkvISTaGK8xSGHjt11LibTzt4JAdndDKIpcMhn4JEgQeeXoW
SJ1chJSUHU7tuqSaA87d1jBzaPAMJqsn8TNUTWFISfXFTY/couwh3iueB7pGTbSU
EMZ/Axa94G9u5Rh4qKZxu5Zgc7V/rTuN19BTWozxHlm4HnOgbLcBy00/CzFBTtGu
EYulgrIJ6GXFaE6kcs46cH8EBgt6xojHWoiP+ap8jzk9JxCi3jjjJ/VxfuCL+psW
VSUiauT0bVxuTxlWdd02I4YgXgf4F8P4gdVN2t+amtk6uz1DAKLNaVt3hagIlfkB
dVIw87lKfzYYk9E2Ct+xFnX2T/RoDylCd2Q7CVrJR1zgLi7ckfE5zLFs3HI72km1
qkuvVVWH3LqtuJwhw60yMJETWxSRBefqnaB4ks3yvO6c2HAi7hbNOJuB67E0CSBk
PuKIbLPIV4d8j0GBiCot1ozIOgmO6UVovrezL0y6M8pggqEPiCseChDU+PSE68Zx
0lCMJziN8aV+DccDZLUYNvo1drWWJZXoCpSyobmAhNIWHcTE3CnZU+UdhYzR/xrs
Tq81AP8DI0uNrvsYKt4kOvgz39kFcgzqxucNh36vn/gDbSuIrUUGas/lZooJeUOz
zsVlnkPpdLybhTnJftgubEaHeT+gqplctZOiNPRE/GqDyCNoHrK+YUqlmaM8pL1b
`protect END_PROTECTED
