`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzY3mmy2hm7wwtg+jnMMfHoID3cLc4yHNMkKUk8PS/l2vYQOjVaIoed5ORMRcXCu
zP7XPPGAFMoQMsw9oF9+Js2FhR/LETKgIZ8taQVZYptuaeGPwXYP2VWTrCdsv2fO
j9Css7Oh00/MaEBjFy5z3idtkfLr+1zD6cDhuCY9SOpt7uYBEAQji61tH+II/HBa
E61emAy7Y+3W7PNeWIbAyonsd57gjtsdBqUIzHEwGhczZ7fd4WRDZS+ngfgQJQ8s
UtcFvk0B4AdnDkbjPzWeo9vSo8cudCvyMyLd/2rXfoB2ZYVKyOKx7fGRCT89bcVD
pMunzcdsfI3BSPtXZnWtm+Lie72tmwJiF+1Y8GgkkO2WmL1VWfDkiWmz1DlQwC4P
oo7cjhkG1DMUx59EV9rgNYbT54aIUc+0h5NIVmuST0kzzWqdYPMf3TQMwY4joVHH
84VQd6GvFczlO+9BlEYkjFjgzC8vyQkuzRoGUkCyR4/sLhCUudZCGW2MJxV4VVBP
CRFFmjEcakaJThsThaTGpGhI8xcSVUqVBYnTeCOfDV7fyizEBFbzc3SkOplxFYxx
uRQmp3vBWcR2manfkWwu/1sweLMLvLihSWR+l+nCpCk4NdjyuAwqqtlq+pt/0OVS
SOoJVe0kenYUJfHjUwJ+kV5m8JnkZxnxcVyv0FaRWwZt+tmxeWtZV8EBCpkBGjun
iSgZvVbE06rhQzBS9o893CW6X4unDkGyShkyDh9dxL7sKq8TNx2muVZlZmdv8cf4
ZH+CsSMjxsepiz96kohWMpWLcaDtx2EHZuVMMCqrsQkCdZbkiVMdCE5EBfrnWl3L
/Q/TOdsKYw2IU3ZeO2RB6TSI4XsHYGJBZSer3EQP7eD33S0iDWWoQbHBmMDc/tW3
09RHAgqtWUPcK6ymY/HGfXnreb18CUgCoZ5WhW3nWLF508V3IXP1WaMrJ58qZ0Fu
QcAWPSn9gD4JGl3k1esVmb8S+sDBUlXdQAEOmUSMPCZPvhs3m0klxvXH1oz2XqCB
Bhz8r6d7RzL4gr699J8vWeJaTWgITEynDaBDDMOpAfEfjv5Cf4DI4EvDfB3axMLK
eEEy2RXgf88tplnFS9zChAvxQ6f8iyRlQo+HLxZpQABMUNDYHVC+9fzri7E20uIf
IwUwiCO8+4LJAlnHRI4kALivZVYSuSezbUXPfZiCne1eZiuZ2+CAwkFEVdYQwPxC
hxX6v8muu3mRidgs7a1d0R1Ul26gB9r/MrF6HS8LH2KxKquRPjnZ70sZ09NElje9
TvWcmeZN+hiQly0Q2V3FL6FPEtfX5ig75HloOcI2OHf36ItGLvR5srzvqkNl0m5b
GxUw7CHpnzek71yTDnOhK0qShwx6IXUQtPdKsA9OMR2p7sK4388DRHDpFRn4UrTQ
vBw0iwPug13xlXADBWfce/EKT2F6T0O1HVtfjopX2yFAZjJkpyYEcVf21TXP7/hI
`protect END_PROTECTED
