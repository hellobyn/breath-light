`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rth1fm2+f3+s13fpDp7xK9szAJqpe8hH+fSKoYFv20qSLenWuAhvqmZBUDUyBP/Q
iOvo0GA/q3iIhjR1A7Q+7c/usQ4IhYWlhWDeGiTp3NBTDbQeavODQvk2G5dBjbEu
XrC24YapFZ4UA8gbmammRbL5xxxI8k+QqopoIV3bb5froA9pdyTRBmg8HlhU6TyZ
vYeSqPmyflxKvUgyclG8883u0HHkQHDBdfTai4e1Fkk/y/ksFoNMjoJLI17o50PO
j6sGV0l11/I2YJf4Zk3cOLGSBv26aI/uUtlR1gPpkWy84rSRTorbUMfRhPo7JI7h
twiEYiItphX1xKfUGL3l71o1gthUZiJ5ATJBSaNNhCQ8B9qSjqBiD4SxKx97S3hD
EBJ5p3jIoJgdh7c8AuYS2tUSFItPROvLa11jyeOLX9EECj3hS1fhTUTc69gZTYjM
7/sc+b9gmW7E4FX7t1s2j7k9oZnIjQukccNqY3lxjPnACcVkTlGslBK18DzbFQvs
6tXngOBSGKwt1uel33gWBHah201hmkgdXpFWjGUdpH7YeGGQfEtQKXhOcIOwTgro
XlEJeNb7O0wXQ6KM6Q0ALNs5uUZ7yWeEQDL3vfR04fcsPa5yd/mOKi9VnbsfELOM
SiPtEOyuDQAc1k2IOZWpc2Uca3EUyDgZ9GNKwRYSd6IU6nLOC1JuFbi4FRCn2Ljy
Q6Ay5X/2P5UipPjxP60T7qz2jeZ6yZFIGXOmkMOW2/JxNHYjdlQwH61ilKxsnX5K
wmArDdk/q+kGeEk+Hb3Op5GJVPTM8HRARcNpHQ2Cw9ghF2STSk/DhSMCpRyI9uTE
a5Ku8CmTNkW5oiBpCCwQgDnZddY0UdwX5PWc4xdzjT1TUrwiUNY6yy14FQuIZXPk
kqXOEr7tfzkIxI9jWyYyzGEwNbe0bakLJsy9Hz84XkqelUK4BNgpskjf7XN/GSnQ
YMUB03fgHX7ml26xh/GL7CYeFl13afTroPfcfACmyVTXUUk0100hrwKMJh7FgrZs
NEElZvmD4ItNROjzAeRTj0cv0O4f6xx12thNIwQVWWD8/TPkb9Dc/02NnRCTNkg/
z1FG42g0z+c7cklKE8O5upMJXaD1nvBcn4MhkXpfFA2BQHrz4PQzjkStV6u3QLBy
QagiSK/w8Kp3Qsmqpx/KK+X8sDj/CPfSWzoxQPhhmt7HHxF8+dbvua8U4GeQrKxX
Thqm7MdphJC0xSbG44UI9Itki200Iw7eQWuf85Goqim+kyjM/iLnDxUa9bpK6bfg
H10aifyavlkH0YZ7VWhuIY5hw2KcpddnkfCZjuLJO2Ndh6rU8JPbIOuLmr6/Xtu8
c1vwT0cEK39Ge8UAQIRn/ppDN+fjvR2QQAaKt0S8um308FIJwF5Bt0xCnBCEyZuE
0RDyexWo7Le+kgRrebML1/jgWekHBONONApKMdhf0vuqcoa/jxkmz7KfKBKwHGVi
`protect END_PROTECTED
