`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3qjckq7auEkYwaH6mzQHamKeHalSF9KgYIt0E28RYZsMruUKecW+H1YuUdj42y8
96lheLg4r5eKuxjRnGwlKSrscjeFJW8caBkW3rpFiT2x6VyRnawqeZSfhW9KLFIb
jVtdZXhqjT8psh5qTS8SXclmvh0ganMdulxt4bK6oEoaV/okrxJQItzHpzoom4Gu
VJqEO3MkqXZhDOa73hlZOYhqLGZsRiko6GGEkvPPpfrMheiETnhRA2klX3JTTeWH
J2MFSzCu9ZAgLwAY/HbMaZb754VsboFK3vBTLK6wmSf28bOsjLHYBDxaHBI0o5D0
z3/kO4nirq0rsl8CobgkWIbcDvaDZbAklqaxXpulfJWXmOFXMdyyA2XOjV0zRvJy
OlzYqQaDNqdE+UKdbv6fZKmWk7m1oB7wakMFWzeypUjzJvfOcA5v2YdassZptjL2
mrIvylLZT68h/Tw5zi6l84WHm6qiierDdHzhv9X0cpMbAOdZoM1MylTfAq6zzgAu
bObrMNHeGXM1Ecn85fL7tYlnOjq83mgwqRysEhKP2D3vaX80nRVpaRS3qhB/u2zc
Qam6h9zUGpQbM8OHd7g6cHSY9RQJvYI/6LmCZ7Iaa8SM5RnQc0OFWR291AnBWF2R
SyIkG3MMa6RkGZeY4fikgXEQqs34t/h0TY9Sv/Xn+j4OnmH34HRjowsvtfwf2ZYV
/V7I6dZXkem41BGkTQGj1Xk5vQ87VF0MDrw44ruyFryczcTg0MCRdch7S5Yp12K9
nEq/WtwGoyGsE52VSCXP1lgjkKM2U1N6DGRFcwUZ5j9LmzqvS94ob9HMVXGmBKh7
xKiPIcSKe8vJONG9BCIC6Vt8zJRg2KlmRp1YTSLlEanbKnEEMRSJjFV8yNq1ix8j
8BQzErDPaqB38izABWOEmGt30edpR+Y148HhK8eYZ9vJ3x30RUC90UnQAs4DlzEO
zK5Y/9ViJvPRryYc6cTn9awtMhIFnlniVmnxzrhfmIFV7sXa5OYnplwdeqv/JpmB
SLFCBTrGyrqFhvGOQ+opvZfd6DJr8u9/qst74wr/xDseMjqQ6LGi3iWgJPGyeRp8
u5yfqiBoStvPorJ9Dcz9V4IPLj64RQsbN1FBcEEbzytmPbcg0nbgoM8iIwJFyqBz
kPKQJt84+IC8s/3QRWLP0Qvo4luisp3K1nTpDmdOnSYkEc65qykWCg/G93DYYdEg
awdESdqTEEonT1rPNwslLLQPq44uI4acHLRLmkJ21GvcyoKQYb6wx5pSmMWF1wEq
FpamdlzuDIiTHT4j6246eZcgFuc/NOm8siK+Vd2ePdY0vAZn9Jr/fsOlKEyzCxsF
4mYsr/gtfueaqbksoTtYq6mfbUTxyYgJn81nznEDWqaNil91w09NTuZprPmtXkeX
xIg/5xheFQbuQn7t8NvwIFRt3O6zAyhzEt8HXdnaOk1ZSp1MNKN7ubQfnvHYKKKM
C9jZJdcbIv/DthGpsQOYaV5hK8Nb4uIATNtURdfVV60wgyLDnXANQDIM9wtBuo77
WPC2nsAhTM7eeMaxKv0nJuGOOyNb1tyCvdjxiNxWNRyGAE4Iom29WqGBqTru6HnK
fJkEj/zwGg35XiC20TeuRKqW2Br7cNlCs88eQ0FZe2mSi1+9lAxmzo/oFhVLpF3e
0E8m/3EiEqZ3NTlinX6zjCI/UALt/jgGJX7KPSxHqDAOSO32w5I1yp/xjiH9HD+d
z6qoAKls//OigLzFMt+ywq1b67KNW0GQrS+Miq8czSUfihnlsCtzRhkMccPfXTyS
eT8pIsTyYkMHFji0DGGXuPCuPrTMt6SSm7vwGySyzriP1xr3HfYcWH/LmF+ZxEJc
zg94JYBj+uB0K6XSNtMTXXwi3PVXPBvsaMrkoDHWEOUPSNZwWb1Vk+e2j6DbL/uo
Fju8PTNgvCmz4yC0rkpWneWb87lI+VcFmjHrSYLb91toYsww4BS+Qj67YmLN2IW6
Q2rLDa9sej4XcTY1U/37O/+MdFzgIG8zZhwrTA4e1dpBtnGq7h5AUhSBsJjkY2r5
stIKJUxh424+X2kkB8DTSQwnBXU70j/DjuSl8KdlNrPNTxySgVxD3HzvuaJBbABe
U0wK3j6YUlxeabDlObc0LkGhiNTRAKe6O+w9eBpFWidwWC/YELrxBUf0s7bAhIlQ
DYwuELZAJ45B7HsIPOGSReO9nsFJw7PpSPO0auB5Jecv2c6jCLUJoE7ICtjLwHCT
bNccsg7ONncwxtRV23imJkj/AWrByZKs+HCFt7eQgeeBf3AuoyNjiQc84tHPqICT
2k/qPQ4HTeYvTLQBU6deQkx9KSEpkAoIgoBjWIhV6DCau2xKOSkqMlZYcqjIwsU+
T/18ltoG+5ttrVRNYOq6nh5fkS3KGdGR0OGcEouYKB1nkjL+Bwt+UYJo+BLTW8fl
nHaf9kqo0TJ3CNsbi0C3Q2qPx0AaVsWqJKDMYwACz5CNE4vC7fg/bHlWNcWvmIah
MLJMskSh9SJCXEHR5Ubq+okeE01GeH4AUi39HmUUvIF7VtDcaEWfIn7agpqnujO4
sPvz/kuu+L/SZITBxa8tQSQWQzIYlpvunIW+jVk1Ja8m1tfQgKU5OmwQL1G3q8pt
JpmHUdiXUNdN8V+pcuGX7D+aGbkHipyqNd2Uu/0SneWnDDRkheno7qucZWyatDvH
RaYnGyiw3xmBYSx0sVx5NDf63f8FnOW+Y/YY3+wooF15r4xkfcjArlZYW5KOirMi
IH3ZFMyusoOtvdeoMnrCJWvBO5AwTCrTrNRY6JoVERmzFpT7ikseUyySt0Hl24H8
CO5hJgyMl7BBLZqpvaUeRcySTOszYlnb+cFKEYpYyxyACKTLM9JF8eZx8twUwYR7
ts5XYJsb1jPjF/Dwc6y41KzZmurM25D3rZ8v8v2yE927dbBSwrJ7QCj9DAWRM6tt
U/w+NHYRWMbkOquUWFK0CMrvjwkM76xOlLnB5Se/S7pgLDooZBsbcBZN0AM6wONC
ddELuri2pz88vASSaixalfPoGnz/4QDqdrcQJ9t6HyhNkI235bcepjc292RnOOJF
mC1qFclJX4u16oPKEfUnrGDdy5HaNat5nklpvg0b8E9XreN+D4Mp6k4xHDKz7c+x
AlDewxhYeBSXPiTpGLAt7zwx2jJl0ejoePneXR5/zYAk5O1Hk9RdLHppCgV/rJGE
Q7E8ecWQNlAueyTmdFMk/OYRECb3VAgtcD4SF0a4YVLizTP5B3+wESeXBRy8Mx4U
ZuXO83ySIGGawRKTMxRbYFi83Jkt1t3DdP2rsGlzXqrhdWh8SuurTOeixnQZQgp9
euM92CgWZi51PDlEtHc1hNNUW/r3B012hgAbu8DXpB9ft4yV6F5/mTlmcG6Qqo2k
cOw8KFougm06XEs9ddzfLlOIXQxVAbUtcgwCVpPY54ouTy5pG3hFvhShVZ1Ge4HY
i9FjrVul66F9+1MTOJpHqZS+nxNWFDN1qTSPWy0b0qf8tgT/0BrpOXK5wXqjv9sl
75+8kzyW1Ft/M2yk4ak1cLhrkxJ7eqErThRrj8YprS95bM9uiF70kIY6jGAiRWHf
ROggk3LEZwX9nSwXhmDDnmz5VrT5vcmH0lDNUqKraVpD+5863uDE3+Z4bNPz0kqW
WCVoqYQwe8PquNVHzkwjlnGniwCtKSPLnIS5nMpjO1j8sIOJnWCL7BckyB8vj0/e
ZJYnK5D4qwM8s06/9oQj1YICIFiGe4ccrpnRKfnzRr75MFHsLidr8mME1NjZtcgr
1ZdyL2Hth9PFIbvg1K0bdNpiIG2ZRk7Y4tT0g9IGuLyDgA+6NBgKKfrAEuDTy+0v
uXOzXatWh3Yr/cZD4XEBAA==
`protect END_PROTECTED
