`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4EnUATdYvvg5A9lKtGhMjIeAYfM5hbTLINv3CfE8ujWIy7hEUxmowBNfRrvPCzvP
fnYYPEQJYNck+jjkCTT3fk4N1BFyJfgOrKSmh5fQc5G0P+aQzT1ws59TzhTh0Roa
Pv+Vy4fY5CIoW/BezkxBw+uVBKtqt3ZvtzQfbUskkWoUwkmDIvzZV+EhQCyN0KL+
hKoIO6yC8b9LjrVxvViI1PumdVO9hdzlaSnSSVZSoQQvc/spbnIXnkVLpvgQ8aS8
UNvMzoRN3G1edOdloLGzS8o+7LN/ZHsfSIYA720t0t+Ekk55UV+ZVolKfrA7QFtM
Hdgg2GEbqNH1En0mmQbC3ufYln76fhxaBmn8gfd15BeUD5jeTuU8+kXn7LHaDfPR
HykIP2rI1k6n/ajWgiXt5nk7v2htHfJ6tOMLSpTligC0LuuEe4LRK5rp18IIF6Q6
yJcVxhMCuI3EHitHhVUICWoiBvCHdo5i0CGSRv5bCnhrUutB1wxMmmbndqggiCKA
IqegPabpTj2l8aZY0HOfHURWU4YRdsrDb1aLL5iNMyX7ngCjYaRrSmwqMPNtczqy
COEYnefIwuZNXkf6NULZgfskAPCoMNw9WcrisgUghVnNCVID/X4AdTFnNQuhdQ2e
`protect END_PROTECTED
