`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u1/rqfCQ/sctS+pV52Otrh/Iqm/ksnAdLs4/cA1x7zK0yxOC2OhuChf8FOiXh7dm
cYow7zAyGyzXrL58mlH7Eo64JuxJ/u7LDIyHqg+7Lkw89pLAkZndFmsHZjJswbnD
Ss7zQ53EuJnjDorISI0dCsMgz8htXCIWEBQvHu3aiEJ9A6+VxFwU9nNc4LZkeki5
p/A1sIHkvjS0FZng8o/8LP60k4xFhpD855Wt7kZFLg0eZFHro+k3f+cZJgF+yChO
flbbieqSjiGhr/vlEOad05z6opHjVuC4Y6svMH6D0rOXEJKa4M2YwRT/eAq/PYfL
l5zHzatNyc0rb0upocKT6sFRylP756dAS6ejJRCj7PykbALbM6H7IgsUVDDYU8iA
/FaeZc/TBUbQBWrHHG0bFhU073qzA4pGRQrCCspcQE/TzsXJmcj49Ok6XC5mO1ZJ
A2E6aqSjsUpCJtKIFOmIr9nTHiZ00yXaZy707be3Sj13smhcjtG0vVG0HfqtjWBJ
g4V5ZVFAlSL2imxJrMGl0eXdEFkr0ZpxjC057hh2o27jIWjDuD8xFeJeV1NNdhcQ
wLk6jpmo2ywfuuM87pgIEkN37K4c32Jk/iVl15mJgXox/hISlHojQ1bO3PpSbu3t
DFcsW1JJAwuckPmjxTpj9Ugf5IkbnB5UXshxqcIWTF8D6m+rt6eOiS8oVnwnXGhA
nijJTtAPjVrmPygjep+g4bGjnJJ3GArDR1H6xmqaxcwlp4P8xtDU85dpFRXnG9tt
7lDc5YgWD2omDdNatEFy6cZe4crpReFl11xwcU8inrU3p4UQSJ6O/ASINr3w6cMw
hyLCgDI+7u9zVObNw2kX/3fs//aufroTS7TABV3TPH9voOxNeQ0FjN5OS+95ij/O
gTxo6ZxbXLUBLUEvtAzcCTyrCDNIHmozTw/wjVjaSsxQZNOLSVMhX4ML8x0Mouhc
8X5cnxVMwXP1PeCEP9n5GX9z3urjoDVL6unqcL1fE1Gfdp6skGT3k59qQqaEPsha
O5twuYmInMoEucBvFP4X+9vzljVn5WZc/WBblFzFiR3BKHJwj41/nznLCUa5tGkm
CBeoiJj36aCjPvEcCbV29KEZC/IP60tsAHkr4aaChC8Fc/katRaa7sPeKUDamNUD
60rCF+kE4g/VU+x0t24aj3AWcLJSeQa5ck6MJwUoq+HFv//E63FDfqSIxyWLcuyV
BhAyBsfmzN7kzQ76sS1ms3Aurpr82U1QDeyNPCwdglWAI9gwg1WcvHAZJk6zLPjb
2UsNzMWxVF0T44g/09IcdP56j+qqNT2eAbDpdKl0wlDLQXIodDnQkYDgN/eE79XD
/xm5JMFkQ0ScEIafBKc8dvd++dKnpImNmCKixLdIfvk=
`protect END_PROTECTED
