`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVgwzZ52JJscWxP3qejXy3q9lRt7EbHExjPZHlr+BBwXsWOZbDIkCnOPJ6Ca/I+K
5BUAIOVUzfTSfaRndqOpXJoOOSOHQZZoMkYAZeITYfsewZ3QBnIcuUPIqJXKSo6f
JZ5Prxv4tVsXaw26x027rg7lcYfwdby704QfkJcHSeU0FBbPZuYU3nnonDa5eASa
2Kip1Uu2mZPFzNQezNo3ZYtdgwfw3Z4av14YyGINN/6IfJRXnjUej6hMSvWnSc9G
GgLSY2YZWvOrkVQq9e3c3CEUvYYv4v5IFRRIHa9zSee0SEXAEOiliItVqUK8vPg4
e1l/kg3r0mpGgEhPZQB6FcVgNiUqmitMKa1gP6opfxW9TVN7iSTIFvrtJaOulJ6+
qdzcB3nmbI0QkWF9ZM5ODM8AYRRQtpqyR/C42Mk3up0k1p5AAGTh12gY6ZohNMKS
gKcTTgISPb43SXmPoypj8YVHIPZn/fuSZvMkZbC0UIcmFXUeII4rYIO/ZRKcuK1s
KPZDzQPvOE6RpLJaHzUc5sBnAgqIQVX9pacwOq5uJ9KvSQYN+hGB6T4tAJ2wGWS0
vBWatkRiFt6IQk2PdbZmg5AGIlnyQjDT6JWZm67Y6J/Bk8K75dYJJBoL99mr99W3
SXoHCCd0fCaZTs6JVTa3z7ZZ8MW2tYpDi9+BsZCF0cTLOMfoB0xVPgZS9b6hGEwc
gsWgnC/XO/28xMcmVUThiswHGqpu/niVYVKxhvz+wdcrrSZnm5+gr4o7zOppDJDo
/1+uTGKOMG4RJkLshTcu54ajzPrCoyZTiS+Ii+Ig75ewlZVUjl3wzPLSlOUY8Atk
bDbwU75XMkX+JltUCKB8c3fNqjmGYx8hoL9joprobYr9rT6iREpyTRiLuya+HKWJ
oSmNvnVneK/UgJTy7UPWGeEFUhZ3ZlxMyUWu4XSAekKTF91E5xe2chHJBaUglKHd
xhyqxyFTLwPX1ctUr7ypChEBYbUs3bpCBNZyW8dMfcvazH79cbXuXKgr0S6g+5ov
czZUGsAFx4K5Ki39Rg5tfpkIzvbLmdwYkz1NzJtgJqITxWbepCBYpJUHZ1cFugUS
sjq5Y3KzYldr6zTaZdXQGuYjSTQJHMSXUDLCKpbP3eQJ4RijO9S00px0GH8JYLvE
TO2tWC8VeOPNQYZB2C/fdT+sWsgxFDRD1CdQAVk3JhpXRdOm91k3R35pK3hamaJF
PRMNb/Ttf25nRdIKhKkEdIo3rV4f94syFj6eGKiHvs6h1NaxhY8I8EE8nC2lzb1O
QzzR4wQD4mvVx/9pR8psqKG9DVFDz1t1KmMAE21UgxqA99w27RQfNA+kQmEWwuIw
brjIa9aoC7+08oShcU2957SsnJd7M3BC/HH0PomvHQqznX7v4FBFaOxVsyok1qjc
HXPRubLgSaagf+acZnB7dtx3SBYf16xmggd8YV0vGgLUd1LlbyFLHPizxCFMSCV6
u7JlzEQRiFZrR40MWeepbAKPv+ZpRgLTsKfo+RnpeFLReHesbyr/p+NOYyIZJ34x
hZ69eUsP/d2I+XF3qo/0nMDW+8OddSfwtl6ik+LXzI3hdyo5fzXZ3V3GbZnKzKhK
`protect END_PROTECTED
