`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEZdbzh4Z+2V3IhlqJycgu8+tH7TjtX7I8cTmIz6T6V5IKaOdEU6U11YKPdqQMMk
eWigxtq6MNq3EjLOvy0gA94jUp+P5//0D54bcNuNtpZKk6pOXcvN1wSTcfwFlRfW
Pl1Oo6D/tCCyYrZviXXn5fyz3mfwRsNIxX/rLTh2KLS1+Kwkyx+lHkEu4hJFzRgg
hsv+UB824Osp/MWGjJU26420JzwItzMIoUAsYyjcasFGAQBY7Da3Y+PV8cNJ0i4N
+mX6ARuDYdAbeooAUhhT3Odt9aWT/7Xfh99GfZ3BQziK+khl6986A4FSawJeJtr0
nvNOAW0UF1KIBhmtggfuMoqfZnv4Y7bOSLPEkxe3NVkeyrGIC2NOvSKCPv5bPOmi
Do5R8rWv2JDUWkMmA6E+p6D9TZ6EwtraG2dOU9r4IPmSVyY2itM1AQd0GzxE+8c3
xqbAOOP+2dGDjLxtcfcONCDSS01QjZiZ0WC1etjgygQ26z957d7FD7r5/Nf4N9es
6ereiGC/mANRwQQK/XqzL17v77ESRS6qBVie/wBS5ik7ERv0E3Ma9taTuh74NTHx
y99uSwAy8Oti0Ehbvh6tQgnQE6raNnRIRJqDLHMRIcga2iYkMa9LMCjMXEuwqSbR
Spad9VXsypzwUjP9OS6Et6FmHs50hTM+mr617v0sIcafyUewSpKQ6BI5alGPuqMX
XdSL6EuXrzTkjA7L1xK2Y+0foLWgjx0SlrgWwagBgG3UJ59b/mWRUURyNUjXQyYf
Dqime+TrGySLGqdR8YB2Mz37xUp1jxsOVZY80QbftFAV0BbiMVPSPWv0ZjbiRAxy
b10HCBcfTK/PLTxat/olQ7A9AQSDLtm8g/q3sC2DhHqA5ReGnwwiOZ4SPxvtVaqh
4NvrSMGXqZOtLBbPGJ4juWLQSKznLNyPDnvAEiLvHjKh+zYK2bOnRrcsgnLHhtbD
peZ3fJCN0tANP/Qt2aMOADDK4ElaDDMZyAhF0rte1OQWHHhNhNYb1UcPfn5hWpfo
atIhdceHSULWYTIT8qw+61GDQWvXDKDIEmr0sp2LFXjtK4rvuIMqQKu/p3GomTDI
714eng3bP2Mes5N/y6S+yLwR7YxtqdcTr/+cfZSKn+y3bVx2RPn3RkNshCP+GLZm
IlaLcQ47U8jJTYKVBY1MUv+YI3bmHhp+QoQfAj1cKjoA9yGzkFmXVzJoxeT+AA3l
q4o0gBWxDU6tzA6HtvPHK/TYt/CBLuKi+HAeBrWH4Dkd4VIonw0scbvs+hRPD8f4
40Tz0ucaPp/MFIyIUFCZNjqaoTPy/33MukNtpHAdup87ZPFeY9QPBEVqnOLrH0Dd
8Z8yIFCAA5JHVnEcP8UJitrb2N1HgzM1lnkEzTyAI5oX1Cat5b072nQWIIczh64W
1wSsdF/meP1jsg2gh5YSo3MMxUOKSmVMEoo5tlJy9mzfNhc8Zvl4g1/ev6gqmb+i
AVdPtR7SEMeNTslnOEUreZ9gvdOHpIPPwU/g6B9OKi4RFZHKheqPQcXfjFQIoBIA
gSkVPZogQcrYj6Vi2DbXa/9nblm+wlY6YH/fGjrXJEAFsnbitxsoyKfy1be64X/I
yAkBJ5x4HhxYzsbA0//fzZCQG4+Bl+n1lJLv7wDK0SuqzaRlLlMjmlQYuU4cWlmG
JTbKJK756K6yXerCjnJdjhlXV83bA7mDeovQ3LNbCrAv5tWqXaVNdpLFoCkK034Y
MnRkIkcf3p8d3D29d/Qj/77OlOU/hP4zT8Rx+9BopIVX7jMCiDxsNPWhTvvIkEWV
fkSzAxeZMAU5HzVrayVr9RLFyB8dhJAhkwvqlRe12OpFyWjkMHdsSt/MhMo9s+46
Tn/zaJvvERZjyzBbophGoFYGAU7gJLwboaeW90Nd8M3enxPHFbVRa52UJJCM57bP
`protect END_PROTECTED
