`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/eaMqf5fatbbSpUWMwDSHMuSJIXnvh/7dti9WPZPQvCtQKTrfG5iwS2lVlx89rrE
bPbIh4MKwcSRU0pqkRZNrVhZ15h6pzohX3VoGyKBt/0q/w3Bq7sNv7DdHCPyld4k
+ryVraWm2uYOMFI86PKxpTb+g15J+9/GzjbklauqQuBxh1L4iv3vH70jT2GVSKLR
4mVxGWOocafWos+AHeXsI60fdo8fLk1MNJ/32FQP0SrlF0kQT0/N216QMlbZUswd
Bwr2/Ec0RenpX/ZI7Fh7dxpeBDaz1hvttNjduaSmopfpKbzjwSItBTO7Vr0jV5Bh
G0l3WTkpF2xE7F9zUSatESevuDAPNYKcGLoIUqSlSFxvtc/5HhqTiAnYthRVGTWW
h3ZyuSU2wBojTpfh5GCNgNjhRRgu206Hy2Xq9geOUtN8biIoYaKZgL1ftto/ta+i
0AihS2IJ479LpbearSP8FFvEUMQ1hAfy3qxM1/vSk1WXoFuvMjKCwTQ2477TDLba
Mt0U53gOUOmsMVx2jBDYW6DBnkggmHvQXrTny3tutw7SL7xHfiXM/m80JAqK0mmi
dGzZQSwtOq9hB5tXfb4f+OQ1EI1G3hdGpvoQmTUwImKHSdFcb62Drd8ymLlT1xm9
bU1R1htTAAIafwd2tAkp+UWv3MN9kazKEKur+HjL841I/K87sTkdJbLqHzgnElTT
PLl8mz2VEveZUEYYMCcTeOaJFakSA4Gm+SneEFj2iTJ8L/dpiNlr63iX3Ie6hjnQ
YifydJBg/qUwTU7O7hMYlZaGPt7bqquJtgsZtJ9ZGhmeoUmmD8jYVQo0VAKm74dZ
tX/GNaT1SZFLrwIG8WwWMWHEYoL+KX/Z+dFal/bX5Xg=
`protect END_PROTECTED
