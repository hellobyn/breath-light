`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAW+4KHQzGLXBtxEKQitNXFxT6i1QzU34HNLT3AijWuepfNGXvq2+Qyk55872Ul9
rShIGf+yjZf5o1OX38L0lAeR37Y00waJXReDnSk1MswfiM+Rzugpv+39H7rGi1je
u0pDZQZ8zs9B/vcbojhk8aU8tMweEbWmVGrdMwmS7fV8lHaXsEKURc2W1h9HtPUU
hTrtiFfJcGfTrKGzkyn+VQrrZWN8UualMR/W9/HrJWV+Wwx5jfte8NFJeKJBTxAR
2jGca/WCIlPGUfDb+KsbhHCTUk72MdMqiSL/f+1bxtXBaZ2hXvg14nVKw4Kdwu3v
DRiUzh7kvQhX9aZ9jfGWpRW8DrWSwUv1L00Whbj+3YZnR79VB9+x9vLNEBghBmCU
mZk/FzLnzwWUdTF1ZvHOoQ/92M2AF8B9/iHOgb7PPeXAwkYFVxQSjynhfNFgiCjL
++KkkUTtD2HoN2gZAl5b/UnKHwsf2Vbrg5nsOzOQpriPSeh5q1HqZ/u8FW0bvPwl
LHfvb5yTcUoLUrpPsLkQCrZMGRr4c38tBewR3m89Ob5TrJ6IKjZW+0URT24pk8pU
JJx1zVujOTGcNArfuExmRCFetQ+uMXiVc8WeMzpxWxaelOFbjHLihyPtIv5YEWB5
tfned1YnKxq1fKXSZpHde1ykxHanuMKuG77X+kAcVJezpeuyURTPOlbCssyznUnb
1wy3vSvdlijZXA+hCin/kAXq7GlGHgNdXAmo0vHB/wmcONkR8Is+M6OiJzLd2TOB
1g0ubMbEiAvmOErqd7w5wpeicDqR4Ybpnrjxk8OsPpmShxqtJNLxhxcbKMrVNg/Z
qVNt9teOvKtbCxBM83L7Xhez1EF4cM5pPZsAg2DqmQlH9VdWGYUu5U0MdXEDVjLu
IhJo1lcwyXo9UIfVUSf6r0LBdyuf1E9eej1lWeZr5VY+ad03ven7IsxiiZDTjapg
m0R2pY3Bxh5Dllbb0jEAvflOEkHOl1qkEFH2HkTvJKLZQ0umRmIBVA779L+3eyOG
CQjyPQ0a71EEx/194iLE6e2ut9Wta3HWv6dl06SnN8zxi1Ebl+iZ9P2jYRaaxEA+
c32m1t+GfuloJaicugpJJl2BX/E0TV3VVG/jDmRVwREix2JOF4rEMfwZoPkU1b43
toAot2vP46wQTcLqjthU+c/DhTOpIZoA23og4AYzOiDmHGJ40Z0Ru0oHAbRHLURK
Jh6hdLm7Fa5/MO6vBkhKXVBcxJYuOPaJvzuonoTkdUD/MQFVH8qnTBXb41ZFxnhn
qwguwfeQgZ68+Cfd2nt68rqVM26Dwuefqaoy+UV9oYGoObvn+AemhK6f7hU7g+yk
Y/s7/dM8Yiho4bPzRQugA5NlMAmcqjQYCmt3tQHMmLZ2b+jdcFiRoWMFuj9/WdjZ
ILdjTuOpulS9a1cpIgG4TW70F0btI29CWcjFPpGyYu+uxN4VzA7Kmr28gEfCXaO3
SdEM0qFzUk0EGpNH5/ne58HI82NOUXEAs/nsUsbhLgvhH0xrs8QOgMT8PFkX0/Ac
SdejQRm3fSeFll/7TXI6jUMiNSXcWoW2cVQn5XFoRA0eqVsAkpNWHGSST9Yzy5qW
cGIChQnjlNFcZf57+t5yA3xfqM+8E9BeWtVwo2txXGCedoTLKOKZ+pZ9MwdrrDNo
pjGJbzepi3r5yELA06D8vZ9Bt60dHQ2/lUifONoBonwJYYljKuMhDdXEKe2rPoL4
8WScqWTP1gVK7Z16KeaKJOz6FWBpdsy6KmjSsoR+CHY1sAPOOnCRWtsGiYcwkMAR
9TsWpdyotGHscDPq1ufUp65X38YqhxnWKBQF08SoHF8qAPUF5oixN6YXaN1+HbFN
BFV9lEgwOMtLEXUi+aguFIVamPcedTKTel3wV04NqJASkGQXeR78lBVYw2yxHxi3
hIOt41WDBr9jqbFesQP+CMrN3AYZsmElKpxKFnHVl+cDbxgA6pdRvehIJDWXknYX
V4U7rZhuonXhQ7vO34z6GDW4MNeDkhz5BpH7g6gHAr4I1kOM1lhntMAyeP2YfvWI
h7oU2F7KUP0PGcGZuLV2xSXMLbetzx3tNdVC5EOz6V9KSk4PIxfheI0yfRAY3Jtj
Yw++DV9rVnQV+OlrffHeXDVAitlWD8ufOBsK/5ep4bX9HMQxviTQPJZAKOECMFuM
fcx7Ers/7ILTon0iD7DaRFAg+0wlB1bqcwQGiBE8w1k5FDrmppMJf7UjrCjWr+Sy
ZIv5ne2VtmOvQ+Z6Bkd6zOaa1H77Lv9erIDESjcoHhwJUonyTAxHOx3FUdPblrxS
VZFwROxdgl8tuX0QfP3j3YNLIFONZJoH0WWEB68DEnGBIfL/uPXtCt0GhFUAWthL
V/u7foC0XfJ6JdeAAttlWcYpnGaDJ6ucEyEg+mmJtFVNoEZEarluDuCsMOyduFNc
EzsfyrX4WfWh/YdLlJr2FP+TXMNQeLSKfgQpHO6KGYLGEnzWFDKSDAVWPpulAWzl
y8T1c99c4fYRMEUrt6mkpXMVHGlgIECw3a8nj7JdPAxBoBw4/SecLoN52nqNHOtc
0FvwqwB2fOPI9lYoQwvqGg2Aj4wKFSlgxTY8U6IorYYaugH/vAZhhYzAcD/8e1jg
Mw6s9ZYbptm7vF/L5hz5RuwbiawLNAym9XcbI98Tp/4N2cjIRoMzFJhUig09UyGo
pA7WhScBejHYGf9nd/iolFjfP524z/ZDTqEUmY3EIg4mcFDFrHjCKLYhpWHcqDNc
ZlRG8704x29sUdd/fua8fgG2G4keLC2xxP2uL00e8TJFcUkWag7MAIzYjCMLEcfh
3M1KSWZjc+IOx12IQof/4VVO+CbB9MVkcpPIrB5CT/pp4dphVfXgn4oD1+u0u3eH
n0AtHovFviRgxlpcU8cXLmNGJcbIfpDD1r/q/ki7JrQasEHug/XRDJJ5NyyAyEzg
HeUYGMWFuECPxVNY1BcrUrRHqLaI9nV5I9XXaESBnSlHqebQFAcr3ecDfjQlQiPU
rGjjGGzmZy8Zx5SvBxQSEwAHlmyWA2UBjI6Hze+EMmCG3UVuOQhE6wUbDfz8McIC
CvwWsPbhE4gyNxNTEbAI3Jrzrr737eIVcGZa7r1mvUuVrEQISFZe4dkfJ+Nxx4kL
HMKNieS+7lTBpezlOsxFN/UyyaqpE05WXtTptb/DcXC53/++kUZR63C8vY5FssXp
1QOTja+DuMJeALoem1voS2kuPGWyYgoR0o0xbV7VBUORLfR+5eB2lZhZHfdDb/dE
I2CFvPETW6VHpj2ZVcosE/c8ewqQzkkP+8T6CLhJNOG6pYDUSCywGLRr6jG1M56B
Juy2WTtgF0L0BMTu7RABLnHcQR8YX7XUm1J7XJrIaObnymlH+tC3p2fH7yJa1q+E
/S/zV8bqBLVAOu05/q4ROfdpwniUr76USTMALjBVnM7qjcztsh2/EDLIGLWJajWV
9VX2GFHlBYRm5lNgshVJCnjfyKPprcsFg4nhJRGL3ExomkHLg1ZJLYi/1SD0POWs
iVj1uz9uAJ91l9xqEoOrkw2E4vMfqXBitUuH/rAXXFD/WVmA6MSWOQbNjWY3aDl9
FXy+EtWzwXRUGXLF3XU1qtG4A9WwRKY7Gj91teLOMxTHMvjLn6E9aQQhPfsNr9Ym
+EcSumw8biEB81K0y5b57Wy98WWoU+YzcqwAcM2DOeSE6sORWUUUDozLdO8H+lL5
ZFianfyZXziBp7+FDIYHrl8Wg5JCjOh1FyrvSz54ZYe2uEFkELpZCrZ+WCvImCrl
5AnG+H4xxEe1Ct0AbEhnaoH7q7e6GOQQ332tolkdHk1LgTa4Ru2j2lXq5P6WGp7e
ZI3E0iIoOmfdXBnpjqC4+9Nb8wLsVdPeA8aBqVWgtt2GhaP2El13zwuSRg55K3Jd
jWo29R0v5jxnaSM491pNixuiA+PBnEousyktNSLlgy6mLMx28PCTHiadWdonJHQA
cCm0pzLj8LApNjsLVpsm8OLaRn+8v9TWNbVM9aOBTC1JmqUOm5ZYh4PL074VcXBn
ou8hf5Mc925nQfKM75tH4TyhMzFPUYhr/PI//DEMKCF7cnjYIS73FpHUkfD33qot
jdre6Q557iMNhkcaIze6kE44uRF86bZLSbL8ZPiS7bqGY5bGwu/tgIR1uABQ12+5
6sbOLJLhEuJIvJ3UuWcBS7EC4KCXqupD1tDev1PXdzPa9/rqKyLa7CDFhBGeKdZ5
/mdfc9zFLUPPgkbtxjhN27p8Lf81nXUVqZJtmEvycGDCy4gOjFZVCZvL0QhCbbSP
jeZvM5oL2hKOOy1CEcd4NFSxWWv8Btu4qN7hmzC9y3ElueQtFQFGftq7fdL+dnX1
3ExSaRyaHJSFuy9hpMOHlz47jgRr5kltBcC4pvPB6wWsLGOjFJ8en0egPpj92KGh
VS7HaVRhfxpMRBikbVRjmMHkwrftWTku90H/QW3Q37iJz5I/5Ad1rcluZbYY37V9
mUtRBkaRbQeEUVoiJ5Ilu2C4yjJlIEFlwWp4WjD0hQj9EBhvlUfTuCut6jBR1cw8
F13wdLt0GvZwSl5F6r1oP6iLIWDn1xcHeEZHhHZ//zc7P5IbI5/F4SjhgUPiRBPl
0ZZhbIio2LOihJ/uuy7LK4Otwj2rOU+PsCSQn558EeZxMHjd/wY6glwE15AYBcti
HpZMxtQcjurLg5QKE/kg5kSqJKLNRwU+LNLEHsfaWVpAdyRlAgoWnYUTIyvMDcKb
SpFa4Wh6MkHb8WT2JZKE5v8N+0L0ryHlwlLly9fePg/Iw4O61hUUtDtwx48mMnTj
ro7EUfs9FdRUbnkrZjY4vo5SKsKaJHxtcnMInDJIvg+/NfGuBW8lDQP4OjokV733
shGnJAjcvwhsEteBO6TluXSU4I/Rc95V03oDjsIkA8chPK1nvICjmAAzpd0RsHvB
`protect END_PROTECTED
