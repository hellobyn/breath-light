`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCrOTp/rsdxbbpmm8iI0OWCvLJ3NgQ9siF+fC+z0jiPzOE7QL4pyzBmy+gQi8Jk3
hrSEr4ZnXR5Vram2+lFZVrzkpasFW9f2yWf60WWN76k7xVRtVLb/FQFTJJXUS6iF
5aRq2cbCFipwp9mDlwPhWXUU8kYgIvHvvMi9BoBy2Agh/6vJxROtKjCv3YUEKhQC
/mi/25dP+jm/YN+2YgAoZHBWu/X9gxWr6sCDKj9MPh9ujdTwprcuzqC0UEe5l5oa
L2zqJlRKFsyPLSMH1e0GLMZ1wfX5LwKgCsctg4GuFFn1sUcYFNDtHPH63I9w9yDv
NQfg90o9OfuNlCjVwvVsX0x9rAtUFqXZz1Sm9jPlID2aF11yvD/h9BMhovs5+j8k
ATPTs3DNYKiiXzXZHYjGYiAnyNobjCVX3Zy+UkQneXAjk8mcMqMsnZ1z3MjGPTuN
y3eH0OMU/4WnQIDgmNzYqbx4WXGvcL/1tVNGpOpaxLqMZgnr9HXKjx6v3Rvb/0GS
eVjYwZNu6pzxpvoLnGN9e8dkDDkY/hFwa5CImmMvZl25cfByBT+d8ZWngeaSQ9v+
pOtFgLIn1vZKz2yQfyJsBhUbcudu2YEAuyJahumzq8TIZNS7jzf1ZBmsxi3DBYwq
WwJT0WATxV+ohGktJbh52cKmVP9Phk+0e61QLowYWkNlXaROOp4rqFUF8d5vjKIL
BZFqm/YYJdfbeSz1kHM1b4qlU4NszPC+5njA2LJsCFeaqX+O/YzLxkuvsFxTX+UG
dBpvCI/VZ4MwY1GmHt5xzx9T1EOD9M04pos39aSuunzA8Qg0TsXiDVbaWLcGq5zZ
xrzbCafmPa9LiDhHQzGqi3SEMnB/9NYunCrp1gONpog2zgnGQWcO+0aGzAG1BCrx
IBUla08JkpyTIJtp+k2UQIWIfH22iAUHaC6cfA8nnkaU0o2+Wsbi+H5vWlzjXlnI
Eyp9shyZtt7a2X9JNp81vNU1ZXlH/sGYG0+TC7Q9MinP+Gq/G/lTSlVhDhVwlhBq
Q3o76MLawDaf+5CItfDaWp9fO3Vcdi3hMchp+ea0qEkZwcGPSPJtuGaIhdTBvdxJ
3+F3jsxjwdiEtMeUsWcq5oiz6h5kRYO5G6muXuraKHfl1SRizwsyUkdYbkOvfcCY
U6M64N8LA8iRfGT9BxBPW60N5zWy/auEVipCne4qAXQP7thaU3lHjhmuMLKR99fi
+DJLPe9UjDzBO3xVCKbIO2krY8qtQ5jlkJ/w1LwMjFtIt29V/idA30fRDTED0RuK
teBMMFlQQUqLZMLqAARvvg==
`protect END_PROTECTED
