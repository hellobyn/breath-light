`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dALK53cJnbAWGfFc0mqUekDsxAJoMXyLZ7YlF5ZjfX8YFvJsKDjZn/dUNq7CDaad
X6fuOKoQYXF1n32nQklXw/H9ACn+4smg1TRBED8o4924Svr+rfvxR0VbpeJ94IIJ
NXUQxxzlLoC+6TqKCOQ4TMh3yqmxz6mZ9y9J7J0DO8sYVYUYQ64vSkEiaCHno9er
fZw4PMvj1sC5S1ubz/uGhAgmqd4RyrLbkluH2vfHFvWXQHLvQc5cIH5ERayU9zyo
MTDhdurzUylpT+Ged6YG+B8zm6Ym7jDRobAVUTo7zjGwlhkjNDijlpnBQRNi/Dmn
Zjx68w1ha6yEPIWg0ConwRdqQ+bk6GLgCQJlrzJFNFxSrwOXv9MZmA7u4MimRSi2
w0LL2BCgzgQMMrdqH6WonykoijqihmFBf6JjgWT5iZ9wTqRZrqxNz3mkPS04uq3y
fnQd49L88yo9w3FOWwBfWgvjzrKUFa0A4M6/9NHeZ0x2KEpsHb58yfwm7Rmf2038
J2l/gbRZbLk3Nifyc6FMeHs6A7DcUH/QOxwKlhWd0Qb/StUuoD5m5eEkRuTjmCx7
g+6v5qUQsM3VWkdwOUrfm9F3lITIZfY3WKE0glQ8YK/EDZe9QdfFSKvKCrdfcgqN
xBaX3jZ81dlBPGg38R+YwJYZeRar9oA7TNJOlK54oKoPPj70DWQTJi9gfCi/hrhw
c3unfPLFMJ+FURVD6NA5kudtk4VASnvysNdcwWaSeo4zOtIZdmf08i9UShzNSf0d
J6l5xkI7vcWLmdpTPKm5sBrZfmSQZII8x6I/+AaNoWSFrkVjvsQ8Vqwhv6MuVqi4
PXIv0bMgX8v4urkT1d5wCoXL+30P/XbH5+qSHQ5M6Cc0c0zy6q/LSFsjX9wReAcV
odMZ18RaLZTbsfE2LzfxNmapgmSyd+vhnu+4BOnypCG0z8dBbAygpdbtYnPlorkh
INSn2Y6nwaBaO0pnwmwvTQ==
`protect END_PROTECTED
