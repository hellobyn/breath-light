`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNO/eUqNq3sPsUJTlmcBpNUbFYh0cE6wBagoDimbu75ncZNWGMY+8bS2EGTyFsSb
XrdIjYxjrWp3z+12ZGM6TtB9MgWoJsShEP+S4d2PizatsoHaPy2itU/AguG42lpN
qIRfVBR3+MBgsOJPrSZ6c8IpLDhZd3tcO71hWjhh+h6V9n5yEu781RAW+jX+2ECI
stOS5pOel1F7TBg05EYvip9UP3ZshcOOiewFJzZnHLcoQHjE/yY1qatYVYWboMP3
7UaN4/o0HbAgFZlgIOoMNZFDwey5QJaWQ/Cvbqt1GhyvzBRDYDNiytDJKMAS4R+y
KvrZxsNb8YIxCdP06W3wvRhJqmB2/ihZdWslXCuSUGGqnXcG5OZakUoSXdakvcHX
vOM8kKnRzYdXZxM2tZPvc241y+7k0XsSfU18BNVuUjzO7OpVU2hok+6Ii0KN0gSz
tQmQrsTtIZxvt+SQE3sZiOEAVSAJrU7fdUqK3aCgt7JH1KSQerDjAJP4Ml9xb5wo
ZEN6SGgCcF1IAmtV+v0bb6FLRixR/kdnJtuukDRLc8hzfRBFDWB24dzMVmwc6c6R
lEDJxWZfbuU7amEeifOhKnOl1bY+4U0aBSL+t51aPv3uzTezz/A/IDH3RwoyE2s6
XpZ9CatqWD2/58hU7WDpMnU+BzbK5iGAAezwINR+n4SZFKwhe8KdxjnQoktWsplx
js5T1u712EF1xG98xS5wXVM3fjmmEA8NUz8k2c4Ag2sM9e/EwvY/wtmiRxzrIpE5
zgGV17idpJzUZaJjYXuEi2bSe8LDUTAl34y8kgqx4XLJr3vl7F5Gv4RdKtxvp9aO
7uUw4nmQS/ISBHPbVkAI8DP5z6dmj6L5e0gqB5KkgPjQPeD6uv445FICxJ/LavBO
rd5ARLWtm7UusfWMsojOWl1s9E5f6RQFxnNeJ1F1vvtC2hT1FfO72qXmijOoFXcH
giTCgsI1QNYODnx6fwuXX4+B5BkbjvbW4YlmHJMkZRvEHbKb5Pm5+zBKUKhx1njY
XA0MBabFqC0Sf9blzU0OASw2Ymap0jC5UXKhEaGUSmfOUhCql922ibHXifyJOoQ2
JnmGDpJqJJPkGqlVmWsKm71IXHf+NoBv+61uhPVz0YJK7J54NHYRW8QdlDeZCsmV
oS0RVVwqhDVoO9gzLjQiC9QcfAxuiOv9CyRwL2cJHust4ZNL+EprsbnY4qV7ZhJt
82DLB9X0NUUU0+L8wV3rUtDiL0dZk+1+Ow4a1THXJO9ar8IOKUvtag3oIXvIiVZ8
`protect END_PROTECTED
