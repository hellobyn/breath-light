`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRTyPldu1ezUDSX5o8D6+2P1oj17s3J/nKA96nENbP3NYWJr9trw9XvP0hZMZsy2
Ud6YEee08YnJCg3tSdehtFX+oXQWqTOc98D4fVHNhftTg6KFdmTkMyHI5xZie62S
Wt2rN50ayBKcRcqaeWCkvVvjsQ368Y5EozXr7rbGp7z6rhsn8Dsfl/K/oidGyAuR
Oes7ZkZ+ZuzwChbQBK4cNH9Oj3rh0NJSXV/wEfEXQiLyYG/jilnKV3sAf23VqP2j
YH8Mi/YbWc7sd3I9vO6GmhoG1J+yYYpltd87V7sc5MEEU7wq7FmxBV3+3lBKW4C9
/xpdOCH3PfNsQhf58JTcvLB4g+fIFrSG3Z8ggs443LZIovTJEwv5vhAKH8pEn5iE
PwJQx2Z/evFZVdbpiNuBOIGBPlcsxQd7hYiKCSyCEwtt5Dk6C5L7uIDCVqpeBugN
C/ZYA1YjWvb399cywo7iFYTkgacbGWCHTeM2tDvbWDwN+1eQmlQ9phxf+a/M4WGs
zSgNU4QV5Q1jGmO0Les8S1FDK9PDjQlBJTngAPT0MpRno85U4yM/Iu7P92K3njtJ
1xEr9OiewUSCS385/0qb62RbgAC+AlLFAvuyJrbMGBsLlSp+498t8cPFgYXqrwsx
XGaWl54KrRciMF6rf4boLuGPc9zCSWYc53Sv6tsAUFhps7DSjKBdVwXBGWAumqhV
xfil96uH8eg0iQIS3o/76jQCH+hc1KBS+8sKqbN0W7yJ7Wi79bFabaqRQaMZU3b3
neM/RmzGTx5NyWg9c7XcsZNvZ/nRyiFS/8cMFf9cM/8tau17oBosF/YAZPE3Twrp
+9EKQDFbhJv6P79G2jRV6anvJ+TDUiVl0cXdrxvqdmQTKSionCUNuriko+PXLGy6
gThTBIcsoSjxuLZGsDBQk2TrwUoOmhyGYVZxe+Up1BzUfWUGGV5QRxewFcussunB
/LPz1pWsYKHoHvylAZqMa6FQ+XMdsT6e5kpAzO1vtk8+M89/WWwOD7w8zS08d8La
I0hABmsTPcWQoqXjbgYEQ1lXQ53TTgZj0Wvs3gpnwVgddzBp14nwZD18ET4ZoZG+
JeqBvJu5qwxeKMeLY0zFePEddF5sg958bK50gBDPdLUfThRX4c4hGOM2/ZdzG3N8
YyAhbxVVlSC4kmEjeVKv9UF5c+3JpLoc58/aljvef1BONtENPxI/h4T23jsT9imJ
tvNEno2NimUY3+qsXYbwOCo3yOlbXt087gTu9mNyX5nyQNWQoY9j0sF0x9TrTP3I
lpeWCs5JRGXWy3s/poT7sDglFUfCaSeCrBRXYpuOzs4EctlLndLpx9tXgZkPG7/Q
/urW3snoNNKKnmPV3TGX4UBR57l8CRlyQ/Q3h2s02Ze88YZiNsrkVW6kX8GrHvBF
YuM6zfSVr9UTrIPUIee0Gum2VpXv7g3W96GqYtIg1+IxtMZTRzYZQQ3fno1HvceW
D4OPzpa7FAXRA3DCEmp+sRMDrcJpCaWrWMX/FmKCJrXU4vPwkU5jiOdAyZMmnvqy
fDBywZ6oFxsHxDeXJK4psqa5UNFAXMJ4sr2+R8bAJ8HsqgqslP/f2BN5xUSiR9PM
bE3U0JQM+NVWkUhoeFrfs17fO2yIDqKBdkOxPCe91vaIyJOghvo8g9zVlHBqphTR
UnlbZa75cQ+apo6FP/pe0jZwJKWTzN7YjUdQZTGeXomxidd5WWTp+z0ScDyN1OBo
Lti5S1z9DmZLSLBrUTJ0hMqr4u7f/LHXqRj2qppT+xG4tqV5hHH/5Bbf2Xt3Pmhx
Zv0p7XteL2x8VpEcDkkx6eDMybsFju64Lqy1dL+8IRc/mseh0v7hI6tJftG/r4I/
o+Tqe9bomN6/bC/8mVGz5oLgjOzMBJwl+gSIBbDfPEFbEu0zAkFCt5NumqdXXlVd
IXQNRejPqv+EIuZ3KNv6PyJQZhKbGeGCpukTwUgwiVUhWND7eAoTTDCBrSWsqm+B
Wnz0t4Q61iBCX8hYCugODXHsqNomsttXybUOxEea6+9VrFlavkhcv2nNeOokFuOw
hkByWvDftS0VJhHiSPoCS4jewLzAkn8Q21xU44r/H5qmSKagiw4wxp6lDDI9rAOV
`protect END_PROTECTED
