`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RO4Z83qOL1sItWsYOZzRnGV7xaUAAohn37gUgfRXlZ+pU1momXTToUQvq1G3B+3K
3EW4otr7zYz9eCmfKtzA50oKRQtua/BLThVyTk6XKrpXtKvShq6Rp6CDS3mGsB5p
UuK54wSpFEkE2Jz6HCZTaNXY0iEZ2rbzEQrsFilpUf7XOHnpda+35Xpbx97QyZcy
y2jeIHnzl6AO4TyHlXXcar5ebHmHlN9qNpI57bi7NlOu37ZeNOJWFX7qdR/5vKu3
fcy0K/kT4xho/aSAICpihgh9HA/q89q1kqnM+/b8q21WZXjSuqVfaD1HOOaKDiOC
vrLTBUCh+4srLB7rvxD9eWH2RNP5Hiagk2Mi3kn5sdCNNh3XxZ/P6THyZeWE05dJ
kAFORp8+a+PNjq9eVd4A6Skqzt3oksCoxy4VycVKj0fgGeW7boNxCq4odMIaAodC
uTADfuqinS+bMntx4hXPglpuyxKypG+FRao+n+RYwbCAQdr15ZXix6onUQuHb+oj
4VAYE4hxKE/ZKN2g3oSnTScJmknm954YMWgCYa15+hZNi1E46DCiTpC6BIET+d8c
0j9AqSW3V/ndQ0rYtw5Qlxu6Z4iPap1zQ+DGF/SMQzwlwo+2yVAvyrHN5Tijctmr
no3joDTNfSVKYmj0gw+sXEgSRsU/bDvfAgWato/U+r7G0a5cKDDgc7zYuXIeMeCP
7PNl5iWp1DLgUf1E4uNceeECJueL/mR9HnZPp5O14OL6VtVSuYNc9Rx0mAUpc+tt
Y1ijysc8fqQbkvCQhZHIKNyyojmiPRL0g2zka7uh49TOPmlpXTQmHxl8EIrOW+f1
udEJ9s541G4s+YD24HTFZRH3EVmVAAZ31876khAJu3phqrPUyiSGaJ57oHPxXAI2
YJZha4Xt5EAKKc8YXd9QcjtuHRsIw0xvYaLwCMVqeqQ=
`protect END_PROTECTED
