`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WuWYA4+hGaaQjKfSfmwW6nnojWyhkxdeKxrlcn/XMRJx4m104d57PcGZFJKfroo3
0YYmcBHun5W32n5cqqcPVc2cGAGxQGFuqwD1MkIbjaBt9NkWT9Pi8lifddRzDCsh
3xL0ZYbT9oUe0Zvt6X+dPKXyB/sclvMYEjWIOMGLZ351PeRkRSVUrjsZ3BQDXTLC
v/sz2JojiP/TfpajRTliMWzcKDWFzkRF/PTHhIRkuDF6diadf33oWeOVJ4cQN7V1
J1Zwjo/QyBkdMtXgVALJrj7O1pQFqCgd9UgoE02f3IEZXdhorWgBSwloFuizCuv0
BzdPH8OhdCRE8DyG/5Lc+ZKAX5F0a+KpswqzQOD3LhVR7txlSI2hUqBy1IGadanR
Mkg11pAt2HzxXEzE1VSA93/lUmZ3CbnwS2uAqdAGyYHgMNY8wURpB9meOEUKhndC
o7KgGpTPJ0RDjBLo0ImviASp+mmB/GWtb3vlomuk3mFh3+K5p05hTMQAaFQbInB4
R4ircIS2+lxQza6yA4h3uPFjOiU0jGKucI5zf2GusezTJpPiHmXybN4hwTixbGST
nDENVHccMTuWBvFtBogrjqOEi8h9lB7KMMRpkrMRTPFodVdM3rCA0GT+g0JKNNEb
wAkeREB5TFga+uaWm5K4xVHgZOeKtaiholirGYyqu+N8urOmq63ZE0kaPnjPgs7I
sQUF05njO6idlPMlRamrbiPeIcAId6RSE6hAuyyPWiK9jtJIQTmy++gVy7GGbJH9
mDuPBBE7IjtXGYzhVbZVeycoQgevOYwWHBTEs5/YZQmNS0Kta0wsuAx2lyp3Na5q
3SISwm+opTQyXIuW3rz+W9pCHLRGx3+kyVipyyfukwSdWNLNXHWcxE/rM34a188X
p7JPpIo1NbETdAkjUjlniuy/jUrtXyD2pqvETpoO8ppZ905cRfVHgdodZ3eaA+sS
7HTTd5f69xMjoH/DKjVlNTQu/bLav87TZHYfkOhSvFDMzW0/iNGdKh8NisKGAHOk
sNKLdzRWwKS3QrsqiaExn+jI2iKUokyFapPejo2JYUEWzP67XTlPRGgIDjREnjgB
GdeJnyD1qqSqXK27i15Lznw4WO0oilwNQCp4ieyNLUzbPlootkfCpdtCjoVhscB6
gwHhnbvpiVvynck5M614bp1nINySJGz2aRWU5H576pe0sib+4NuNwiDhdhVigIo+
C3PPqHLBKKcdWPjJe01PJiqua+dSsnN1MtVcQBeCmYG5omJWoIMlT0iz2/YzIJUu
AI6DSmisT+ssIzJntwaPyGHl2MGRruiwsPielnWLDTGkAehtKcMsHDZSvT8HgKT7
`protect END_PROTECTED
