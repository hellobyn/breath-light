`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waYvWsMFz+4pCRFJ/OL7PrLBGvnHXs644KrYJmtnBCY0fOY2Td56op87wF905TzN
yHy8/KpZH+iki2owMarhseSbrVTOJjg9abY8q/gDyy7hbgCa2gR3T5ZYRml1WCIb
0zg7Tjf+XKdgSQHJkcxsjhTeIrw+Z61wS5pVbLK6N1ha1hVGTvIK1r+FKyzvMEPb
JWkQWIsF4sWT1Y6EyVRGutyFHbwhPVqGbRqUqp1SJfXH4W1cLgB0pncQXspXmty9
NOtaG3KmtJcP3u8uG4vP6HZ7CU0SjD9IgZzPM3DdgZTu0k5sZEtoap5yZaD6Vf0z
vEHTeaJtlfVVEXMPxEHD8Y+i9XoIwl2dRhs67a8FkrydYrjE2OCR/KKgEAiMgtz2
kzLsoiGQj+kSI0kZQq32fiBtxGsSqoBIDM4AsyejrwMtg/WhH9qZ7k5PHhZCfo9r
e49RpOwxuUvj6iTjGdTMagSfjktNago7/Qs2u2a3OWRSpO9Pf0AAYkHvOZ9JCNZg
u0PNt0knu7mfd44OyxJoTSAKc3OGrTjJnvHSnM1RNYGdkKpR+L5NfbABUJumPU5G
lWdEkcudbxYMROQpr0an1jUtjfvtuhRc+AyIzbjH6eHaOvCWpliPixCbx3gP+JP8
`protect END_PROTECTED
