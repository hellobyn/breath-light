`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eE7y7jPdBoWlOD1tBxhLwZufq8gqrkC/gXnCP3LIbRomJ6y7MOaoNmZY7IPH6Twf
gxroNcXN83Rw8zBH6hzmIE47hraECMRaEKMQkirHa8ytMOGAIh3Ju1EgOlDSsYEl
gOAt+wo3pW++E2X5KVpgX7OkGosXxy8sG33hl9oLd5gCIyRJR09Z2OXda98/xXq7
YLaQVgQNOu/NjVIqAeIzjRcAOTjZdRJ/eOt9R0sGoHmXd5pO9mVQdq3Ndukn7cLt
/XniUfo+BJDNC9dd9C2shQ8ZMZIdUBMkDuxDCz9rmA0lD8F681/Ut61yuqoCd37/
jYzMOpw4QMW1JdDq1V1zKLM3t3hJaxfPh1p+xvtUKvm2hsoBBABpEewsFeUvF1Og
cA2N+qdeHt2FBNtA/8GmHaMXapvTteCVkEd+RlhiFeaUr8gJmNE2zkH4NbuQty2c
2Dp/2DrQQzsZrcJqLiwL9urSRd94dctXgcEM4pLhKIb/VmNpSojicmEdjeBec71u
Jn/fTQ+TwxZLZ35kR1Y0b8hEokIuOFy/ryfXcTLmeG6BatLmSkgWsxzUQiPzsBUm
J/lhSbzR5HXEeiep9VFgPTMnF/95/4QKq/kJXPJqxZE1qsJofJGFV0KdEOeubHkr
nNsOQF2Ugx4ogrnHGTGnCddxL2XTcuAoo+Lqs+2bATYP1MvJIDMX52TQrQg5Ag7g
r4QEN32rd/2s0C7FuQMq37ZYiXLyzz10Q3eqBBJXhBAICEsSAzRl0FuXcYDvG7za
boEUR1GOGWMiuRkQ7DR9M+4u/89/0PlwcXr+ODeWGJRH3Fv7AtFK7gRaYaa+U2IS
QBOWagfydi81x19P1hLb7niJxuNXP+e2HTnVK0iL1Aly5Wl9FlnJG/7Hc+gilNgG
/OVmM9XQum93V3O7NrV+ckGZrjmFswP0cP3ZcOiIY6d0TOawbNeFxlYyajU0HsGX
Vih5adp7U7YO65kKKxeRcqJ2r/F8SsIVKi0oYkaXlAeF48M6Ja43B4qngWNfz6qP
2/NlVx3dKrk+jPuYKMlTfRsU1KHewFoshI+PFXG1QRaNSclCfck1Jdv+m/NDRcJd
nZGCaL97zN8K9lcpMIj3UJUBVrDHq65u5yRJ/GYcLJ74Dzs8apvkW95wasfohxyH
15U5/tPeuhQ0pXWmlLhxVP5oSwGaGCBYFVcI2dFrwMjzsnwx6diZrZP//Skesvqk
+qEEvoHwIC6Y+Bfy5YP1zSGMzL7RO8yIbsSl354CIXIaICygy7X14M5lns4PPoYK
wlWLsN6/g1jk74XxVfurIQDVJ2S6xW6rtDSpvcDnrxqdL6b2kfpKStAf5g+970es
PiEE7AJiCCfqjx+R+22haM5+qztK5vkGsJtQmbwaxf5u+5YyyqbHXJFnvjG+FfJ8
igvTkRhF97aCmO3bta6d7fDXdkqUzsnODWzs8OSfpfYuGuSmL051skT8sjlsZKQr
yFOiJ58kikMhCQHOluakvdLM5SPWU0I21u0KVu1sfRMLqFAfRXWU9ifScF8oUJqU
8i4/P3c7waorvgQYnJTvP05uzbCkJgmrjXUFyY6EVfxtes04kc9wElA6gTiMtGMv
196AOqG9Bw/1EfCrKbYdwbTOUmuHpbL/lpxfsZqdu6BPTNOmAJyu5chUIoYYLBgv
+C29c+MLqXzlcrk+acWOIEbo9hMALlidysdWRiBnmmOoNxr1dMz05AbhiK2YgdP7
eaehx/JI7hAcKMGsdFIEmRnhAj1D87SFvIgaVGTmP/yfT1Gaw4I3Xg+0Drgetkzc
wj1Z0+5k15vb/E14+TUPqKUeTCySRE8I2z3pEgByQD6I0fMv73Vmeo8BfFXPMRzG
rAsLSqfGkQ48Ka5B5Vt6gX1y2rgYzmMIgR1oX63HWPCQBIoz/82gwdij0BQ0WLrT
VtD7shnyUhvyGgZo1ugOEC+rmVAaHKGpZZiUrmPBtl8p/geT2+0xWpzrxsKrHSuX
pUjfhpezHDHMocIoXEIX53KVeZwazEmT+H5/KjFnCwk010zXvCCWFRq5Z5SasH7A
55gnMc/WVxFcb0nIPezaxTPyvwjiu9l4XzfH4BenK8y/adE430rxbssXDWs/MyqO
Sa8ghsjX5xDnh3W8dgLuYjXsKJEr/YwKSCsSMim/kuvJqC1NLhfvsWm0ERMi6n+n
lA2K4ZMvruunWGHe/ZtkvvJJD1BthDPbWOCk6jaNie5xeGGTKBb7gGPsOuPKLlWA
NCaeOG+1la7KXbVzy6806EpmEeLFh/3FyYaZK9YIlHF9ZFzrMlHYe+r5+KnJ+WMK
wPFYKszPyuRZlq0AavQKWnH4Bf0XMKsb/Be/Qg47IMK3VjoWnJdgib+zTpBJB0QH
Z1xYxfweCW66zqecvflzfwDq/sUgqpGz3ByZD4e/A0WaDf55SJzxKrezNOCNzmNk
7erPdAqog8mk/CESdMuTu6nBuX2PWBWZRBSSBPOrpUiCqA1tEl9qz2Kv4LOqzkY7
u9YNgoG8uiGuSROfWDv5+T851xAPmcDKlRsa6GMGSAMmeuNmhe3N7ZAGSSt9bhsU
7+nI0t/J2z8grCHR2R5Dk04Nj477rzhujxxw1Cz7PIsecDQXuDdwG5u+89Tc1q/r
AVzAPydFpkdopXrniMHnyQUXpKQ+BajDiKbgFaKiF6u3waukHeWLQCiz1f3rmfF9
+w+pnfjVmnnzTtLHwcjz/ZkZjbzcbe4mK386SM4V+FAHJKUfPkrkjyjab4GcmZVh
uzXV9zdiFZOXc0EKq3HIlJFSCqA+qY2eoQuSqou3lTteEnckJC6nQJeqdGEbJNLU
8oAk/K+4jxqzid7jVqkkSyR1LphQhXD3rmFFLPy+ugsyjhVDTvZ/QxZJUPbOoVo4
uqpPCRCzjksZnNUmAt1ICJ5ZX/u11ZLub3NUtYLiQ3ZcokfBRJ2TeOMX5bIJHOpi
eS9w9DB5CN6zf8dsExNM4l9/GCjB/BR7cCEFJqZbfSXrQYrychNasv81ISUDcLzj
xzAOWieX62XdrvKBdzxKYgNUWJ2Xw8v4f/nUA7xcEPLMN9p57TI0AYjdLYNciyoC
RZG2c7tTm+DpAwJEQHkgGRdmR8Z+LSBg0031La/SjjeFco+3xlUh8MLS96cX6E7N
i/oabrDWYwU1cZGIgGt9GMRBeEBhQWM4PXL5IFrj5MHGBMOZigZZ5xGMqOM71sXf
mAdo3z9h0MUupx2dT5yX+bbE92h2EaG4y+qHPGecXXTVT9amlG34Agh2ALcDk6Ux
GxhxRNxc34OJRaUf1KmVJQN20VzsTldyA4UwwWaXYDu2beuvy38o25ksnqJPAiXG
3OGBluTGF6YKKiSsmQhoDvTqP3hWdnJObqtLrX68R6e4oQWoiiMXFdgrvHgXBPj7
lGxHdtTLKHxbBtoElIBkVqi3yi8XkLEQqERfWW8OF6p7uoXMlZMCwA0AEKfAru7Y
8DLnb87Cv17m9yk4qxucOfn9/5cXOaVT1bJ/FkvQ0EAPrSATWnzCAmAnT2cTbkgr
z6AxLD+NsMITZONXQg61wTKpD1EgkQyh5+lT43pZkPvl3HVSKF9+BsdpSE2TsfKO
+BvOHpOsFxQ1vupsQem9ciCi1ceUUxsniltUl4nLlJ4r2Jrod4RmDoDumj2FJ1c3
i8yu5Xs0aJA3CLIIXU1kKgEId+DDkU9m0nEIyOHf7NU4XM3SidseeV4rcAuLF0f5
U1EnfAUx7SJEDDnBCWZ9bSbGzJ9DbV31Kg/DQ50+p3E+bV206N11Dv/lxcA8RVM7
WjG5HYj5xh5sALTTYjUN40c0QYD5hgR3soz0E79VHOtVC1p4+Xl6VVM2HgvzjE4h
ABakf0c0vaf8w/sooZqRurthnmStMfADB1Vnd2OG2+DmJgDbA2AEHrKjjnuDf6cI
9gkD+aBFeMqw1PDOhUsC9UoGjJiLOS9fKLo92xTHgXiLZd+OJD3OGyBP3JaSmzj1
hwHizHqQiVpql637ONCfWUmD/L71sqk/5/rEtvfRbOJDD+qwlDTFpCWIUK4h9YsK
kMOou6BPoHOxEJ8bOW8L8Q==
`protect END_PROTECTED
