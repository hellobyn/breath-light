`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3yYbGfIVM0vQbwED2GXQKv7daTiAR5YepcbXjg/QV+bhJx2iLkPWrz0xPYqR7Dq
/rk+ckXFuAHLjXdRDCuTRVaXR1g8PnEPvXUuGGuAb9emhfoZttMnfHRygtU0HUy4
JM4qonWMU0Kd8Z66HiTdMWHLQfLIAP/4WkKBPIE0hUqr1V4PJd3dI9iYtx2OhDgU
1m/OhrCI7WE+GMXvt86jRsfExHn790cSx8CvhihIM+sEnrq9CWYIp31I+pFqYSH+
BBmnrU3CRoYIXmSyXWYGOZd2PNEzlHKS6uyUU4xSDf7gPd53xcgUNJvc04pw44Rl
HpmsnGbOcYcCsftpPwcHloLZougUU9t7ULJHPlgagYE2GeygB7o1IR5ijCVowRNA
8PnC+G6Ihel+zLh1mrgxdqwkzmC6KgV7apQM97RKXnZUTNfZS05721SW+CHtZ0yY
DNW+CvxHP+iZ/Kl5RcJnV59ibEWLSClzOy9HBwDDKMA7nKCBoCRXcMz4pBRVYY3W
IEPDRv6P7ykg8uNoDh/LZORCiIQ5yJ4vUfrg1dSE9mbU7vUMts4wciamO4DvMKz2
Gto4MQRL9ziXwgUMRG+yTLeaXdDPChE1XQD+vNwzTAdgV9lcmQPhM5ecF8mORY8K
z56G0pbeWSO3dbkGCbJeQQyeDoxeQENHMHavbgblHh00Tsmbie+FXL+a2daxlFn7
VYpGU3sty/LBZqZcn+aqD7iFhb+qq23O3/U8f4cM/fDkOanrjr+Oy8CnteN9MDm/
fpKtVbJpHM7ltAGsyrd4gly5tUBI8Qy6dx2VRUMZ+Uzjo9qH5ONXQLHo3xrGUYdO
repTQZq+P8jGpMqjb/kiSCek6KoFVTDAZRFLMjykuzyO89GPjlCEF6G/A8sYlIHy
jq0oSE3FImIn7I2Gd/DG9JdokXehAdaj0Pa7hG0dwnTypZx5X4hasvatdWleT0FZ
O2QYHI4uCJNHTaIkfgBO7jobis+ohrMkPD/Dqrywuowt5eNR59MJ9BiCrAM/yOTl
u+QiJ8n08v7XaWoDLMB1FBbU58gplENe+JZwFOVbno0IIXtk3zvGtusUuhR7IDQN
f/N8jkoTQSdGByWtoKTbjJ0eNCASE/uOVIThMo8cb++uR0+adF+3OZ0fw7hw4wFa
qbwkXlfLhgbEQv7pR570JY0VjbPPpzBuMgEUvOfyZA/pG7x7hOPMgOCSISUcGUFE
oBZBlAD0UZJAqdGNT/nYEmJlLM07aDFHy1/QonMqhKeKbbh/1mVJFebuAr098GAZ
Q5yyE2taKu/3nQRohPg1awALiLaApBCnorHq9Zlaczm32GmFBoZ77DijgzE47PbK
sMEblYho9QjP9GsqK1WLRW+12TH94QkGw0hxGP/a7q/C/QlQ3wyH5ulKsxTmCiBo
NSGfe1CxijcNUSEZd3ceT1aDt8OxeDjtoFk9Hfrn1/Q=
`protect END_PROTECTED
