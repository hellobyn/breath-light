`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBGGYZDySseU5aITZaod2E7fUlcKIW63gMssv/PSRddfvlk54+jGgt3Kdyb7oNU+
bt1GtydjlTVyzl9VSI9OB7qnMOijuuvNPGVZgHnR99jdur3RMMabgM/qkccvF09f
qL6R5kiRPiCRdB/5OVl9vQXk55ok7IhBI9wL2gWul4x7KPOeyvb8+nYOzYBB8K1J
BNWuZRi8jz7CgisLdW3lUqDlrqiVKBVbDSUXGsfrPCo9c/qpIGVC0mkAglc3vzaw
9u9DBYp5zegypAEHUG2b3Q+SnxBm3XsXaTcd2qZeORcd+dvF93RT2quAZ14miTLC
m+d3ZPYGcWO1CkURs6luJe3j0wfThtd1kEwAOSYpg5h88K+iGOg0sjGErxGUrRjg
xiTY3G8qTCKBrPEUEukQWAKLkXRJxochvSKTBSONIUdXbdVMQNw+IvGZgm9O3qAO
9wRxmyHGyH+F9CxYhtiquEdUWRS17oIQgdoGTLefl4E=
`protect END_PROTECTED
