`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdHVeoxVSS2utt8QgyRNBL7NT28jUppZSOU8rcApVITSylRnLD0MxGxypJTmvC18
6I1lReKphBooKID0CQ7KuYOXrFwbzQy8KcOJv8igG2KZXJ5O0ze61wZEdQBPbbBJ
EZsh4ipZc5ApB9MHjbqGlIHiv9Z4O8UdfHO/kwMpbsu1TH/396iI+/g3HVDZ7hjo
x8oD726hp41aXGr5nJS4UUxZa1cCSgVValY6vHImiq5d9smT+p1CAnm9LwtEfKFI
PwVP240zh8n45cEW4EZxjM1mL2ns0ScocfxJq4cCo2MYyLDIysqaZpjP8Ivk1d5B
1SHlIICMQv4XivCIl6vPU6QnmBKokr78HwVwS3vwOvlBFvzggECxKKFs8dWFsFKQ
LBUe1jlgtOi8qiLNWfvxz178kGdpEoVDALpfBCKzLykiTkIG8k80akHi4JNbs9Pz
XVzgPD/mJ6TyFDNW4Y/aYDvgp+8JBTwB0JK382ftGHeCuvehzPIbp8upBp5yUTX4
yUDkfaPS6/irDaSwAVlGaOtrePB7YOrEYUMNodRbX4dzpKgWZ1M3ziXRYLiicQ9z
bZCtwbRXaeunnenGHcPfoyCLbPKwJqJeKwWRloDSNgE=
`protect END_PROTECTED
