`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlnE8KG88xc2eeOhqPTzUZX/cUNoprVwGq1jlFDzv5bJogdO40SF1sec6ZTUbobk
Q/PIrUYVfRDKA1c9RjVxagbAAwlED+Mxe23gegaNYORIanpGOEC9MLSGJV0SK1Ta
TdQ4Xzo/byc9wsNC4vcAoCpcQZlozKYz5omWICHbch9yJO3fKbi9J9Kl/cccXjCF
osg0IWAeU3ioTFyS6KBlqhSV6SOI/qmj9UhfS2onRt/LT6/ZCDPB2KUzCVIeeWcI
mxjAKGSSGKS1H/Dim+RQNxojHsqQS2uT4lOpNgb2Icxx+icshpV7g2L8K8uC0LM4
wo9ln+kT4EA46RDMCRmD5XhDHcP9l6sb12oYGR4/WNo5Argg1H9lk3rDp+Y0uW86
NHLyhFo3fyZtYNFsDjt12A==
`protect END_PROTECTED
