`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kB3FaGw0n5LonVD+ccIFlK0h4H3SYIrbuUaPfkdZ11QWMmtZ44sY/6uums8jmiYZ
Xt5aKIXCm74cxBsYmYFaIzmVub5+hNoLlsaJ0DTbrDoc45euqobm82RpW8Od7YRd
t9QRSO5ukL1CjRMGR+Y/Prb8Nuhoy4/IX26AYFMvNMIAtaJW7BcX5z9Dp+Mtxjah
58z480J9syJX9Mk5AYaFcYxCze5hSIsAguuapj/FyRbigZRSayRVKdYCl/me+AHk
ZHZCs7y/N3wEE/q1RtaXnOJkaX/68L749hP3Or8yN2+DAeJB1ZbKaGl93vENDZ2c
ADQMTd1VWAAsfa5IFNDrsrUKa31zLXdUYyRE2dmYVV6iZrq3OKvFuJpX0umjEI0w
Za3nO25HLNVSdvS1ed8cgQG3M9U1pvEGlO1bNmBSwPPY0G0dcnXnjsg+6XnM2oeS
DboxIfRrxCGJDw+WuP9x2UjZUPZlgaMlB1e9GUUdexsTeEcKYEtPytHv3Cuo0Fm4
LKBjxdqPoKsiPJ87CZY0EdmR0xtWwQ6IB3fW96qoPl2CndYXCty3cHZaWXKDiC5x
p6Nbm9EBolS6lRHMiJHb2DjTAOngMOCglhv7XHz6Veb7RtvgFDWz+a9SZsbpkSBE
WA1KxyK9EYaKscsUXMasAwm2uHTK1nXGRT31Hrl9dmlAhjBtZPCC6Q8nSKXM5+7K
4x2gQwnh9hFnfMHXuegBimxu7CkaIsQj14CTUPGrglSXbtCamvDwRRVusx76E1WO
CNTBH0TTaBXtxO16VRa+1DQB6H/aVlUbQEsn15YTc2XlmlSwMOLHNDoIzUXHKSCt
mRIyN/S2HJJtFBY9t/qRoXP/vzPrkqUZ9vEc4NjUnuuVMw1QaTOQva1Nrkn5PGa0
X1l2Lb2BnYw63vo14prX+zw8N6/oWQZ0y/mKNGv7nzxIs9JU8tqWgaUl0UlQYIhQ
08mLu9pN1FoLN8X6Ns6LhRDUaHKsuHOYcuVPhaBuh0abfEXcd4EHWLIrvlf2WhKc
EhmELu9u5EYWrPjonGoa9F5XoW1SkRAHH4tZxAv0TBiehqhuKxlxaYjSo8JCdjwj
YhHKzOk4iEauqBmBVVqm8j7+W1ZegJYo6cWUYHo6hcElDvU2F+pJ/vUbVY4w4BpM
ujc3/Pvvk7AqUcVfu5l+rzV/JYf45SK1skDUYBdXJbZlsbgXvIPDv9djZi1NOMnL
91468rfY48BhLgTsMl2VVCwc1jM9ARSSYs0Uoj5jZKwPM1Zl+5Mk2kOqpfPcFO53
`protect END_PROTECTED
