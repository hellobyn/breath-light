`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0SmvdNdjjn3Q3tUbRsRcPURkvJwMlkIuGtVgtrkAYJD9gvNV5Qf9/pYU1gWbSlG0
SNb+Fut/CksW8emauChgJJGnY7Ysr50Rudn0DNm8vOZTsFZWtwYcg3hSGduPg4hw
zmHT6asMGENzgsja62rxrBji+rA0VhOFYFUtKvD8uKdTU+qMxlm48t/o36YHeUP3
SSwFytmjLsNSYar2nMPx9eMH9FQKO3r+SaSfN6kfmNAgoMOqBz22PAT7E6OPL5vd
aaD4p8jeTGC7PcX0DuWW0XdoIHam9fNCz2CbNpB9QMerBeS1JdzZ3ox6jmV3L70C
euUZFXYyoSO4R2bdJg1JWnf2kaMMVywO9JhbsSRVGr/MS9d1apEE4LuxXBMn4ate
8cKbHCEA/hH2mMrV1/RhPw7JRWNtp42nYbODFwxZ8OZpm/lxNZ1g5j7ztsPzUpeI
oZvDWkmKFH4diVCuAsTjsMsj9CCmfOGlnzqWv1187rvKS7+n94sIabBHI3ZIzbTd
/9cjR8oRd7wJj/x3feGNvtGf2pGODWbBiSu00/xksMcc5cYg8bzkgqmXFbr0Xkq2
tcUBML7BqtWrOmMR6ettaZcuG21liFo8Zfu6cSHyBLMXhZIpoHpx2KJXsf8b5vw8
grAJyxS3Wv+deW58g1z47wD0HM4LTYGY6ojd8+95d9OVi8gb5eO1r3zgzrunAJKF
VgXw8D9QvTvbQli2yUmmI1cVNtpwjuq9/3tAndwDILz0WaU4L9JdrOVMuI2t3CdJ
xzGvkKp22VXkureD4e+/uN+l81PwWeq/JaXbsFer5nvByWiZOXen9i9aUPunNEh1
ro3tm24NdXF9kQc7HtGXQmf5a4Yi5hXuusC7EhM5fIK9uZm+CzgVTk9/AQ86/rmu
OoYRaeCwiXULpGIzksQ5WLfCiy6NFB+JLvqUxlMQKoO7ZH5evsqzGh6NWaO2+GoJ
ML3EAHuAcfXgTSZIfv7jZLeY1zShrLlnXtjGdrKbXNSFHt1qruOFfWnHcXGmsnUS
RpOofcRjDKoJOJ/UpcQpKa9Uv/PYt/bd7SuYgM4QNalbWcFeRY0DZn7xSPQBu5J0
liIyQmQhhF2IxybHoiTr/csoe1lZmlTzUUm/HiUB1BVIfnPW60tL7hkuhR1B+etL
VMXFKNWGNLsaIBKDX9g83vlK+geZmlaEAF7aw6nW+UgtbVCTaPIf9gWpA9fQy8hB
Zh7ceKMp4PR8ElcR2CTjYqw8HXLYr/pu5WQKbBoYDmwcCqEEZawSuVoV4/9dW9M9
rpSa1Mufoijja0LguM+50y4h4A76KcjXNexNFg0ok7g0stDXm7G5t05aF9c1rNAc
fmwpUtoOg7eECjtfVHXFwlTPjoyqNbs/+gYin2jRKWdgXZXeze9YUis8CKxOeGsy
9+O5JQ6/NQmd8/Zo8rQ2jkPg1GqF8cslJ0JbjPVMsSO0qtGfojpYf6trxNdJoGmb
9t63LJXDWG6x57ZYoDrGMg3lp0MjBIlvzNufI5jNynX8hdzv/y8Mg3mwbuEpzvFD
MKkm6CF0uX0/8zfR3G5GfjTjhXTzx/mcrweoFMU9HT7cZXf9VRugBzr4CzjF8V1F
fsrMxq4Cdh6iiDAngmLdQ9pWhM1ZMdUZzBRB/+BUt5o=
`protect END_PROTECTED
